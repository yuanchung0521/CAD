module c54321 (N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413, N1414, N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503, N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513, N1514, N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563, N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612, N1613, N1614, N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664, N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734, N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804, N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1823, N1824, N1825, N1826, N1827, N1828, N1829, N1830, N1831, N1832, N1833, N1834, N1835, N1836, N1837, N1838, N1839, N1840, N1841, N1842, N1843, N1844, N1845, N1846, N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854, N1855, N1856, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1885, N1886, N1887, N1888, N1889, N1890, N1891, N1892, N1893, N1894, N1895, N1896, N1897, N1898, N1899, N1900, N1901, N1902, N1903, N1904, N1905, N1906, N1907, N1908, N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918, N1919, N1920, N1921, N1922, N1923, N1924, N1925, N1926, N1927, N1928, N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1947, N1948, N1949, N1950, N1951, N1952, N1953, N1954, N1955, N1956, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1964, N1965, N1966, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976, N1977, N1978, N1979, N1980, N1981, N1982, N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, N1991, N1992, N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, N2001, N2002, N2003, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044, N2045, N2046, N2047, N2048, N2049, N2050, N2051, N2052, N2053, N2054, N2055, N2056, N2057, N2058, N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079, N2080, N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2089, N2090, N2091, N2092, N2093, N2094, N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102, N2103, N2104, N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112, N2113, N2114, N2115, N2116, N2117, N2118, N2119, N2120, N2121, N2122, N2123, N2124, N2125, N2126, N2127, N2128, N2129, N2130, N2131, N2132, N2133, N2134, N2135, N2136, N2137, N2138, N2139, N2140, N2141, N2142, N2143, N2144, N2145, N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153, N2154, N2155, N2156, N2157, N2158, N2159, N2160, N2161, N2162, N2163, N2164, N2165, N2166, N2167, N2168, N2169, N2170, N2171, N2172, N2173, N2174, N2175, N2176, N2177, N2178, N2179, N2180, N2181, N2182, N2183, N2184, N2185, N2186, N2187, N2188, N2189, N2190, N2191, N2192, N2193, N2194, N2195, N2196, N2197, N2198, N2199, N2200, N2201, N2202, N2203, N2204, N2205, N2206, N2207, N2208, N2209, N2210, N2211, N2212, N2213, N2214, N2215, N2216, N2217, N2218, N2219, N2220, N2221, N2222, N2223, N2224, N2225, N2226, N2227, N2228, N2229, N2230, N2231, N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259, N2260, N2261, N2262, N2263, N2264, N2265, N2266, N2267, N2268, N2269, N2270, N2271, N2272, N2273, N2274, N2275, N2276, N2277, N2278, N2279, N2280, N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2288, N2289, N2290, N2291, N2292, N2293, N2294, N2295, N2296, N2297, N2298, N2299, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2369, N2370, N2371, N2372, N2373, N2374, N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393, N2394, N2395, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414, N2415, N2416, N2417, N2418, N2419, N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435, N2436, N2437, N2438, N2439, N2440, N2441, N2442, N2443, N2444, N2445, N2446, N2447, N2448, N2449, N2450, N2451, N2452, N2453, N2454, N2455, N2456, N2457, N2458, N2459, N2460, N2461, N2462, N2463, N2464, N2465, N2466, N2467, N2468, N2469, N2470, N2471, N2472, N2473, N2474, N2475, N2476, N2477, N2478, N2479, N2480, N2481, N2482, N2483, N2484, N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494, N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504, N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514, N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, N2542, N2543, N2544, N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2554, N2555, N2556, N2557, N2558, N2559, N2560, N2561, N2562, N2563, N2564, N2565, N2566, N2567, N2568, N2569, N2570, N2571, N2572, N2573, N2574, N2575, N2576, N2577, N2578, N2579, N2580, N2581, N2582, N2583, N2584, N2585, N2586, N2587, N2588, N2589, N2590, N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2623, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2648, N2649, N2650, N2651, N2652, N2653, N2654, N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2682, N2683, N2684, N2685, N2686, N2687, N2688, N2689, N2690, N2691, N2692, N2693, N2694, N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2704, N2705, N2706, N2707, N2708, N2709, N2710, N2711, N2712, N2713, N2714, N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2723, N2724, N2725, N2726, N2727, N2728, N2729, N2730, N2731, N2732, N2733, N2734, N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744, N2745, N2746, N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754, N2755, N2756, N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764, N2765, N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2788, N2789, N2790, N2791, N2792, N2793, N2794, N2795, N2796, N2797, N2798, N2799, N2800, N2801, N2802, N2803, N2804, N2805, N2806, N2807, N2808, N2809, N2810, N2811, N2812, N2813, N2814, N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859, N2860, N2861, N2862, N2863, N2864, N2865, N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, N3165, N3166, N3167, N3168, N3169, N3170, N3171, N3172, N3173, N3174, N3175, N3176, N3177, N3178, N3179, N3180, N3181, N3182, N3183, N3184, N3185, N3186, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196, N3197, N3198, N3199, N3200, N3201, N3202, N3203, N3204, N3205, N3206, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266, N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, N3338, N3339, N3340, N3341, N3342, N3343, N3344, N3345, N3346, N3347, N3348, N3349, N3350, N3351, N3352, N3353, N3354, N3355, N3356, N3357, N3358, N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3376, N3377, N3378, N3379, N3380, N3381, N3382, N3383, N3384, N3385, N3386, N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394, N3395, N3396, N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3417, N3418, N3419, N3420, N3421, N3422, N3423, N3424, N3425, N3426, N3427, N3428, N3429, N3430, N3431, N3432, N3433, N3434, N3435, N3436, N3437, N3438, N3439, N3440, N3441, N3442, N3443, N3444, N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, N3457, N3458, N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3467, N3468, N3469, N3470, N3471, N3472, N3473, N3474, N3475, N3476, N3477, N3478, N3479, N3480, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494, N3495, N3496, N3497, N3498, N3499, N3500, N3501, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514, N3515, N3516, N3517, N3518, N3519, N3520, N3521, N3522, N3523, N3524, N3525, N3526, N3527, N3528, N3529, N3530, N3531, N3532, N3533, N3534, N3535, N3536, N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544, N3545, N3546, N3547, N3548, N3549, N3550, N3551, N3552, N3553, N3554, N3555, N3556, N3557, N3558, N3559, N3560, N3561, N3562, N3563, N3564, N3565, N3566, N3567, N3568, N3569, N3570, N3571, N3572, N3573, N3574, N3575, N3576, N3577, N3578, N3579, N3580, N3581, N3582, N3583, N3584, N3585, N3586, N3587, N3588, N3589, N3590, N3591, N3592, N3593, N3594, N3595, N3596, N3597, N3598, N3599, N3600, N3601, N3602, N3603, N3604, N3605, N3606, N3607, N3608, N3609, N3610, N3611, N3612, N3613, N3614, N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3687, N3688, N3689, N3690, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3698, N3699, N3700, N3701, N3702, N3703, N3704, N3705, N3706, N3707, N3708, N3709, N3710, N3711, N3712, N3713, N3714, N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3733, N3734, N3735, N3736, N3737, N3738, N3739, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3772, N3773, N3774, N3775, N3776, N3777, N3778, N3779, N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, N3790, N3791, N3792, N3793, N3794, N3795, N3796, N3797, N3798, N3799, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, N3808, N3809, N3810, N3811, N3812, N3813, N3814, N3815, N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3823, N3824, N3825, N3826, N3827, N3828, N3829, N3830, N3831, N3832, N3833, N3834, N3835, N3836, N3837, N3838, N3839, N3840, N3841, N3842, N3843, N3844, N3845, N3846, N3847, N3848, N3849, N3850, N3851, N3852, N3853, N3854, N3855, N3856, N3857, N3858, N3859, N3860, N3861, N3862, N3863, N3864, N3865, N3866, N3867, N3868, N3869, N3870, N3871, N3872, N3873, N3874, N3875, N3876, N3877, N3878, N3879, N3880, N3881, N3882, N3883, N3884, N3885, N3886, N3887, N3888, N3889, N3890, N3891, N3892, N3893, N3894, N3895, N3896, N3897, N3898, N3899, N3900, N3901, N3902, N3903, N3904, N3905, N3906, N3907, N3908, N3909, N3910, N3911, N3912, N3913, N3914, N3915, N3916, N3917, N3918, N3919, N3920, N3921, N3922, N3923, N3924, N3925, N3926, N3927, N3928, N3929, N3930, N3931, N3932, N3933, N3934, N3935, N3936, N3937, N3938, N3939, N3940, N3941, N3942, N3943, N3944, N3945, N3946, N3947, N3948, N3949, N3950, N3951, N3952, N3953, N3954, N3955, N3956, N3957, N3958, N3959, N3960, N3961, N3962, N3963, N3964, N3965, N3966, N3967, N3968, N3969, N3970, N3971, N3972, N3973, N3974, N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3985, N3986, N3987, N3988, N3989, N3990, N3991, N3992, N3993, N3994, N3995, N3996, N3997, N3998, N3999, N4000, N4001, N4002, N4003, N4004, N4005, N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014, N4015, N4016, N4017, N4018, N4019, N4020, N4021, N4022, N4023, N4024, N4025, N4026, N4027, N4028, N4029, N4030, N4031, N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040, N4041, N4042, N4043, N4044, N4045, N4046, N4047, N4048, N4049, N4050, N4051, N4052, N4053, N4054, N4055, N4056, N4057, N4058, N4059, N4060, N4061, N4062, N4063, N4064, N4065, N4066, N4067, N4068, N4069, N4070, N4071, N4072, N4073, N4074, N4075, N4076, N4077, N4078, N4079, N4080, N4081, N4082, N4083, N4084, N4085, N4086, N4087, N4088, N4089, N4090, N4091, N4092, N4093, N4094, N4095, N4096, N4097, N4098, N4099, N4100, N4101, N4102, N4103, N4104, N4105, N4106, N4107, N4108, N4109, N4110, N4111, N4112, N4113, N4114, N4115, N4116, N4117, N4118, N4119, N4120, N4121, N4122, N4123, N4124, N4125, N4126, N4127, N4128, N4129, N4130, N4131, N4132, N4133, N4134, N4135, N4136, N4137, N4138, N4139, N4140, N4141, N4142, N4143, N4144, N4145, N4146, N4147, N4148, N4149, N4150, N4151, N4152, N4153, N4154, N4155, N4156, N4157, N4158, N4159, N4160, N4161, N4162, N4163, N4164, N4165, N4166, N4167, N4168, N4169, N4170, N4171, N4172, N4173, N4174, N4175, N4176, N4177, N4178, N4179, N4180, N4181, N4182, N4183, N4184, N4185, N4186, N4187, N4188, N4189, N4190, N4191, N4192, N4193, N4194, N4195, N4196, N4197, N4198, N4199, N4200, N4201, N4202, N4203, N4204, N4205, N4206, N4207, N4208, N4209, N4210, N4211, N4212, N4213, N4214, N4215, N4216, N4217, N4218, N4219, N4220, N4221, N4222, N4223, N4224, N4225, N4226, N4227, N4228, N4229, N4230, N4231, N4232, N4233, N4234, N4235, N4236, N4237, N4238, N4239, N4240, N4241, N4242, N4243, N4244, N4245, N4246, N4247, N4248, N4249, N4250, N4251, N4252, N4253, N4254, N4255, N4256, N4257, N4258, N4259, N4260, N4261, N4262, N4263, N4264, N4265, N4266, N4267, N4268, N4269, N4270, N4271, N4272, N4273, N4274, N4275, N4276, N4277, N4278, N4279, N4280, N4281, N4282, N4283, N4284, N4285, N4286, N4287, N4288, N4289, N4290, N4291, N4292, N4293, N4294, N4295, N4296, N4297, N4298, N4299, N4300, N4301, N4302, N4303, N4304, N4305, N4306, N4307, N4308, N4309, N4310, N4311, N4312, N4313, N4314, N4315, N4316, N4317, N4318, N4319, N4320, N4321, N4322, N4323, N4324, N4325, N4326, N4327, N4328, N4329, N4330, N4331, N4332, N4333, N4334, N4335, N4336, N4337, N4338, N4339, N4340, N4341, N4342, N4343, N4344, N4345, N4346, N4347, N4348, N4349, N4350, N4351, N4352, N4353, N4354, N4355, N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363, N4364, N4365, N4366, N4367, N4368, N4369, N4370, N4371, N4372, N4373, N4374, N4375, N4376, N4377, N4378, N4379, N4380, N4381, N4382, N4383, N4384, N4385, N4386, N4387, N4388, N4389, N4390, N4391, N4392, N4393, N4394, N4395, N4396, N4397, N4398, N4399, N4400, N4401, N4402, N4403, N4404, N4405, N4406, N4407, N4408, N4409, N4410, N4411, N4412, N4413, N4414, N4415, N4416, N4417, N4418, N4419, N4420, N4421, N4422, N4423, N4424, N4425, N4426, N4427, N4428, N4429, N4430, N4431, N4432, N4433, N4434, N4435, N4436, N4437, N4438, N4439, N4440, N4441, N4442, N4443, N4444, N4445, N4446, N4447, N4448, N4449, N4450, N4451, N4452, N4453, N4454, N4455, N4456, N4457, N4458, N4459, N4460, N4461, N4462, N4463, N4464, N4465, N4466, N4467, N4468, N4469, N4470, N4471, N4472, N4473, N4474, N4475, N4476, N4477, N4478, N4479, N4480, N4481, N4482, N4483, N4484, N4485, N4486, N4487, N4488, N4489, N4490, N4491, N4492, N4493, N4494, N4495, N4496, N4497, N4498, N4499, N4500, N4501, N4502, N4503, N4504, N4505, N4506, N4507, N4508, N4509, N4510, N4511, N4512, N4513, N4514, N4515, N4516, N4517, N4518, N4519, N4520, N4521, N4522, N4523, N4524, N4525, N4526, N4527, N4528, N4529, N4530, N4531, N4532, N4533, N4534, N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543, N4544, N4545, N4546, N4547, N4548, N4549, N4550, N4551, N4552, N4553, N4554, N4555, N4556, N4557, N4558, N4559, N4560, N4561, N4562, N4563, N4564, N4565, N4566, N4567, N4568, N4569, N4570, N4571, N4572, N4573, N4574, N4575, N4576, N4577, N4578, N4579, N4580, N4581, N4582, N4583, N4584, N4585, N4586, N4587, N4588, N4589, N4590, N4591, N4592, N4593, N4594, N4595, N4596, N4597, N4598, N4599, N4600, N4601, N4602, N4603, N4604, N4605, N4606, N4607, N4608, N4609, N4610, N4611, N4612, N4613, N4614, N4615, N4616, N4617, N4618, N4619, N4620, N4621, N4622, N4623, N4624, N4625, N4626, N4627, N4628, N4629, N4630, N4631, N4632, N4633, N4634, N4635, N4636, N4637, N4638, N4639, N4640, N4641, N4642, N4643, N4644, N4645, N4646, N4647, N4648, N4649, N4650, N4651, N4652, N4653, N4654, N4655, N4656, N4657, N4658, N4659, N4660, N4661, N4662, N4663, N4664, N4665, N4666, N4667, N4668, N4669, N4670, N4671, N4672, N4673, N4674, N4675, N4676, N4677, N4678, N4679, N4680, N4681, N4682, N4683, N4684, N4685, N4686, N4687, N4688, N4689, N4690, N4691, N4692, N4693, N4694, N4695, N4696, N4697, N4698, N4699, N4700, N4701, N4702, N4703, N4704, N4705, N4706, N4707, N4708, N4709, N4710, N4711, N4712, N4713, N4714, N4715, N4716, N4717, N4718, N4719, N4720, N4721, N4722, N4723, N4724, N4725, N4726, N4727, N4728, N4729, N4730, N4731, N4732, N4733, N4734, N4735, N4736, N4737, N4738, N4739, N4740, N4741, N4742, N4743, N4744, N4745, N4746, N4747, N4748, N4749, N4750, N4751, N4752, N4753, N4754, N4755, N4756, N4757, N4758, N4759, N4760, N4761, N4762, N4763, N4764, N4765, N4766, N4767, N4768, N4769, N4770, N4771, N4772, N4773, N4774, N4775, N4776, N4777, N4778, N4779, N4780, N4781, N4782, N4783, N4784, N4785, N4786, N4787, N4788, N4789, N4790, N4791, N4792, N4793, N4794, N4795, N4796, N4797, N4798, N4799, N4800, N4801, N4802, N4803, N4804, N4805, N4806, N4807, N4808, N4809, N4810, N4811, N4812, N4813, N4814, N4815, N4816, N4817, N4818, N4819, N4820, N4821, N4822, N4823, N4824, N4825, N4826, N4827, N4828, N4829, N4830, N4831, N4832, N4833, N4834, N4835, N4836, N4837, N4838, N4839, N4840, N4841, N4842, N4843, N4844, N4845, N4846, N4847, N4848, N4849, N4850, N4851, N4852, N4853, N4854, N4855, N4856, N4857, N4858, N4859, N4860, N4861, N4862, N4863, N4864, N4865, N4866, N4867, N4868, N4869, N4870, N4871, N4872, N4873, N4874, N4875, N4876, N4877, N4878, N4879, N4880, N4881, N4882, N4883, N4884, N4885, N4886, N4887, N4888, N4889, N4890, N4891, N4892, N4893, N4894, N4895, N4896, N4897, N4898, N4899, N4900, N4901, N4902, N4903, N4904, N4905, N4906, N4907, N4908, N4909, N4910, N4911, N4912, N4913, N4914, N4915, N4916, N4917, N4918, N4919, N4920, N4921, N4922, N4923, N4924, N4925, N4926, N4927, N4928, N4929, N4930, N4931, N4932, N4933, N4934, N4935, N4936, N4937, N4938, N4939, N4940, N4941, N4942, N4943, N4944, N4945, N4946, N4947, N4948, N4949, N4950, N4951, N4952, N4953, N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4962, N4963, N4964, N4965, N4966, N4967, N4968, N4969, N4970, N4971, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N4988, N4989, N4990, N4991, N4992, N4993, N4994, N4995, N4996, N4997, N4998, N4999, N5000, N5001, N5002, N5003, N5004, N5005, N5006, N5007, N5008, N5009, N5010, N5011, N5012, N5013, N5014, N5015, N5016, N5017, N5018, N5019, N5020, N5021, N5022, N5023, N5024, N5025, N5026, N5027, N5028, N5029, N5030, N5031, N5032, N5033, N5034, N5035, N5036, N5037, N5038, N5039, N5040, N5041, N5042, N5043, N5044, N5045, N5046, N5047, N5048, N5049, N5050, N5051, N5052, N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062, N5063, N5064, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5074, N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083, N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093, N5094, N5095, N5096, N5097, N5098, N5099, N5100, N5101, N5102, N5103, N5104, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113, N5114, N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123, N5124, N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, N5134, N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144, N5145, N5146, N5147, N5148, N5149, N5150, N5151, N5152, N5153, N5154, N5155, N5156, N5157, N5158, N5159, N5160, N5161, N5162, N5163, N5164, N5165, N5166, N5167, N5168, N5169, N5170, N5171, N5172, N5173, N5174, N5175, N5176, N5177, N5178, N5179, N5180, N5181, N5182, N5183, N5184, N5185, N5186, N5187, N5188, N5189, N5190, N5191, N5192, N5193, N5194, N5195, N5196, N5197, N5198, N5199, N5200, N5201, N5202, N5203, N5204, N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212, N5213, N5214, N5215, N5216, N5217, N5218, N5219, N5220, N5221, N5222, N5223, N5224, N5225, N5226, N5227, N5228, N5229, N5230, N5231, N5232, N5233, N5234, N5235, N5236, N5237, N5238, N5239, N5240, N5241, N5242, N5243, N5244, N5245, N5246, N5247, N5248, N5249, N5250, N5251, N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262, N5263, N5264, N5265, N5266, N5267, N5268, N5269, N5270, N5271, N5272, N5273, N5274, N5275, N5276, N5277, N5278, N5279, N5280, N5281, N5282, N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290, N5291, N5292, N5293, N5294, N5295, N5296, N5297, N5298, N5299, N5300, N5301, N5302, N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310, N5311, N5312, N5313, N5314, N5315, N5316, N5317, N5318, N5319, N5320, N5321, N5322, N5323, N5324, N5325, N5326, N5327, N5328, N5329, N5330, N5331, N5332, N5333, N5334, N5335, N5336, N5337, N5338, N5339, N5340, N5341, N5342, N5343, N5344, N5345, N5346, N5347, N5348, N5349, N5350, N5351, N5352, N5353, N5354, N5355, N5356, N5357, N5358, N5359, N5360, N5361, N5362, N5363, N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5372, N5373, N5374, N5375, N5376, N5377, N5378, N5379, N5380, N5381, N5382, N5383, N5384, N5385, N5386, N5387, N5388, N5389, N5390, N5391, N5392, N5393, N5394, N5395, N5396, N5397, N5398, N5399, N5400, N5401, N5402, N5403, N5404, N5405, N5406, N5407, N5408, N5409, N5410, N5411, N5412, N5413, N5414, N5415, N5416, N5417, N5418, N5419, N5420, N5421, N5422, N5423, N5424, N5425, N5426, N5427, N5428, N5429, N5430, N5431, N5432, N5433, N5434, N5435, N5436, N5437, N5438, N5439, N5440, N5441, N5442, N5443, N5444, N5445, N5446, N5447, N5448, N5449, N5450, N5451, N5452, N5453, N5454, N5455, N5456, N5457, N5458, N5459, N5460, N5461, N5462, N5463, N5464, N5465, N5466, N5467, N5468, N5469, N5470, N5471, N5472, N5473, N5474, N5475, N5476, N5477, N5478, N5479, N5480, N5481, N5482, N5483, N5484, N5485, N5486, N5487, N5488, N5489, N5490, N5491, N5492, N5493, N5494, N5495, N5496, N5497, N5498, N5499, N5500, N5501, N5502, N5503, N5504, N5505, N5506, N5507, N5508, N5509, N5510, N5511, N5512, N5513, N5514, N5515, N5516, N5517, N5518, N5519, N5520, N5521, N5522, N5523, N5524, N5525, N5526, N5527, N5528, N5529, N5530, N5531, N5532, N5533, N5534, N5535, N5536, N5537, N5538, N5539, N5540, N5541, N5542, N5543, N5544, N5545, N5546, N5547, N5548, N5549, N5550, N5551, N5552, N5553, N5554, N5555, N5556, N5557, N5558, N5559, N5560, N5561, N5562, N5563, N5564, N5565, N5566, N5567, N5568, N5569, N5570, N5571, N5572, N5573, N5574, N5575, N5576, N5577, N5578, N5579, N5580, N5581, N5582, N5583, N5584, N5585, N5586, N5587, N5588, N5589, N5590, N5591, N5592, N5593, N5594, N5595, N5596, N5597, N5598, N5599, N5600, N5601, N5602, N5603, N5604, N5605, N5606, N5607, N5608, N5609, N5610, N5611, N5612, N5613, N5614, N5615, N5616, N5617, N5618, N5619, N5620, N5621, N5622, N5623, N5624, N5625, N5626, N5627, N5628, N5629, N5630, N5631, N5632, N5633, N5634, N5635, N5636, N5637, N5638, N5639, N5640, N5641, N5642, N5643, N5644, N5645, N5646, N5647, N5648, N5649, N5650, N5651, N5652, N5653, N5654, N5655, N5656, N5657, N5658, N5659, N5660, N5661, N5662, N5663, N5664, N5665, N5666, N5667, N5668, N5669, N5670, N5671, N5672, N5673, N5674, N5675, N5676, N5677, N5678, N5679, N5680, N5681, N5682, N5683, N5684, N5685, N5686, N5687, N5688, N5689, N5690, N5691, N5692, N5693, N5694, N5695, N5696, N5697, N5698, N5699, N5700, N5701, N5702, N5703, N5704, N5705, N5706, N5707, N5708, N5709, N5710, N5711, N5712, N5713, N5714, N5715, N5716, N5717, N5718, N5719, N5720, N5721, N5722, N5723, N5724, N5725, N5726, N5727, N5728, N5729, N5730, N5731, N5732, N5733, N5734, N5735, N5736, N5737, N5738, N5739, N5740, N5741, N5742, N5743, N5744, N5745, N5746, N5747, N5748, N5749, N5750, N5751, N5752, N5753, N5754, N5755, N5756, N5757, N5758, N5759, N5760, N5761, N5762, N5763, N5764, N5765, N5766, N5767, N5768, N5769, N5770, N5771, N5772, N5773, N5774, N5775, N5776, N5777, N5778, N5779, N5780, N5781, N5782, N5783, N5784, N5785, N5786, N5787, N5788, N5789, N5790, N5791, N5792, N5793, N5794, N5795, N5796, N5797, N5798, N5799, N5800, N5801, N5802, N5803, N5804, N5805, N5806, N5807, N5808, N5809, N5810, N5811, N5812, N5813, N5814, N5815, N5816, N5817, N5818, N5819, N5820, N5821, N5822, N5823, N5824, N5825, N5826, N5827, N5828, N5829, N5830, N5831, N5832, N5833, N5834, N5835, N5836, N5837, N5838, N5839, N5840, N5841, N5842, N5843, N5844, N5845, N5846, N5847, N5848, N5849, N5850, N5851, N5852, N5853, N5854, N5855, N5856, N5857, N5858, N5859, N5860, N5861, N5862, N5863, N5864, N5865, N5866, N5867, N5868, N5869, N5870, N5871, N5872, N5873, N5874, N5875, N5876, N5877, N5878, N5879, N5880, N5881, N5882, N5883, N5884, N5885, N5886, N5887, N5888, N5889, N5890, N5891, N5892, N5893, N5894, N5895, N5896, N5897, N5898, N5899, N5900, N5901, N5902, N5903, N5904, N5905, N5906, N5907, N5908, N5909, N5910, N5911, N5912, N5913, N5914, N5915, N5916, N5917, N5918, N5919, N5920, N5921, N5922, N5923, N5924, N5925, N5926, N5927, N5928, N5929, N5930, N5931, N5932, N5933, N5934, N5935, N5936, N5937, N5938, N5939, N5940, N5941, N5942, N5943, N5944, N5945, N5946, N5947, N5948, N5949, N5950, N5951, N5952, N5953, N5954, N5955, N5956, N5957, N5958, N5959, N5960, N5961, N5962, N5963, N5964, N5965, N5966, N5967, N5968, N5969, N5970, N5971, N5972, N5973, N5974, N5975, N5976, N5977, N5978, N5979, N5980, N5981, N5982, N5983, N5984, N5985, N5986, N5987, N5988, N5989, N5990, N5991, N5992, N5993, N5994, N5995, N5996, N5997, N5998, N5999, N6000, N6001, N6002, N6003, N6004, N6005, N6006, N6007, N6008, N6009, N6010, N6011, N6012, N6013, N6014, N6015, N6016, N6017, N6018, N6019, N6020, N6021, N6022, N6023, N6024, N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032, N6033, N6034, N6035, N6036, N6037, N6038, N6039, N6040, N6041, N6042, N6043, N6044, N6045, N6046, N6047, N6048, N6049, N6050, N6051, N6052, N6053, N6054, N6055, N6056, N6057, N6058, N6059, N6060, N6061, N6062, N6063, N6064, N6065, N6066, N6067, N6068, N6069, N6070, N6071, N6072, N6073, N6074, N6075, N6076, N6077, N6078, N6079, N6080, N6081, N6082, N6083, N6084, N6085, N6086, N6087, N6088, N6089, N6090, N6091, N6092, N6093, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6109, N6110, N6111, N6112, N6113, N6114, N6115, N6116, N6117, N6118, N6119, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134, N6135, N6136, N6137, N6138, N6139, N6140, N6141, N6142, N6143, N6144, N6145, N6146, N6147, N6148, N6149, N6150, N6151, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6165, N6166, N6167, N6168, N6169, N6170, N6171, N6172, N6173, N6174, N6175, N6176, N6177, N6178, N6179, N6180, N6181, N6182, N6183, N6184, N6185, N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6195, N6196, N6197, N6198, N6199, N6200, N6201, N6202, N6203, N6204, N6205, N6206, N6207, N6208, N6209, N6210, N6211, N6212, N6213, N6214, N6215, N6216, N6217, N6218, N6219, N6220, N6221, N6222, N6223, N6224, N6225, N6226, N6227, N6228, N6229, N6230, N6231, N6232, N6233, N6234, N6235, N6236, N6237, N6238, N6239, N6240, N6241, N6242, N6243, N6244, N6245, N6246, N6247, N6248, N6249, N6250, N6251, N6252, N6253, N6254, N6255, N6256, N6257, N6258, N6259, N6260, N6261, N6262, N6263, N6264, N6265, N6266, N6267, N6268, N6269, N6270, N6271, N6272, N6273, N6274, N6275, N6276, N6277, N6278, N6279, N6280, N6281, N6282, N6283, N6284, N6285, N6286, N6287, N6288, N6289, N6290, N6291, N6292, N6293, N6294, N6295, N6296, N6297, N6298, N6299, N6300, N6301, N6302, N6303, N6304, N6305, N6306, N6307, N6308, N6309, N6310, N6311, N6312, N6313, N6314, N6315, N6316, N6317, N6318, N6319, N6320, N6321, N6322, N6323, N6324, N6325, N6326, N6327, N6328, N6329, N6330, N6331, N6332, N6333, N6334, N6335, N6336, N6337, N6338, N6339, N6340, N6341, N6342, N6343, N6344, N6345, N6346, N6347, N6348, N6349, N6350, N6351, N6352, N6353, N6354, N6355, N6356, N6357, N6358, N6359, N6360, N6361, N6362, N6363, N6364, N6365, N6366, N6367, N6368, N6369, N6370, N6371, N6372, N6373, N6374, N6375, N6376, N6377, N6378, N6379, N6380, N6381, N6382, N6383, N6384, N6385, N6386, N6387, N6388, N6389, N6390, N6391, N6392, N6393, N6394, N6395, N6396, N6397, N6398, N6399, N6400, N6401, N6402, N6403, N6404, N6405, N6406, N6407, N6408, N6409, N6410, N6411, N6412, N6413, N6414, N6415, N6416, N6417, N6418, N6419, N6420, N6421, N6422, N6423, N6424, N6425, N6426, N6427, N6428, N6429, N6430, N6431, N6432, N6433, N6434, N6435, N6436, N6437, N6438, N6439, N6440, N6441, N6442, N6443, N6444, N6445, N6446, N6447, N6448, N6449, N6450, N6451, N6452, N6453, N6454, N6455, N6456, N6457, N6458, N6459, N6460, N6461, N6462, N6463, N6464, N6465, N6466, N6467, N6468, N6469, N6470, N6471, N6472, N6473, N6474, N6475, N6476, N6477, N6478, N6479, N6480, N6481, N6482, N6483, N6484, N6485, N6486, N6487, N6488, N6489, N6490, N6491, N6492, N6493, N6494, N6495, N6496, N6497, N6498, N6499, N6500, N6501, N6502, N6503, N6504, N6505, N6506, N6507, N6508, N6509, N6510, N6511, N6512, N6513, N6514, N6515, N6516, N6517, N6518, N6519, N6520, N6521, N6522, N6523, N6524, N6525, N6526, N6527, N6528, N6529, N6530, N6531, N6532, N6533, N6534, N6535, N6536, N6537, N6538, N6539, N6540, N6541, N6542, N6543, N6544, N6545, N6546, N6547, N6548, N6549, N6550, N6551, N6552, N6553, N6554, N6555, N6556, N6557, N6558, N6559, N6560, N6561, N6562, N6563, N6564, N6565, N6566, N6567, N6568, N6569, N6570, N6571, N6572, N6573, N6574, N6575, N6576, N6577, N6578, N6579, N6580, N6581, N6582, N6583, N6584, N6585, N6586, N6587, N6588, N6589, N6590, N6591, N6592, N6593, N6594, N6595, N6596, N6597, N6598, N6599, N6600, N6601, N6602, N6603, N6604, N6605, N6606, N6607, N6608, N6609, N6610, N6611, N6612, N6613, N6614, N6615, N6616, N6617, N6618, N6619, N6620, N6621, N6622, N6623, N6624, N6625, N6626, N6627, N6628, N6629, N6630, N6631, N6632, N6633, N6634, N6635, N6636, N6637, N6638, N6639, N6640, N6641, N6642, N6643, N6644, N6645, N6646, N6647, N6648, N6649, N6650, N6651, N6652, N6653, N6654, N6655, N6656, N6657, N6658, N6659, N6660, N6661, N6662, N6663, N6664, N6665, N6666, N6667, N6668, N6669, N6670, N6671, N6672, N6673, N6674, N6675, N6676, N6677, N6678, N6679, N6680, N6681, N6682, N6683, N6684, N6685, N6686, N6687, N6688, N6689, N6690, N6691, N6692, N6693, N6694, N6695, N6696, N6697, N6698, N6699, N6700, N6701, N6702, N6703, N6704, N6705, N6706, N6707, N6708, N6709, N6710, N6711, N6712, N6713, N6714, N6715, N6716, N6717, N6718, N6719, N6720, N6721, N6722, N6723, N6724, N6725, N6726, N6727, N6728, N6729, N6730, N6731, N6732, N6733, N6734, N6735, N6736, N6737, N6738, N6739, N6740, N6741, N6742, N6743, N6744, N6745, N6746, N6747, N6748, N6749, N6750, N6751, N6752, N6753, N6754, N6755, N6756, N6757, N6758, N6759, N6760, N6761, N6762, N6763, N6764, N6765, N6766, N6767, N6768, N6769, N6770, N6771, N6772, N6773, N6774, N6775, N6776, N6777, N6778, N6779, N6780, N6781, N6782, N6783, N6784, N6785, N6786, N6787, N6788, N6789, N6790, N6791, N6792, N6793, N6794, N6795, N6796, N6797, N6798, N6799, N6800, N6801, N6802, N6803, N6804, N6805, N6806, N6807, N6808, N6809, N6810, N6811, N6812, N6813, N6814, N6815, N6816, N6817, N6818, N6819, N6820, N6821, N6822, N6823, N6824, N6825, N6826, N6827, N6828, N6829, N6830, N6831, N6832, N6833, N6834, N6835, N6836, N6837, N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6845, N6846, N6847, N6848, N6849, N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857, N6858, N6859, N6860, N6861, N6862, N6863, N6864, N6865, N6866, N6867, N6868, N6869, N6870, N6871, N6872, N6873, N6874, N6875, N6876, N6877, N6878, N6879, N6880, N6881, N6882, N6883, N6884, N6885, N6886, N6887, N6888, N6889, N6890, N6891, N6892, N6893, N6894, N6895, N6896, N6897, N6898, N6899, N6900, N6901, N6902, N6903, N6904, N6905, N6906, N6907, N6908, N6909, N6910, N6911, N6912, N6913, N6914, N6915, N6916, N6917, N6918, N6919, N6920, N6921, N6922, N6923, N6924, N6925, N6926, N6927, N6928, N6929, N6930, N6931, N6932, N6933, N6934, N6935, N6936, N6937, N6938, N6939, N6940, N6941, N6942, N6943, N6944, N6945, N6946, N6947, N6948, N6949, N6950, N6951, N6952, N6953, N6954, N6955, N6956, N6957, N6958, N6959, N6960, N6961, N6962, N6963, N6964, N6965, N6966, N6967, N6968, N6969, N6970, N6971, N6972, N6973, N6974, N6975, N6976, N6977, N6978, N6979, N6980, N6981, N6982, N6983, N6984, N6985, N6986, N6987, N6988, N6989, N6990, N6991, N6992, N6993, N6994, N6995, N6996, N6997, N6998, N6999, N7000, N7001, N7002, N7003, N7004, N7005, N7006, N7007, N7008, N7009, N7010, N7011, N7012, N7013, N7014, N7015, N7016, N7017, N7018, N7019, N7020, N7021, N7022, N7023, N7024, N7025, N7026, N7027, N7028, N7029, N7030, N7031, N7032, N7033, N7034, N7035, N7036, N7037, N7038, N7039, N7040, N7041, N7042, N7043, N7044, N7045, N7046, N7047, N7048, N7049, N7050, N7051, N7052, N7053, N7054, N7055, N7056, N7057, N7058, N7059, N7060, N7061, N7062, N7063, N7064, N7065, N7066, N7067, N7068, N7069, N7070, N7071, N7072, N7073, N7074, N7075, N7076, N7077, N7078, N7079, N7080, N7081, N7082, N7083, N7084, N7085, N7086, N7087, N7088, N7089, N7090, N7091, N7092, N7093, N7094, N7095, N7096, N7097, N7098, N7099, N7100, N7101, N7102, N7103, N7104, N7105, N7106, N7107, N7108, N7109, N7110, N7111, N7112, N7113, N7114, N7115, N7116, N7117, N7118, N7119, N7120, N7121, N7122, N7123, N7124, N7125, N7126, N7127, N7128, N7129, N7130, N7131, N7132, N7133, N7134, N7135, N7136, N7137, N7138, N7139, N7140, N7141, N7142, N7143, N7144, N7145, N7146, N7147, N7148, N7149, N7150, N7151, N7152, N7153, N7154, N7155, N7156, N7157, N7158, N7159, N7160, N7161, N7162, N7163, N7164, N7165, N7166, N7167, N7168, N7169, N7170, N7171, N7172, N7173, N7174, N7175, N7176, N7177, N7178, N7179, N7180, N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188, N7189, N7190, N7191, N7192, N7193, N7194, N7195, N7196, N7197, N7198, N7199, N7200, N7201, N7202, N7203, N7204, N7205, N7206, N7207, N7208, N7209, N7210, N7211, N7212, N7213, N7214, N7215, N7216, N7217, N7218, N7219, N7220, N7221, N7222, N7223, N7224, N7225, N7226, N7227, N7228, N7229, N7230, N7231, N7232, N7233, N7234, N7235, N7236, N7237, N7238, N7239, N7240, N7241, N7242, N7243, N7244, N7245, N7246, N7247, N7248, N7249, N7250, N7251, N7252, N7253, N7254, N7255, N7256, N7257, N7258, N7259, N7260, N7261, N7262, N7263, N7264, N7265, N7266, N7267, N7268, N7269, N7270, N7271, N7272, N7273, N7274, N7275, N7276, N7277, N7278, N7279, N7280, N7281, N7282, N7283, N7284, N7285, N7286, N7287, N7288, N7289, N7290, N7291, N7292, N7293, N7294, N7295, N7296, N7297, N7298, N7299, N7300, N7301, N7302, N7303, N7304, N7305, N7306, N7307, N7308, N7309, N7310, N7311, N7312, N7313, N7314, N7315, N7316, N7317, N7318, N7319, N7320, N7321, N7322, N7323, N7324, N7325, N7326, N7327, N7328, N7329, N7330, N7331, N7332, N7333, N7334, N7335, N7336, N7337, N7338, N7339, N7340, N7341, N7342, N7343, N7344, N7345, N7346, N7347, N7348, N7349, N7350, N7351, N7352, N7353, N7354, N7355, N7356, N7357, N7358, N7359, N7360, N7361, N7362, N7363, N7364, N7365, N7366, N7367, N7368, N7369, N7370, N7371, N7372, N7373, N7374, N7375, N7376, N7377, N7378, N7379, N7380, N7381, N7382, N7383, N7384, N7385, N7386, N7387, N7388, N7389, N7390, N7391, N7392, N7393, N7394, N7395, N7396, N7397, N7398, N7399, N7400, N7401, N7402, N7403, N7404, N7405, N7406, N7407, N7408, N7409, N7410, N7411, N7412, N7413, N7414, N7415, N7416, N7417, N7418, N7419, N7420, N7421, N7422, N7423, N7424, N7425, N7426, N7427, N7428, N7429, N7430, N7431, N7432, N7433, N7434, N7435, N7436, N7437, N7438, N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447, N7448, N7449, N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7457, N7458, N7459, N7460, N7461, N7462, N7463, N7464, N7465, N7466, N7467, N7468, N7469, N7470, N7471, N7472, N7473, N7474, N7475, N7476, N7477, N7478, N7479, N7480, N7481, N7482, N7483, N7484, N7485, N7486, N7487, N7488, N7489, N7490, N7491, N7492, N7493, N7494, N7495, N7496, N7497, N7498, N7499, N7500, N7501, N7502, N7503, N7504, N7505, N7506, N7507, N7508, N7509, N7510, N7511, N7512, N7513, N7514, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7523, N7524, N7525, N7526, N7527, N7528, N7529, N7530, N7531, N7532, N7533, N7534, N7535, N7536, N7537, N7538, N7539, N7540, N7541, N7542, N7543, N7544, N7545, N7546, N7547, N7548, N7549, N7550, N7551, N7552, N7553, N7554, N7555, N7556, N7557, N7558, N7559, N7560, N7561, N7562, N7563, N7564, N7565, N7566, N7567, N7568, N7569, N7570, N7571, N7572, N7573, N7574, N7575, N7576, N7577, N7578, N7579, N7580, N7581, N7582, N7583, N7584, N7585, N7586, N7587, N7588, N7589, N7590, N7591, N7592, N7593, N7594, N7595, N7596, N7597, N7598, N7599, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7608, N7609, N7610, N7611, N7612, N7613, N7614, N7615, N7616, N7617, N7618, N7619, N7620, N7621, N7622, N7623, N7624, N7625, N7626, N7627, N7628, N7629, N7630, N7631, N7632, N7633, N7634, N7635, N7636, N7637, N7638, N7639, N7640, N7641, N7642, N7643, N7644, N7645, N7646, N7647, N7648, N7649, N7650, N7651, N7652, N7653, N7654, N7655, N7656, N7657, N7658, N7659, N7660, N7661, N7662, N7663, N7664, N7665, N7666, N7667, N7668, N7669, N7670, N7671, N7672, N7673, N7674, N7675, N7676, N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684, N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692, N7693, N7694, N7695, N7696, N7697, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7708, N7709, N7710, N7711, N7712, N7713, N7714, N7715, N7716, N7717, N7718, N7719, N7720, N7721, N7722, N7723, N7724, N7725, N7726, N7727, N7728, N7729, N7730, N7731, N7732, N7733, N7734, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7743, N7744, N7745, N7746, N7747, N7748, N7749, N7750, N7751, N7752, N7753, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N7762, N7763, N7764, N7765, N7766, N7767, N7768, N7769, N7770, N7771, N7772, N7773, N7774, N7775, N7776, N7777, N7778, N7779, N7780, N7781, N7782, N7783, N7784, N7785, N7786, N7787, N7788, N7789, N7790, N7791, N7792, N7793, N7794, N7795, N7796, N7797, N7798, N7799, N7800, N7801, N7802, N7803, N7804, N7805, N7806, N7807, N7808, N7809, N7810, N7811, N7812, N7813, N7814, N7815, N7816, N7817, N7818, N7819, N7820, N7821, N7822, N7823, N7824, N7825, N7826, N7827, N7828, N7829, N7830, N7831, N7832, N7833, N7834, N7835, N7836, N7837, N7838, N7839, N7840, N7841, N7842, N7843, N7844, N7845, N7846, N7847, N7848, N7849, N7850, N7851, N7852, N7853, N7854, N7855, N7856, N7857, N7858, N7859, N7860, N7861, N7862, N7863, N7864, N7865, N7866, N7867, N7868, N7869, N7870, N7871, N7872, N7873, N7874, N7875, N7876, N7877, N7878, N7879, N7880, N7881, N7882, N7883, N7884, N7885, N7886, N7887, N7888, N7889, N7890, N7891, N7892, N7893, N7894, N7895, N7896, N7897, N7898, N7899, N7900, N7901, N7902, N7903, N7904, N7905, N7906, N7907, N7908, N7909, N7910, N7911, N7912, N7913, N7914, N7915, N7916, N7917, N7918, N7919, N7920, N7921, N7922, N7923, N7924, N7925, N7926, N7927, N7928, N7929, N7930, N7931, N7932, N7933, N7934, N7935, N7936, N7937, N7938, N7939, N7940, N7941, N7942, N7943, N7944, N7945, N7946, N7947, N7948, N7949, N7950, N7951, N7952, N7953, N7954, N7955, N7956, N7957, N7958, N7959, N7960, N7961, N7962, N7963, N7964, N7965, N7966, N7967, N7968, N7969, N7970, N7971, N7972, N7973, N7974, N7975, N7976, N7977, N7978, N7979, N7980, N7981, N7982, N7983, N7984, N7985, N7986, N7987, N7988, N7989, N7990, N7991, N7992, N7993, N7994, N7995, N7996, N7997, N7998, N7999, N8000, N8001, N8002, N8003, N8004, N8005, N8006, N8007, N8008, N8009, N8010, N8011, N8012, N8013, N8014, N8015, N8016, N8017, N8018, N8019, N8020, N8021, N8022, N8023, N8024, N8025, N8026, N8027, N8028, N8029, N8030, N8031, N8032, N8033, N8034, N8035, N8036, N8037, N8038, N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8046, N8047, N8048, N8049, N8050, N8051, N8052, N8053, N8054, N8055, N8056, N8057, N8058, N8059, N8060, N8061, N8062, N8063, N8064, N8065, N8066, N8067, N8068, N8069, N8070, N8071, N8072, N8073, N8074, N8075, N8076, N8077, N8078, N8079, N8080, N8081, N8082, N8083, N8084, N8085, N8086, N8087, N8088, N8089, N8090, N8091, N8092, N8093, N8094, N8095, N8096, N8097, N8098, N8099, N8100, N8101, N8102, N8103, N8104, N8105, N8106, N8107, N8108, N8109, N8110, N8111, N8112, N8113, N8114, N8115, N8116, N8117, N8118, N8119, N8120, N8121, N8122, N8123, N8124, N8125, N8126, N8127, N8128, N8129, N8130, N8131, N8132, N8133, N8134, N8135, N8136, N8137, N8138, N8139, N8140, N8141, N8142, N8143, N8144, N8145, N8146, N8147, N8148, N8149, N8150, N8151, N8152, N8153, N8154, N8155, N8156, N8157, N8158, N8159, N8160, N8161, N8162, N8163, N8164, N8165, N8166, N8167, N8168, N8169, N8170, N8171, N8172, N8173, N8174, N8175, N8176, N8177, N8178, N8179, N8180, N8181, N8182, N8183, N8184, N8185, N8186, N8187, N8188, N8189, N8190, N8191, N8192, N8193, N8194, N8195, N8196, N8197, N8198, N8199, N8200, N8201, N8202, N8203, N8204, N8205, N8206, N8207, N8208, N8209, N8210, N8211, N8212, N8213, N8214, N8215, N8216, N8217, N8218, N8219, N8220, N8221, N8222, N8223, N8224, N8225, N8226, N8227, N8228, N8229, N8230, N8231, N8232, N8233, N8234, N8235, N8236, N8237, N8238, N8239, N8240, N8241, N8242, N8243, N8244, N8245, N8246, N8247, N8248, N8249, N8250, N8251, N8252, N8253, N8254, N8255, N8256, N8257, N8258, N8259, N8260, N8261, N8262, N8263, N8264, N8265, N8266, N8267, N8268, N8269, N8270, N8271, N8272, N8273, N8274, N8275, N8276, N8277, N8278, N8279, N8280, N8281, N8282, N8283, N8284, N8285, N8286, N8287, N8288, N8289, N8290, N8291, N8292, N8293, N8294, N8295, N8296, N8297, N8298, N8299, N8300, N8301, N8302, N8303, N8304, N8305, N8306, N8307, N8308, N8309, N8310, N8311, N8312, N8313, N8314, N8315, N8316, N8317, N8318, N8319, N8320, N8321, N8322, N8323, N8324, N8325, N8326, N8327, N8328, N8329, N8330, N8331, N8332, N8333, N8334, N8335, N8336, N8337, N8338, N8339, N8340, N8341, N8342, N8343, N8344, N8345, N8346, N8347, N8348, N8349, N8350, N8351, N8352, N8353, N8354, N8355, N8356, N8357, N8358, N8359, N8360, N8361, N8362, N8363, N8364, N8365, N8366, N8367, N8368, N8369, N8370, N8371, N8372, N8373, N8374, N8375, N8376, N8377, N8378, N8379, N8380, N8381, N8382, N8383, N8384, N8385, N8386, N8387, N8388, N8389, N8390, N8391, N8392, N8393, N8394, N8395, N8396, N8397, N8398, N8399, N8400, N8401, N8402, N8403, N8404, N8405, N8406, N8407, N8408, N8409, N8410, N8411, N8412, N8413, N8414, N8415, N8416, N8417, N8418, N8419, N8420, N8421, N8422, N8423, N8424, N8425, N8426, N8427, N8428, N8429, N8430, N8431, N8432, N8433, N8434, N8435, N8436, N8437, N8438, N8439, N8440, N8441, N8442, N8443, N8444, N8445, N8446, N8447, N8448, N8449, N8450, N8451, N8452, N8453, N8454, N8455, N8456, N8457, N8458, N8459, N8460, N8461, N8462, N8463, N8464, N8465, N8466, N8467, N8468, N8469, N8470, N8471, N8472, N8473, N8474, N8475, N8476, N8477, N8478, N8479, N8480, N8481, N8482, N8483, N8484, N8485, N8486, N8487, N8488, N8489, N8490, N8491, N8492, N8493, N8494, N8495, N8496, N8497, N8498, N8499, N8500, N8501, N8502, N8503, N8504, N8505, N8506, N8507, N8508, N8509, N8510, N8511, N8512, N8513, N8514, N8515, N8516, N8517, N8518, N8519, N8520, N8521, N8522, N8523, N8524, N8525, N8526, N8527, N8528, N8529, N8530, N8531, N8532, N8533, N8534, N8535, N8536, N8537, N8538, N8539, N8540, N8541, N8542, N8543, N8544, N8545, N8546, N8547, N8548, N8549, N8550, N8551, N8552, N8553, N8554, N8555, N8556, N8557, N8558, N8559, N8560, N8561, N8562, N8563, N8564, N8565, N8566, N8567, N8568, N8569, N8570, N8571, N8572, N8573, N8574, N8575, N8576, N8577, N8578, N8579, N8580, N8581, N8582, N8583, N8584, N8585, N8586, N8587, N8588, N8589, N8590, N8591, N8592, N8593, N8594, N8595, N8596, N8597, N8598, N8599, N8600, N8601, N8602, N8603, N8604, N8605, N8606, N8607, N8608, N8609, N8610, N8611, N8612, N8613, N8614, N8615, N8616, N8617, N8618, N8619, N8620, N8621, N8622, N8623, N8624, N8625, N8626, N8627, N8628, N8629, N8630, N8631, N8632, N8633, N8634, N8635, N8636, N8637, N8638, N8639, N8640, N8641, N8642, N8643, N8644, N8645, N8646, N8647, N8648, N8649, N8650, N8651, N8652, N8653, N8654, N8655, N8656, N8657, N8658, N8659, N8660, N8661, N8662, N8663, N8664, N8665, N8666, N8667, N8668, N8669, N8670, N8671, N8672, N8673, N8674, N8675, N8676, N8677, N8678, N8679, N8680, N8681, N8682, N8683, N8684, N8685, N8686, N8687, N8688, N8689, N8690, N8691, N8692, N8693, N8694, N8695, N8696, N8697, N8698, N8699, N8700, N8701, N8702, N8703, N8704, N8705, N8706, N8707, N8708, N8709, N8710, N8711, N8712, N8713, N8714, N8715, N8716, N8717, N8718, N8719, N8720, N8721, N8722, N8723, N8724, N8725, N8726, N8727, N8728, N8729, N8730, N8731, N8732, N8733, N8734, N8735, N8736, N8737, N8738, N8739, N8740, N8741, N8742, N8743, N8744, N8745, N8746, N8747, N8748, N8749, N8750, N8751, N8752, N8753, N8754, N8755, N8756, N8757, N8758, N8759, N8760, N8761, N8762, N8763, N8764, N8765, N8766, N8767, N8768, N8769, N8770, N8771, N8772, N8773, N8774, N8775, N8776, N8777, N8778, N8779, N8780, N8781, N8782, N8783, N8784, N8785, N8786, N8787, N8788, N8789, N8790, N8791, N8792, N8793, N8794, N8795, N8796, N8797, N8798, N8799, N8800, N8801, N8802, N8803, N8804, N8805, N8806, N8807, N8808, N8809, N8810, N8811, N8812, N8813, N8814, N8815, N8816, N8817, N8818, N8819, N8820, N8821, N8822, N8823, N8824, N8825, N8826, N8827, N8828, N8829, N8830, N8831, N8832, N8833, N8834, N8835, N8836, N8837, N8838, N8839, N8840, N8841, N8842, N8843, N8844, N8845, N8846, N8847, N8848, N8849, N8850, N8851, N8852, N8853, N8854, N8855, N8856, N8857, N8858, N8859, N8860, N8861, N8862, N8863, N8864, N8865, N8866, N8867, N8868, N8869, N8870, N8871, N8872, N8873, N8874, N8875, N8876, N8877, N8878, N8879, N8880, N8881, N8882, N8883, N8884, N8885, N8886, N8887, N8888, N8889, N8890, N8891, N8892, N8893, N8894, N8895, N8896, N8897, N8898, N8899, N8900, N8901, N8902, N8903, N8904, N8905, N8906, N8907, N8908, N8909, N8910, N8911, N8912, N8913, N8914, N8915, N8916, N8917, N8918, N8919, N8920, N8921, N8922, N8923, N8924, N8925, N8926, N8927, N8928, N8929, N8930, N8931, N8932, N8933, N8934, N8935, N8936, N8937, N8938, N8939, N8940, N8941, N8942, N8943, N8944, N8945, N8946, N8947, N8948, N8949, N8950, N8951, N8952, N8953, N8954, N8955, N8956, N8957, N8958, N8959, N8960, N8961, N8962, N8963, N8964, N8965, N8966, N8967, N8968, N8969, N8970, N8971, N8972, N8973, N8974, N8975, N8976, N8977, N8978, N8979, N8980, N8981, N8982, N8983, N8984, N8985, N8986, N8987, N8988, N8989, N8990, N8991, N8992, N8993, N8994, N8995, N8996, N8997, N8998, N8999, N9000, N9001, N9002, N9003, N9004, N9005, N9006, N9007, N9008, N9009, N9010, N9011, N9012, N9013, N9014, N9015, N9016, N9017, N9018, N9019, N9020, N9021, N9022, N9023, N9024, N9025, N9026, N9027, N9028, N9029, N9030, N9031, N9032, N9033, N9034, N9035, N9036, N9037, N9038, N9039, N9040, N9041, N9042, N9043, N9044, N9045, N9046, N9047, N9048, N9049, N9050, N9051, N9052, N9053, N9054, N9055, N9056, N9057, N9058, N9059, N9060, N9061, N9062, N9063, N9064, N9065, N9066, N9067, N9068, N9069, N9070, N9071, N9072, N9073, N9074, N9075, N9076, N9077, N9078, N9079, N9080, N9081, N9082, N9083, N9084, N9085, N9086, N9087, N9088, N9089, N9090, N9091, N9092, N9093, N9094, N9095, N9096, N9097, N9098, N9099, N9100, N9101, N9102, N9103, N9104, N9105, N9106, N9107, N9108, N9109, N9110, N9111, N9112, N9113, N9114, N9115, N9116, N9117, N9118, N9119, N9120, N9121, N9122, N9123, N9124, N9125, N9126, N9127, N9128, N9129, N9130, N9131, N9132, N9133, N9134, N9135, N9136, N9137, N9138, N9139, N9140, N9141, N9142, N9143, N9144, N9145, N9146, N9147, N9148, N9149, N9150, N9151, N9152, N9153, N9154, N9155, N9156, N9157, N9158, N9159, N9160, N9161, N9162, N9163, N9164, N9165, N9166, N9167, N9168, N9169, N9170, N9171, N9172, N9173, N9174, N9175, N9176, N9177, N9178, N9179, N9180, N9181, N9182, N9183, N9184, N9185, N9186, N9187, N9188, N9189, N9190, N9191, N9192, N9193, N9194, N9195, N9196, N9197, N9198, N9199, N9200, N9201, N9202, N9203, N9204, N9205, N9206, N9207, N9208, N9209, N9210, N9211, N9212, N9213, N9214, N9215, N9216, N9217, N9218, N9219, N9220, N9221, N9222, N9223, N9224, N9225, N9226, N9227, N9228, N9229, N9230, N9231, N9232, N9233, N9234, N9235, N9236, N9237, N9238, N9239, N9240, N9241, N9242, N9243, N9244, N9245, N9246, N9247, N9248, N9249, N9250, N9251, N9252, N9253, N9254, N9255, N9256, N9257, N9258, N9259, N9260, N9261, N9262, N9263, N9264, N9265, N9266, N9267, N9268, N9269, N9270, N9271, N9272, N9273, N9274, N9275, N9276, N9277, N9278, N9279, N9280, N9281, N9282, N9283, N9284, N9285, N9286, N9287, N9288, N9289, N9290, N9291, N9292, N9293, N9294, N9295, N9296, N9297, N9298, N9299, N9300, N9301, N9302, N9303, N9304, N9305, N9306, N9307, N9308, N9309, N9310, N9311, N9312, N9313, N9314, N9315, N9316, N9317, N9318, N9319, N9320, N9321, N9322, N9323, N9324, N9325, N9326, N9327, N9328, N9329, N9330, N9331, N9332, N9333, N9334, N9335, N9336, N9337, N9338, N9339, N9340, N9341, N9342, N9343, N9344, N9345, N9346, N9347, N9348, N9349, N9350, N9351, N9352, N9353, N9354, N9355, N9356, N9357, N9358, N9359, N9360, N9361, N9362, N9363, N9364, N9365, N9366, N9367, N9368, N9369, N9370, N9371, N9372, N9373, N9374, N9375, N9376, N9377, N9378, N9379, N9380, N9381, N9382, N9383, N9384, N9385, N9386, N9387, N9388, N9389, N9390, N9391, N9392, N9393, N9394, N9395, N9396, N9397, N9398, N9399, N9400, N9401, N9402, N9403, N9404, N9405, N9406, N9407, N9408, N9409, N9410, N9411, N9412, N9413, N9414, N9415, N9416, N9417, N9418, N9419, N9420, N9421, N9422, N9423, N9424, N9425, N9426, N9427, N9428, N9429, N9430, N9431, N9432, N9433, N9434, N9435, N9436, N9437, N9438, N9439, N9440, N9441, N9442, N9443, N9444, N9445, N9446, N9447, N9448, N9449, N9450, N9451, N9452, N9453, N9454, N9455, N9456, N9457, N9458, N9459, N9460, N9461, N9462, N9463, N9464, N9465, N9466, N9467, N9468, N9469, N9470, N9471, N9472, N9473, N9474, N9475, N9476, N9477, N9478, N9479, N9480, N9481, N9482, N9483, N9484, N9485, N9486, N9487, N9488, N9489, N9490, N9491, N9492, N9493, N9494, N9495, N9496, N9497, N9498, N9499, N9500, N9501, N9502, N9503, N9504, N9505, N9506, N9507, N9508, N9509, N9510, N9511, N9512, N9513, N9514, N9515, N9516, N9517, N9518, N9519, N9520, N9521, N9522, N9523, N9524, N9525, N9526, N9527, N9528, N9529, N9530, N9531, N9532, N9533, N9534, N9535, N9536, N9537, N9538, N9539, N9540, N9541, N9542, N9543, N9544, N9545, N9546, N9547, N9548, N9549, N9550, N9551, N9552, N9553, N9554, N9555, N9556, N9557, N9558, N9559, N9560, N9561, N9562, N9563, N9564, N9565, N9566, N9567, N9568, N9569, N9570, N9571, N9572, N9573, N9574, N9575, N9576, N9577, N9578, N9579, N9580, N9581, N9582, N9583, N9584, N9585, N9586, N9587, N9588, N9589, N9590, N9591, N9592, N9593, N9594, N9595, N9596, N9597, N9598, N9599, N9600, N9601, N9602, N9603, N9604, N9605, N9606, N9607, N9608, N9609, N9610, N9611, N9612, N9613, N9614, N9615, N9616, N9617, N9618, N9619, N9620, N9621, N9622, N9623, N9624, N9625, N9626, N9627, N9628, N9629, N9630, N9631, N9632, N9633, N9634, N9635, N9636, N9637, N9638, N9639, N9640, N9641, N9642, N9643, N9644, N9645, N9646, N9647, N9648, N9649, N9650, N9651, N9652, N9653, N9654, N9655, N9656, N9657, N9658, N9659, N9660, N9661, N9662, N9663, N9664, N9665, N9666, N9667, N9668, N9669, N9670, N9671, N9672, N9673, N9674, N9675, N9676, N9677, N9678, N9679, N9680, N9681, N9682, N9683, N9684, N9685, N9686, N9687, N9688, N9689, N9690, N9691, N9692, N9693, N9694, N9695, N9696, N9697, N9698, N9699, N9700, N9701, N9702, N9703, N9704, N9705, N9706, N9707, N9708, N9709, N9710, N9711, N9712, N9713, N9714, N9715, N9716, N9717, N9718, N9719, N9720, N9721, N9722, N9723, N9724, N9725, N9726, N9727, N9728, N9729, N9730, N9731, N9732, N9733, N9734, N9735, N9736, N9737, N9738, N9739, N9740, N9741, N9742, N9743, N9744, N9745, N9746, N9747, N9748, N9749, N9750, N9751, N9752, N9753, N9754, N9755, N9756, N9757, N9758, N9759, N9760, N9761, N9762, N9763, N9764, N9765, N9766, N9767, N9768, N9769, N9770, N9771, N9772, N9773, N9774, N9775, N9776, N9777, N9778, N9779, N9780, N9781, N9782, N9783, N9784, N9785, N9786, N9787, N9788, N9789, N9790, N9791, N9792, N9793, N9794, N9795, N9796, N9797, N9798, N9799, N9800, N9801, N9802, N9803, N9804, N9805, N9806, N9807, N9808, N9809, N9810, N9811, N9812, N9813, N9814, N9815, N9816, N9817, N9818, N9819, N9820, N9821, N9822, N9823, N9824, N9825, N9826, N9827, N9828, N9829, N9830, N9831, N9832, N9833, N9834, N9835, N9836, N9837, N9838, N9839, N9840, N9841, N9842, N9843, N9844, N9845, N9846, N9847, N9848, N9849, N9850, N9851, N9852, N9853, N9854, N9855, N9856, N9857, N9858, N9859, N9860, N9861, N9862, N9863, N9864, N9865, N9866, N9867, N9868, N9869, N9870, N9871, N9872, N9873, N9874, N9875, N9876, N9877, N9878, N9879, N9880, N9881, N9882, N9883, N9884, N9885, N9886, N9887, N9888, N9889, N9890, N9891, N9892, N9893, N9894, N9895, N9896, N9897, N9898, N9899, N9900, N9901, N9902, N9903, N9904, N9905, N9906, N9907, N9908, N9909, N9910, N9911, N9912, N9913, N9914, N9915, N9916, N9917, N9918, N9919, N9920, N9921, N9922, N9923, N9924, N9925, N9926, N9927, N9928, N9929, N9930, N9931, N9932, N9933, N9934, N9935, N9936, N9937, N9938, N9939, N9940, N9941, N9942, N9943, N9944, N9945, N9946, N9947, N9948, N9949, N9950, N9951, N9952, N9953, N9954, N9955, N9956, N9957, N9958, N9959, N9960, N9961, N9962, N9963, N9964, N9965, N9966, N9967, N9968, N9969, N9970, N9971, N9972, N9973, N9974, N9975, N9976, N9977, N9978, N9979, N9980, N9981, N9982, N9983, N9984, N9985, N9986, N9987, N9988, N9989, N9990, N9991, N9992, N9993, N9994, N9995, N9996, N9997, N9998, N9999, N10000, N10001, N10002, N10003, N10004, N10005, N10006, N10007, N10008, N10009, N10010, N10011, N10012, N10013, N10014, N10015, N10016, N10017, N10018, N10019, N10020, N10021, N10022, N10023, N10024, N10025, N10026, N10027, N10028, N10029, N10030, N10031, N10032, N10033, N10034, N10035, N10036, N10037, N10038, N10039, N10040, N10041, N10042, N10043, N10044, N10045, N10046, N10047, N10048, N10049, N10050, N10051, N10052, N10053, N10054, N10055, N10056, N10057, N10058, N10059, N10060, N10061, N10062, N10063, N10064, N10065, N10066, N10067, N10068, N10069, N10070, N10071, N10072, N10073, N10074, N10075, N10076, N10077, N10078, N10079, N10080, N10081, N10082, N10083, N10084, N10085, N10086, N10087, N10088, N10089, N10090, N10091, N10092, N10093, N10094, N10095, N10096, N10097, N10098, N10099, N10100, N10101, N10102, N10103, N10104, N10105, N10106, N10107, N10108, N10109, N10110, N10111, N10112, N10113, N10114, N10115, N10116, N10117, N10118, N10119, N10120, N10121, N10122, N10123, N10124, N10125, N10126, N10127, N10128, N10129, N10130, N10131, N10132, N10133, N10134, N10135, N10136, N10137, N10138, N10139, N10140, N10141, N10142, N10143, N10144, N10145, N10146, N10147, N10148, N10149, N10150, N10151, N10152, N10153, N10154, N10155, N10156, N10157, N10158, N10159, N10160, N10161, N10162, N10163, N10164, N10165, N10166, N10167, N10168, N10169, N10170, N10171, N10172, N10173, N10174, N10175, N10176, N10177, N10178, N10179, N10180, N10181, N10182, N10183, N10184, N10185, N10186, N10187, N10188, N10189, N10190, N10191, N10192, N10193, N10194, N10195, N10196, N10197, N10198, N10199, N10200, N10201, N10202, N10203, N10204, N10205, N10206, N10207, N10208, N10209, N10210, N10211, N10212, N10213, N10214, N10215, N10216, N10217, N10218, N10219, N10220, N10221, N10222, N10223, N10224, N10225, N10226, N10227, N10228, N10229, N10230, N10231, N10232, N10233, N10234, N10235, N10236, N10237, N10238, N10239, N10240, N10241, N10242, N10243, N10244, N10245, N10246, N10247, N10248, N10249, N10250, N10251, N10252, N10253, N10254, N10255, N10256, N10257, N10258, N10259, N10260, N10261, N10262, N10263, N10264, N10265, N10266, N10267, N10268, N10269, N10270, N10271, N10272, N10273, N10274, N10275, N10276, N10277, N10278, N10279, N10280, N10281, N10282, N10283, N10284, N10285, N10286, N10287, N10288, N10289, N10290, N10291, N10292, N10293, N10294, N10295, N10296, N10297, N10298, N10299, N10300, N10301, N10302, N10303, N10304, N10305, N10306, N10307, N10308, N10309, N10310, N10311, N10312, N10313, N10314, N10315, N10316, N10317, N10318, N10319, N10320, N10321, N10322, N10323, N10324, N10325, N10326, N10327, N10328, N10329, N10330, N10331, N10332, N10333, N10334, N10335, N10336, N10337, N10338, N10339, N10340, N10341, N10342, N10343, N10344, N10345, N10346, N10347, N10348, N10349, N10350, N10351, N10352, N10353, N10354, N10355, N10356, N10357, N10358, N10359, N10360, N10361, N10362, N10363, N10364, N10365, N10366, N10367, N10368, N10369, N10370, N10371, N10372, N10373, N10374, N10375, N10376, N10377, N10378, N10379, N10380, N10381, N10382, N10383, N10384, N10385, N10386, N10387, N10388, N10389, N10390, N10391, N10392, N10393, N10394, N10395, N10396, N10397, N10398, N10399, N10400, N10401, N10402, N10403, N10404, N10405, N10406, N10407, N10408, N10409, N10410, N10411, N10412, N10413, N10414, N10415, N10416, N10417, N10418, N10419, N10420, N10421, N10422, N10423, N10424, N10425, N10426, N10427, N10428, N10429, N10430, N10431, N10432, N10433, N10434, N10435, N10436, N10437, N10438, N10439, N10440, N10441, N10442, N10443, N10444, N10445, N10446, N10447, N10448, N10449, N10450, N10451, N10452, N10453, N10454, N10455, N10456, N10457, N10458, N10459, N10460, N10461, N10462, N10463, N10464, N10465, N10466, N10467, N10468, N10469, N10470, N10471, N10472, N10473, N10474, N10475, N10476, N10477, N10478, N10479, N10480, N10481, N10482, N10483, N10484, N10485, N10486, N10487, N10488, N10489, N10490, N10491, N10492, N10493, N10494, N10495, N10496, N10497, N10498, N10499, N10500, N10501, N10502, N10503, N10504, N10505, N10506, N10507, N10508, N10509, N10510, N10511, N10512, N10513, N10514, N10515, N10516, N10517, N10518, N10519, N10520, N10521, N10522, N10523, N10524, N10525, N10526, N10527, N10528, N10529, N10530, N10531, N10532, N10533, N10534, N10535, N10536, N10537, N10538, N10539, N10540, N10541, N10542, N10543, N10544, N10545, N10546, N10547, N10548, N10549, N10550, N10551, N10552, N10553, N10554, N10555, N10556, N10557, N10558, N10559, N10560, N10561, N10562, N10563, N10564, N10565, N10566, N10567, N10568, N10569, N10570, N10571, N10572, N10573, N10574, N10575, N10576, N10577, N10578, N10579, N10580, N10581, N10582, N10583, N10584, N10585, N10586, N10587, N10588, N10589, N10590, N10591, N10592, N10593, N10594, N10595, N10596, N10597, N10598, N10599, N10600, N10601, N10602, N10603, N10604, N10605, N10606, N10607, N10608, N10609, N10610, N10611, N10612, N10613, N10614, N10615, N10616, N10617, N10618, N10619, N10620, N10621, N10622, N10623, N10624, N10625, N10626, N10627, N10628, N10629, N10630, N10631, N10632, N10633, N10634, N10635, N10636, N10637, N10638, N10639, N10640, N10641, N10642, N10643, N10644, N10645, N10646, N10647, N10648, N10649, N10650, N10651, N10652, N10653, N10654, N10655, N10656, N10657, N10658, N10659, N10660, N10661, N10662, N10663, N10664, N10665, N10666, N10667, N10668, N10669, N10670, N10671, N10672, N10673, N10674, N10675, N10676, N10677, N10678, N10679, N10680, N10681, N10682, N10683, N10684, N10685, N10686, N10687, N10688, N10689, N10690, N10691, N10692, N10693, N10694, N10695, N10696, N10697, N10698, N10699, N10700, N10701, N10702, N10703, N10704, N10705, N10706, N10707, N10708, N10709, N10710, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10719, N10720, N10721, N10722, N10723, N10724, N10725, N10726, N10727, N10728, N10729, N10730, N10731, N10732, N10733, N10734, N10735, N10736, N10737, N10738, N10739, N10740, N10741, N10742, N10743, N10744, N10745, N10746, N10747, N10748, N10749, N10750, N10751, N10752, N10753, N10754, N10755, N10756, N10757, N10758, N10759, N10760, N10761, N10762, N10763, N10764, N10765, N10766, N10767, N10768, N10769, N10770, N10771, N10772, N10773, N10774, N10775, N10776, N10777, N10778, N10779, N10780, N10781, N10782, N10783, N10784, N10785, N10786, N10787, N10788, N10789, N10790, N10791, N10792, N10793, N10794, N10795, N10796, N10797, N10798, N10799, N10800, N10801, N10802, N10803, N10804, N10805, N10806, N10807, N10808, N10809, N10810, N10811, N10812, N10813, N10814, N10815, N10816, N10817, N10818, N10819, N10820, N10821, N10822, N10823, N10824, N10825, N10826, N10827, N10828, N10829, N10830, N10831, N10832, N10833, N10834, N10835, N10836, N10837, N10838, N10839, N10840, N10841, N10842, N10843, N10844, N10845, N10846, N10847, N10848, N10849, N10850, N10851, N10852, N10853, N10854, N10855, N10856, N10857, N10858, N10859, N10860, N10861, N10862, N10863, N10864, N10865, N10866, N10867, N10868, N10869, N10870, N10871, N10872, N10873, N10874, N10875, N10876, N10877, N10878, N10879, N10880, N10881, N10882, N10883, N10884, N10885, N10886, N10887, N10888, N10889, N10890, N10891, N10892, N10893, N10894, N10895, N10896, N10897, N10898, N10899, N10900, N10901, N10902, N10903, N10904, N10905, N10906, N10907, N10908, N10909, N10910, N10911, N10912, N10913, N10914, N10915, N10916, N10917, N10918, N10919, N10920, N10921, N10922, N10923, N10924, N10925, N10926, N10927, N10928, N10929, N10930, N10931, N10932, N10933, N10934, N10935, N10936, N10937, N10938, N10939, N10940, N10941, N10942, N10943, N10944, N10945, N10946, N10947, N10948, N10949, N10950, N10951, N10952, N10953, N10954, N10955, N10956, N10957, N10958, N10959, N10960, N10961, N10962, N10963, N10964, N10965, N10966, N10967, N10968, N10969, N10970, N10971, N10972, N10973, N10974, N10975, N10976, N10977, N10978, N10979, N10980, N10981, N10982, N10983, N10984, N10985, N10986, N10987, N10988, N10989, N10990, N10991, N10992, N10993, N10994, N10995, N10996, N10997, N10998, N10999, N11000, N11001, N11002, N11003, N11004, N11005, N11006, N11007, N11008, N11009, N11010, N11011, N11012, N11013, N11014, N11015, N11016, N11017, N11018, N11019, N11020, N11021, N11022, N11023, N11024, N11025, N11026, N11027, N11028, N11029, N11030, N11031, N11032, N11033, N11034, N11035, N11036, N11037, N11038, N11039, N11040, N11041, N11042, N11043, N11044, N11045, N11046, N11047, N11048, N11049, N11050, N11051, N11052, N11053, N11054, N11055, N11056, N11057, N11058, N11059, N11060, N11061, N11062, N11063, N11064, N11065, N11066, N11067, N11068, N11069, N11070, N11071, N11072, N11073, N11074, N11075, N11076, N11077, N11078, N11079, N11080, N11081, N11082, N11083, N11084, N11085, N11086, N11087, N11088, N11089, N11090, N11091, N11092, N11093, N11094, N11095, N11096, N11097, N11098, N11099, N11100, N11101, N11102, N11103, N11104, N11105, N11106, N11107, N11108, N11109, N11110, N11111, N11112, N11113, N11114, N11115, N11116, N11117, N11118, N11119, N11120, N11121, N11122, N11123, N11124, N11125, N11126, N11127, N11128, N11129, N11130, N11131, N11132, N11133, N11134, N11135, N11136, N11137, N11138, N11139, N11140, N11141, N11142, N11143, N11144, N11145, N11146, N11147, N11148, N11149, N11150, N11151, N11152, N11153, N11154, N11155, N11156, N11157, N11158, N11159, N11160, N11161, N11162, N11163, N11164, N11165, N11166, N11167, N11168, N11169, N11170, N11171, N11172, N11173, N11174, N11175, N11176, N11177, N11178, N11179, N11180, N11181, N11182, N11183, N11184, N11185, N11186, N11187, N11188, N11189, N11190, N11191, N11192, N11193, N11194, N11195, N11196, N11197, N11198, N11199, N11200, N11201, N11202, N11203, N11204, N11205, N11206, N11207, N11208, N11209, N11210, N11211, N11212, N11213, N11214, N11215, N11216, N11217, N11218, N11219, N11220, N11221, N11222, N11223, N11224, N11225, N11226, N11227, N11228, N11229, N11230, N11231, N11232, N11233, N11234, N11235, N11236, N11237, N11238, N11239, N11240, N11241, N11242, N11243, N11244, N11245, N11246, N11247, N11248, N11249, N11250, N11251, N11252, N11253, N11254, N11255, N11256, N11257, N11258, N11259, N11260, N11261, N11262, N11263, N11264, N11265, N11266, N11267, N11268, N11269, N11270, N11271, N11272, N11273, N11274, N11275, N11276, N11277, N11278, N11279, N11280, N11281, N11282, N11283, N11284, N11285, N11286, N11287, N11288, N11289, N11290, N11291, N11292, N11293, N11294, N11295, N11296, N11297, N11298, N11299, N11300, N11301, N11302, N11303, N11304, N11305, N11306, N11307, N11308, N11309, N11310, N11311, N11312, N11313, N11314, N11315, N11316, N11317, N11318, N11319, N11320, N11321, N11322, N11323, N11324, N11325, N11326, N11327, N11328, N11329, N11330, N11331, N11332, N11333, N11334, N11335, N11336, N11337, N11338, N11339, N11340, N11341, N11342, N11343, N11344, N11345, N11346, N11347, N11348, N11349, N11350, N11351, N11352, N11353, N11354, N11355, N11356, N11357, N11358, N11359, N11360, N11361, N11362, N11363, N11364, N11365, N11366, N11367, N11368, N11369, N11370, N11371, N11372, N11373, N11374, N11375, N11376, N11377, N11378, N11379, N11380, N11381, N11382, N11383, N11384, N11385, N11386, N11387, N11388, N11389, N11390, N11391, N11392, N11393, N11394, N11395, N11396, N11397, N11398, N11399, N11400, N11401, N11402, N11403, N11404, N11405, N11406, N11407, N11408, N11409, N11410, N11411, N11412, N11413, N11414, N11415, N11416, N11417, N11418, N11419, N11420, N11421, N11422, N11423, N11424, N11425, N11426, N11427, N11428, N11429, N11430, N11431, N11432, N11433, N11434, N11435, N11436, N11437, N11438, N11439, N11440, N11441, N11442, N11443, N11444, N11445, N11446, N11447, N11448, N11449, N11450, N11451, N11452, N11453, N11454, N11455, N11456, N11457, N11458, N11459, N11460, N11461, N11462, N11463, N11464, N11465, N11466, N11467, N11468, N11469, N11470, N11471, N11472, N11473, N11474, N11475, N11476, N11477, N11478, N11479, N11480, N11481, N11482, N11483, N11484, N11485, N11486, N11487, N11488, N11489, N11490, N11491, N11492, N11493, N11494, N11495, N11496, N11497, N11498, N11499, N11500, N11501, N11502, N11503, N11504, N11505, N11506, N11507, N11508, N11509, N11510, N11511, N11512, N11513, N11514, N11515, N11516, N11517, N11518, N11519, N11520, N11521, N11522, N11523, N11524, N11525, N11526, N11527, N11528, N11529, N11530, N11531, N11532, N11533, N11534, N11535, N11536, N11537, N11538, N11539, N11540, N11541, N11542, N11543, N11544, N11545, N11546, N11547, N11548, N11549, N11550, N11551, N11552, N11553, N11554, N11555, N11556, N11557, N11558, N11559, N11560, N11561, N11562, N11563, N11564, N11565, N11566, N11567, N11568, N11569, N11570, N11571, N11572, N11573, N11574, N11575, N11576, N11577, N11578, N11579, N11580, N11581, N11582, N11583, N11584, N11585, N11586, N11587, N11588, N11589, N11590, N11591, N11592, N11593, N11594, N11595, N11596, N11597, N11598, N11599, N11600, N11601, N11602, N11603, N11604, N11605, N11606, N11607, N11608, N11609, N11610, N11611, N11612, N11613, N11614, N11615, N11616, N11617, N11618, N11619, N11620, N11621, N11622, N11623, N11624, N11625, N11626, N11627, N11628, N11629, N11630, N11631, N11632, N11633, N11634, N11635, N11636, N11637, N11638, N11639, N11640, N11641, N11642, N11643, N11644, N11645, N11646, N11647, N11648, N11649, N11650, N11651, N11652, N11653, N11654, N11655, N11656, N11657, N11658, N11659, N11660, N11661, N11662, N11663, N11664, N11665, N11666, N11667, N11668, N11669, N11670, N11671, N11672, N11673, N11674, N11675, N11676, N11677, N11678, N11679, N11680, N11681, N11682, N11683, N11684, N11685, N11686, N11687, N11688, N11689, N11690, N11691, N11692, N11693, N11694, N11695, N11696, N11697, N11698, N11699, N11700, N11701, N11702, N11703, N11704, N11705, N11706, N11707, N11708, N11709, N11710, N11711, N11712, N11713, N11714, N11715, N11716, N11717, N11718, N11719, N11720, N11721, N11722, N11723, N11724, N11725, N11726, N11727, N11728, N11729, N11730, N11731, N11732, N11733, N11734, N11735, N11736, N11737, N11738, N11739, N11740, N11741, N11742, N11743, N11744, N11745, N11746, N11747, N11748, N11749, N11750, N11751, N11752, N11753, N11754, N11755, N11756, N11757, N11758, N11759, N11760, N11761, N11762, N11763, N11764, N11765, N11766, N11767, N11768, N11769, N11770, N11771, N11772, N11773, N11774, N11775, N11776, N11777, N11778, N11779, N11780, N11781, N11782, N11783, N11784, N11785, N11786, N11787, N11788, N11789, N11790, N11791, N11792, N11793, N11794, N11795, N11796, N11797, N11798, N11799, N11800, N11801, N11802, N11803, N11804, N11805, N11806, N11807, N11808, N11809, N11810, N11811, N11812, N11813, N11814, N11815, N11816, N11817, N11818, N11819, N11820, N11821, N11822, N11823, N11824, N11825, N11826, N11827, N11828, N11829, N11830, N11831, N11832, N11833, N11834, N11835, N11836, N11837, N11838, N11839, N11840, N11841, N11842, N11843, N11844, N11845, N11846, N11847, N11848, N11849, N11850, N11851, N11852, N11853, N11854, N11855, N11856, N11857, N11858, N11859, N11860, N11861, N11862, N11863, N11864, N11865, N11866, N11867, N11868, N11869, N11870, N11871, N11872, N11873, N11874, N11875, N11876, N11877, N11878, N11879, N11880, N11881, N11882, N11883, N11884, N11885, N11886, N11887, N11888, N11889, N11890, N11891, N11892, N11893, N11894, N11895, N11896, N11897, N11898, N11899, N11900, N11901, N11902, N11903, N11904, N11905, N11906, N11907, N11908, N11909, N11910, N11911, N11912, N11913, N11914, N11915, N11916, N11917, N11918, N11919, N11920, N11921, N11922, N11923, N11924, N11925, N11926, N11927, N11928, N11929, N11930, N11931, N11932, N11933, N11934, N11935, N11936, N11937, N11938, N11939, N11940, N11941, N11942, N11943, N11944, N11945, N11946, N11947, N11948, N11949, N11950, N11951, N11952, N11953, N11954, N11955, N11956, N11957, N11958, N11959, N11960, N11961, N11962, N11963, N11964, N11965, N11966, N11967, N11968, N11969, N11970, N11971, N11972, N11973, N11974, N11975, N11976, N11977, N11978, N11979, N11980, N11981, N11982, N11983, N11984, N11985, N11986, N11987, N11988, N11989, N11990, N11991, N11992, N11993, N11994, N11995, N11996, N11997, N11998, N11999, N12000, N12001, N12002, N12003, N12004, N12005, N12006, N12007, N12008, N12009, N12010, N12011, N12012, N12013, N12014, N12015, N12016, N12017, N12018, N12019, N12020, N12021, N12022, N12023, N12024, N12025, N12026, N12027, N12028, N12029, N12030, N12031, N12032, N12033, N12034, N12035, N12036, N12037, N12038, N12039, N12040, N12041, N12042, N12043, N12044, N12045, N12046, N12047, N12048, N12049, N12050, N12051, N12052, N12053, N12054, N12055, N12056, N12057, N12058, N12059, N12060, N12061, N12062, N12063, N12064, N12065, N12066, N12067, N12068, N12069, N12070, N12071, N12072, N12073, N12074, N12075, N12076, N12077, N12078, N12079, N12080, N12081, N12082, N12083, N12084, N12085, N12086, N12087, N12088, N12089, N12090, N12091, N12092, N12093, N12094, N12095, N12096, N12097, N12098, N12099, N12100, N12101, N12102, N12103, N12104, N12105, N12106, N12107, N12108, N12109, N12110, N12111, N12112, N12113, N12114, N12115, N12116, N12117, N12118, N12119, N12120, N12121, N12122, N12123, N12124, N12125, N12126, N12127, N12128, N12129, N12130, N12131, N12132, N12133, N12134, N12135, N12136, N12137, N12138, N12139, N12140, N12141, N12142, N12143, N12144, N12145, N12146, N12147, N12148, N12149, N12150, N12151, N12152, N12153, N12154, N12155, N12156, N12157, N12158, N12159, N12160, N12161, N12162, N12163, N12164, N12165, N12166, N12167, N12168, N12169, N12170, N12171, N12172, N12173, N12174, N12175, N12176, N12177, N12178, N12179, N12180, N12181, N12182, N12183, N12184, N12185, N12186, N12187, N12188, N12189, N12190, N12191, N12192, N12193, N12194, N12195, N12196, N12197, N12198, N12199, N12200, N12201, N12202, N12203, N12204, N12205, N12206, N12207, N12208, N12209, N12210, N12211, N12212, N12213, N12214, N12215, N12216, N12217, N12218, N12219, N12220, N12221, N12222, N12223, N12224, N12225, N12226, N12227, N12228, N12229, N12230, N12231, N12232, N12233, N12234, N12235, N12236, N12237, N12238, N12239, N12240, N12241, N12242, N12243, N12244, N12245, N12246, N12247, N12248, N12249, N12250, N12251, N12252, N12253, N12254, N12255, N12256, N12257, N12258, N12259, N12260, N12261, N12262, N12263, N12264, N12265, N12266, N12267, N12268, N12269, N12270, N12271, N12272, N12273, N12274, N12275, N12276, N12277, N12278, N12279, N12280, N12281, N12282, N12283, N12284, N12285, N12286, N12287, N12288, N12289, N12290, N12291, N12292, N12293, N12294, N12295, N12296, N12297, N12298, N12299, N12300, N12301, N12302, N12303, N12304, N12305, N12306, N12307, N12308, N12309, N12310, N12311, N12312, N12313, N12314, N12315, N12316, N12317, N12318, N12319, N12320, N12321, N12322, N12323, N12324, N12325, N12326, N12327, N12328, N12329, N12330, N12331, N12332, N12333, N12334, N12335, N12336, N12337, N12338, N12339, N12340, N12341, N12342, N12343, N12344, N12345, N12346, N12347, N12348, N12349, N12350, N12351, N12352, N12353, N12354, N12355, N12356, N12357, N12358, N12359, N12360, N12361, N12362, N12363, N12364, N12365, N12366, N12367, N12368, N12369, N12370, N12371, N12372, N12373, N12374, N12375, N12376, N12377, N12378, N12379, N12380, N12381, N12382, N12383, N12384, N12385, N12386, N12387, N12388, N12389, N12390, N12391, N12392, N12393, N12394, N12395, N12396, N12397, N12398, N12399, N12400, N12401, N12402, N12403, N12404, N12405, N12406, N12407, N12408, N12409, N12410, N12411, N12412, N12413, N12414, N12415, N12416, N12417, N12418, N12419, N12420, N12421, N12422, N12423, N12424, N12425, N12426, N12427, N12428, N12429, N12430, N12431, N12432, N12433, N12434, N12435, N12436, N12437, N12438, N12439, N12440, N12441, N12442, N12443, N12444, N12445, N12446, N12447, N12448, N12449, N12450, N12451, N12452, N12453, N12454, N12455, N12456, N12457, N12458, N12459, N12460, N12461, N12462, N12463, N12464, N12465, N12466, N12467, N12468, N12469, N12470, N12471, N12472, N12473, N12474, N12475, N12476, N12477, N12478, N12479, N12480, N12481, N12482, N12483, N12484, N12485, N12486, N12487, N12488, N12489, N12490, N12491, N12492, N12493, N12494, N12495, N12496, N12497, N12498, N12499, N12500, N12501, N12502, N12503, N12504, N12505, N12506, N12507, N12508, N12509, N12510, N12511, N12512, N12513, N12514, N12515, N12516, N12517, N12518, N12519, N12520, N12521, N12522, N12523, N12524, N12525, N12526, N12527, N12528, N12529, N12530, N12531, N12532, N12533, N12534, N12535, N12536, N12537, N12538, N12539, N12540, N12541, N12542, N12543, N12544, N12545, N12546, N12547, N12548, N12549, N12550, N12551, N12552, N12553, N12554, N12555, N12556, N12557, N12558, N12559, N12560, N12561, N12562, N12563, N12564, N12565, N12566, N12567, N12568, N12569, N12570, N12571, N12572, N12573, N12574, N12575, N12576, N12577, N12578, N12579, N12580, N12581, N12582, N12583, N12584, N12585, N12586, N12587, N12588, N12589, N12590, N12591, N12592, N12593, N12594, N12595, N12596, N12597, N12598, N12599, N12600, N12601, N12602, N12603, N12604, N12605, N12606, N12607, N12608, N12609, N12610, N12611, N12612, N12613, N12614, N12615, N12616, N12617, N12618, N12619, N12620, N12621, N12622, N12623, N12624, N12625, N12626, N12627, N12628, N12629, N12630, N12631, N12632, N12633, N12634, N12635, N12636, N12637, N12638, N12639, N12640, N12641, N12642, N12643, N12644, N12645, N12646, N12647, N12648, N12649, N12650, N12651, N12652, N12653, N12654, N12655, N12656, N12657, N12658, N12659, N12660, N12661, N12662, N12663, N12664, N12665, N12666, N12667, N12668, N12669, N12670, N12671, N12672, N12673, N12674, N12675, N12676, N12677, N12678, N12679, N12680, N12681, N12682, N12683, N12684, N12685, N12686, N12687, N12688, N12689, N12690, N12691, N12692, N12693, N12694, N12695, N12696, N12697, N12698, N12699, N12700, N12701, N12702, N12703, N12704, N12705, N12706, N12707, N12708, N12709, N12710, N12711, N12712, N12713, N12714, N12715, N12716, N12717, N12718, N12719, N12720, N12721, N12722, N12723, N12724, N12725, N12726, N12727, N12728, N12729, N12730, N12731, N12732, N12733, N12734, N12735, N12736, N12737, N12738, N12739, N12740, N12741, N12742, N12743, N12744, N12745, N12746, N12747, N12748, N12749, N12750, N12751, N12752, N12753, N12754, N12755, N12756, N12757, N12758, N12759, N12760, N12761, N12762, N12763, N12764, N12765, N12766, N12767, N12768, N12769, N12770, N12771, N12772, N12773, N12774, N12775, N12776, N12777, N12778, N12779, N12780, N12781, N12782, N12783, N12784, N12785, N12786, N12787, N12788, N12789, N12790, N12791, N12792, N12793, N12794, N12795, N12796, N12797, N12798, N12799, N12800, N12801, N12802, N12803, N12804, N12805, N12806, N12807, N12808, N12809, N12810, N12811, N12812, N12813, N12814, N12815, N12816, N12817, N12818, N12819, N12820, N12821, N12822, N12823, N12824, N12825, N12826, N12827, N12828, N12829, N12830, N12831, N12832, N12833, N12834, N12835, N12836, N12837, N12838, N12839, N12840, N12841, N12842, N12843, N12844, N12845, N12846, N12847, N12848, N12849, N12850, N12851, N12852, N12853, N12854, N12855, N12856, N12857, N12858, N12859, N12860, N12861, N12862, N12863, N12864, N12865, N12866, N12867, N12868, N12869, N12870, N12871, N12872, N12874, N12877, N12881, N12891, N12892, N12897, N12899, N12905, N12908, N12911, N12916, N12918, N12920, N12924, N12925, N12931, N12933, N12943, N12949, N12952, N12958, N12965, N12969, N12973, N12980, N12981, N12991, N12995, N12996, N13008, N13015, N13021, N13023, N13024, N13028, N13033, N13035, N13040, N13043, N13065, N13071, N13084, N13096, N13110, N13118, N13120, N13123, N13124, N13132, N13144, N13154, N13157, N13165, N13168, N13170, N13182, N13189, N13200, N13206, N13211, N13217, N13225, N13228, N13233, N13241, N13242, N13250, N13257, N13276, N13277, N13283, N13307, N13309, N13310, N13326, N13327, N13330, N13339, N13342, N13348, N13353, N13360, N13361, N13362, N13369, N13373, N13376, N13377, N13381, N13396, N13408, N13410, N13415, N13420, N13421, N13431, N13434, N13442, N13443, N13444, N13446, N13448, N13456, N13457, N13458, N13465, N13466, N13482, N13483, N13490, N13492, N13505, N13512, N13514, N13517, N13524, N13527, N13533, N13536, N13547, N13548, N13551, N13556, N13563, N13566, N13577, N13589, N13594, N13595, N13608, N13610, N13611, N13612, N13615, N13616, N13628, N13633, N13647, N13650, N13651, N13663, N13666, N13673, N13674, N13679, N13681, N13684, N13686, N13691, N13699, N13700, N13707, N13711, N13718, N13719, N13734, N13737, N13741, N13742, N13761, N13767, N13770, N13775, N13776, N13781, N13785, N13789, N13803, N13806, N13809, N13811, N13819, N13820, N13828, N13838, N13842, N13844, N13847, N13852, N13858, N13867, N13869, N13870, N13873, N13880, N13885, N13893, N13896, N13901, N13905, N13906, N13910, N13915, N13920, N13921, N13929, N13932, N13934, N13941, N13956, N13959, N13965, N13969, N13972, N13991, N14000, N14005, N14018, N14019, N14033, N14034, N14037, N14040, N14045, N14052, N14056, N14060, N14079, N14084, N14087, N14100, N14101, N14104, N14107, N14113, N14119, N14124, N14125, N14126, N14147, N14151, N14158, N14159, N14161, N14165, N14171, N14174, N14180, N14185, N14186, N14187, N14203, N14205, N14207, N14208, N14212, N14214, N14215, N14216, N14217, N14219, N14222, N14234, N14243, N14269, N14274, N14275, N14280, N14288, N14289, N14291, N14296, N14298, N14311, N14318, N14321, N14337, N14347, N14352, N14354, N14355, N14359, N14361, N14368, N14382, N14385, N14416, N14417, N14424, N14428, N14429, N14433, N14436, N14441, N14443, N14444, N14453, N14455, N14462, N14469, N14471, N14480, N14481, N14490, N14499, N14502, N14507, N14515, N14518, N14519, N14528, N14546, N14553, N14563, N14568, N14570, N14577, N14578, N14594, N14600, N14603, N14604, N14606, N14608, N14613, N14623, N14637, N14638, N14653, N14663, N14666, N14671, N14679, N14680, N14685, N14691, N14694, N14698, N14709, N14715, N14725, N14733, N14736, N14744, N14752, N14755, N14756, N14767, N14775, N14783, N14785, N14791, N14812, N14824, N14826, N14831, N14837, N14839, N14840, N14848, N14849, N14850, N14863, N14867, N14876, N14881, N14890, N14898, N14899, N14920, N14922, N14931, N14936, N14939, N14947, N14953, N14958, N14961, N14968, N14969, N14971, N14978, N14991, N14992, N15002, N15005, N15006, N15013, N15015, N15018, N15032, N15035, N15038, N15071, N15075, N15078, N15085, N15090, N15100, N15101, N15104, N15105, N15107, N15110, N15111, N15114, N15126, N15134, N15144, N15148, N15152, N15156, N15158, N15169, N15170, N15171, N15173, N15174, N15183, N15185, N15199, N15201, N15209, N15214, N15217, N15224, N15228, N15233, N15249, N15254, N15255, N15257, N15259, N15260, N15274, N15278, N15291, N15294, N15296, N15303, N15304, N15307, N15308, N15310, N15313, N15317, N15319, N15323, N15331, N15346, N15353, N15354, N15362, N15366, N15379, N15390, N15402, N15403, N15410, N15422, N15434, N15442, N15444, N15453, N15455, N15469, N15473, N15485, N15489, N15494, N15496, N15497, N15500, N15501, N15504, N15513, N15516, N15519, N15520, N15522, N15529, N15532, N15534, N15537, N15540, N15541, N15543, N15545, N15550, N15556, N15561, N15564, N15572, N15575, N15591, N15592, N15600, N15622, N15638, N15643, N15646, N15653, N15660, N15664, N15670, N15673, N15677, N15678, N15680, N15691, N15693, N15705, N15708, N15709, N15711, N15715, N15719, N15722, N15724, N15738, N15740, N15741, N15748, N15756, N15761, N15766, N15774, N15788, N15793, N15795, N15798, N15799, N15818, N15819, N15823, N15828, N15831, N15835, N15836, N15837, N15844, N15847, N15852, N15854, N15878, N15889, N15890, N15893, N15908, N15910, N15916, N15929, N15934, N15948, N15951, N15963, N15969, N15970, N15975, N15984, N15991, N16008, N16009, N16010, N16012, N16014, N16020, N16022, N16026, N16029, N16035, N16036, N16042, N16046, N16050, N16057, N16058, N16060, N16068, N16079, N16081, N16095, N16110, N16111, N16112, N16113, N16116, N16118, N16121, N16123, N16133, N16138, N16142, N16154, N16160, N16170, N16177, N16183, N16191, N16193, N16197, N16198, N16201, N16202, N16210, N16215, N16231, N16233, N16255, N16256, N16266, N16274, N16278, N16282, N16283, N16289, N16290, N16301, N16303, N16323, N16326, N16328, N16330, N16332, N16334, N16341, N16353, N16364, N16367, N16379, N16385, N16394, N16398, N16400, N16402, N16403, N16409, N16416, N16417, N16421, N16428, N16442, N16450, N16453, N16457, N16458, N16462, N16466, N16474, N16480, N16487, N16494, N16499, N16516, N16519, N16527, N16529, N16533, N16537, N16551, N16556, N16560, N16565, N16571, N16576, N16578, N16582, N16586, N16591, N16592, N16598, N16601, N16602, N16616, N16629, N16631, N16632, N16634, N16642, N16645, N16649, N16666, N16667, N16674, N16677, N16682, N16684, N16687, N16695, N16709, N16717, N16725, N16730, N16738, N16742, N16747, N16760, N16765, N16782, N16796, N16797, N16801, N16803, N16806, N16809, N16814, N16818, N16828, N16830, N16839, N16841, N16846, N16847, N16848, N16854, N16867, N16871, N16879, N16883, N16891, N16906, N16911, N16920, N16925, N16939, N16940, N16942, N16949, N16954, N16956, N16971, N16981, N16984, N16990, N16996, N16999, N17002, N17004, N17017, N17018, N17019, N17024, N17041, N17043, N17052, N17053, N17063, N17066, N17076, N17082, N17083, N17091, N17095, N17098, N17102, N17106, N17107, N17110, N17115, N17124, N17127, N17141, N17148, N17156, N17169, N17181, N17182, N17183, N17188, N17191, N17193, N17203, N17209, N17210, N17214, N17216, N17219, N17221, N17223, N17236, N17243, N17250, N17251, N17252, N17255, N17260, N17264, N17274, N17278, N17285, N17291, N17301, N17304, N17310, N17318, N17323, N17335, N17337, N17342, N17360, N17362, N17367, N17369, N17375, N17384, N17393, N17397, N17399, N17400, N17413, N17425, N17428, N17431, N17444, N17445, N17446, N17451, N17459, N17460, N17464, N17480, N17482, N17494, N17495, N17512, N17521, N17523, N17526, N17529, N17536, N17537, N17542, N17544, N17548, N17550, N17555, N17571, N17578, N17579, N17582, N17586, N17590, N17591, N17593, N17601, N17604, N17609, N17612, N17614, N17619, N17633, N17642, N17649, N17650, N17662, N17665, N17673, N17674, N17675, N17685, N17686, N17701, N17707, N17709, N17711, N17719, N17723, N17727, N17728, N17735, N17745, N17749, N17753, N17766, N17770, N17794, N17800, N17804, N17806, N17832, N17838, N17843, N17847, N17852, N17858, N17885, N17888, N17894, N17895, N17897, N17903, N17905, N17908, N17911, N17912, N17917, N17918, N17922, N17925, N17927, N17931, N17934, N17935, N17943, N17944, N17945, N17948, N17966, N17971, N17972, N17983, N17993, N17997, N17999, N18005, N18007, N18010, N18016, N18022, N18027, N18029, N18042, N18054, N18058, N18060, N18081, N18097, N18101, N18109, N18110, N18112, N18120, N18126, N18138, N18144, N18149, N18153, N18157, N18159, N18166, N18172, N18173, N18174, N18189, N18201, N18203, N18219, N18234, N18240, N18245, N18249, N18261, N18264, N18267, N18271, N18279, N18281, N18285, N18303, N18310, N18322, N18338, N18339, N18350, N18351, N18354, N18362, N18364, N18372, N18375, N18379, N18400, N18416, N18420, N18430, N18436, N18445, N18461, N18464, N18467, N18484, N18488, N18493, N18495, N18502, N18506, N18510, N18519, N18524, N18526, N18528, N18544, N18549, N18561, N18563, N18566, N18576, N18578, N18583, N18587, N18619, N18622, N18627, N18641, N18649, N18665, N18668, N18671, N18685, N18688, N18693, N18723, N18724, N18730, N18737, N18739, N18741, N18743, N18751, N18754, N18776, N18781, N18783, N18799, N18805, N18820, N18822, N18825, N18834, N18838, N18848, N18850, N18855, N18866, N18867, N18881, N18883, N18884, N18887, N18899, N18907, N18912, N18919, N18921, N18924, N18929, N18937, N18939, N18944, N18949, N18955, N18971, N18980, N18981, N18983, N18984, N18988, N18991, N18999, N19007, N19008, N19011, N19017, N19033, N19038, N19048, N19051, N19056, N19057, N19058, N19063, N19066, N19068, N19070, N19076, N19087, N19088, N19095, N19097, N19100, N19104, N19105, N19108, N19109, N19112, N19113, N19116, N19129, N19130, N19139, N19160, N19174, N19175, N19178, N19182, N19187, N19190, N19194, N19207, N19209, N19212, N19213, N19215, N19220, N19224, N19241, N19242, N19246, N19247, N19248, N19251, N19265, N19274, N19277, N19279, N19296, N19303, N19306, N19314, N19324, N19326, N19329, N19334, N19340, N19341, N19346, N19347, N19350, N19375, N19380, N19386, N19388, N19399, N19402, N19409, N19430, N19445, N19447, N19457, N19459, N19474, N19481, N19482, N19484, N19493, N19499, N19524, N19527, N19531, N19532, N19534, N19536, N19537, N19543, N19549, N19561, N19564, N19567, N19568, N19570, N19577, N19583, N19585, N19593, N19596, N19617, N19622, N19623, N19630, N19633, N19657, N19658, N19668, N19670, N19673, N19676, N19678, N19686, N19693, N19696, N19714, N19729, N19743, N19744, N19746, N19747, N19748, N19751, N19763, N19780, N19785, N19816, N19819, N19822, N19823, N19824, N19829, N19832, N19839, N19844, N19851, N19852, N19859, N19864, N19870, N19871, N19872, N19881, N19892, N19893, N19897, N19905, N19909, N19918, N19920, N19921, N19927, N19937, N19938, N19939, N19942, N19948, N19951, N19953, N19960, N19968, N19969, N19978, N19986, N19988, N19995, N19998, N20002, N20003, N20007, N20010, N20018, N20019, N20036, N20042, N20047, N20048, N20055, N20057, N20059, N20060, N20066, N20068, N20069, N20072, N20074, N20077, N20082, N20087, N20089, N20099, N20105, N20108, N20119, N20123, N20125, N20135, N20138, N20146, N20154, N20158, N20164, N20186, N20189, N20190, N20191, N20192, N20197, N20199, N20203, N20208, N20217, N20218, N20227, N20249, N20270, N20277, N20278, N20279, N20281, N20284, N20286, N20287, N20291, N20292, N20295, N20299, N20300, N20309, N20314, N20333, N20345, N20354, N20359, N20360, N20367, N20369, N20376, N20394, N20396, N20403, N20404, N20407, N20408, N20409, N20411, N20413, N20422, N20425, N20429, N20445, N20455, N20458, N20479, N20484, N20493, N20495, N20507, N20508, N20515, N20522, N20523, N20533, N20534, N20536, N20541, N20545, N20547, N20567, N20576, N20577, N20586, N20588, N20594, N20598, N20601, N20602, N20604, N20606, N20607, N20610, N20613, N20618, N20619, N20629, N20637, N20638, N20640, N20650, N20652, N20653, N20661, N20663, N20668, N20680, N20685, N20692, N20703, N20710, N20727, N20744, N20747, N20748, N20771, N20773, N20776, N20783, N20787, N20791, N20799, N20803, N20806, N20807, N20808, N20816, N20818, N20823, N20824, N20843, N20851, N20863, N20864, N20870, N20873, N20874, N20888, N20893, N20900, N20902, N20906, N20911, N20916, N20921, N20924, N20933, N20935, N20938, N20941, N20952, N20958, N20963, N20970, N20971, N21001, N21019, N21022, N21023, N21024, N21036, N21037, N21038, N21041, N21050, N21051, N21064, N21065, N21074, N21085, N21086, N21094, N21095, N21096, N21106, N21115, N21116, N21119, N21122, N21134, N21140, N21145, N21150, N21157, N21161, N21170, N21191, N21192, N21203, N21206, N21211, N21213, N21214, N21217, N21219, N21226, N21227, N21228, N21231, N21235, N21238, N21241, N21248, N21251, N21252, N21254, N21257, N21261, N21264, N21270, N21274, N21276, N21284, N21285, N21287, N21291, N21292, N21296, N21302, N21304, N21306, N21307, N21316, N21323, N21325, N21327, N21330, N21331, N21332, N21333, N21334, N21336, N21349, N21350, N21352, N21354, N21356, N21357, N21362, N21368, N21371, N21372, N21377, N21382, N21386, N21388, N21395, N21397, N21399, N21402, N21404, N21406, N21416, N21421, N21426, N21432, N21433, N21438, N21445, N21450, N21452, N21457, N21459, N21465, N21466, N21467, N21468, N21469, N21470, N21481, N21483, N21485, N21491, N21498, N21503, N21509, N21516, N21518, N21521, N21523, N21527, N21530, N21537, N21538, N21540, N21546, N21547, N21555, N21561, N21562, N21566, N21567, N21569, N21571, N21582, N21584, N21585, N21586, N21590, N21591, N21597, N21598, N21607, N21609, N21610, N21611, N21613, N21617, N21622, N21624, N21629, N21631, N21636, N21637, N21641, N21654, N21669, N21672, N21675, N21684, N21685, N21686, N21687, N21688, N21692, N21694, N21698, N21705, N21712, N21715, N21717, N21719, N21721, N21727, N21739, N21741, N21742, N21745, N21746, N21753, N21758, N21769, N21770, N21772, N21773, N21781, N21786, N21788, N21795, N21796, N21797, N21798, N21813, N21833, N21835, N21842, N21852, N21857, N21860, N21862, N21864, N21868, N21869, N21871, N21876, N21882, N21885, N21889, N21891, N21898, N21902, N21908, N21909, N21914, N21916, N21918, N21930, N21935, N21943, N21954, N21957, N21958, N21959, N21964, N21966, N21971, N21978, N21982, N21983, N21987, N21989, N21991, N21994, N21995, N21996, N21998, N21999, N22003, N22008, N22014, N22018, N22019, N22023, N22024, N22026, N22029, N22032, N22037, N22040, N22043, N22049, N22052, N22053, N22058, N22059, N22060, N22064, N22066, N22067, N22068, N22069, N22070, N22071, N22073, N22076, N22077, N22080, N22081, N22084, N22100, N22102, N22104, N22105, N22116, N22117, N22121, N22123, N22126, N22132, N22140, N22142, N22145, N22147, N22150, N22157, N22161, N22167, N22173, N22177, N22183, N22185, N22186, N22188, N22191, N22197, N22199, N22204, N22206, N22213, N22215, N22217, N22218, N22221, N22222, N22223, N22225, N22234, N22235, N22237, N22240, N22241, N22243, N22244, N22248, N22249, N22251, N22257, N22262, N22263, N22266, N22272, N22284, N22287, N22302, N22303, N22307, N22311, N22312, N22315, N22317, N22324, N22327, N22329, N22330, N22332, N22334, N22340, N22341, N22342, N22343, N22344, N22350, N22354, N22363, N22365, N22368, N22372, N22377, N22380, N22382, N22391, N22397, N22398, N22400, N22401, N22420, N22424, N22430, N22432, N22435, N22439, N22440, N22446, N22454, N22460, N22467, N22470, N22472, N22473, N22488, N22489, N22490, N22495, N22498, N22503, N22510, N22511, N22512, N22516, N22517, N22520, N22521, N22523, N22528, N22537, N22541, N22547, N22549, N22551, N22552, N22560, N22561, N22563, N22568, N22578, N22589, N22595, N22597, N22606, N22618, N22621, N22622, N22629, N22631, N22634, N22638, N22648, N22650, N22656, N22659, N22664, N22676, N22677, N22682, N22683, N22684, N22693, N22694, N22699, N22704, N22705, N22706, N22709, N22714, N22715, N22724, N22727, N22730, N22737, N22749, N22761, N22764, N22769, N22779, N22780, N22782, N22783, N22790, N22792, N22794, N22797, N22804, N22806, N22809, N22810, N22818, N22819, N22821, N22822, N22823, N22824, N22827, N22829, N22831, N22834, N22840, N22842, N22846, N22850, N22860, N22861, N22873, N22876, N22880, N22884, N22888, N22893, N22895, N22900, N22901, N22902, N22911, N22914, N22916, N22918, N22920, N22922, N22934, N22941, N22942, N22947, N22951, N22955, N22959, N22968, N22978, N22980, N22984, N22991, N22994, N22997, N22998, N23000, N23001, N23007, N23008, N23009, N23018, N23019, N23026, N23028, N23029, N23032, N23038, N23054, N23056, N23057, N23058, N23059, N23064, N23068, N23072, N23076, N23081, N23086, N23087, N23090, N23092, N23093, N23101, N23102, N23110, N23111, N23112, N23114, N23116, N23117, N23121, N23126, N23129, N23133, N23135, N23137, N23141, N23142, N23147, N23148, N23157, N23159, N23165, N23170, N23178, N23186, N23188, N23194, N23196, N23197, N23198, N23199, N23201, N23214, N23217, N23218, N23221, N23222, N23223, N23224, N23225, N23228, N23231, N23232, N23241, N23244, N23245, N23246, N23247, N23251, N23259, N23261, N23262, N23269, N23277, N23280, N23283, N23287, N23289, N23297, N23300, N23312, N23315, N23316, N23320, N23324, N23331, N23336, N23349, N23351, N23359, N23365, N23366, N23367, N23369, N23370, N23374, N23376, N23378, N23390, N23391, N23392, N23395, N23397, N23406, N23413, N23415, N23420, N23433, N23439, N23447, N23455, N23456, N23457, N23458, N23459, N23468, N23475, N23478, N23481, N23482, N23486, N23489, N23492, N23493, N23494, N23506, N23508, N23515, N23517, N23521, N23522, N23528, N23535, N23537, N23540, N23547, N23554, N23558, N23559, N23560, N23563, N23567, N23575, N23579, N23587, N23588, N23590, N23592, N23594, N23597, N23600, N23602, N23607, N23610, N23611, N23613, N23622, N23630, N23634, N23636, N23641, N23646, N23655, N23656, N23660, N23661, N23667, N23671, N23675, N23680, N23685, N23693, N23699, N23700, N23701, N23702, N23705, N23708, N23712, N23732, N23738, N23739, N23746, N23749, N23755, N23758, N23759, N23760, N23769, N23770, N23771, N23772, N23774, N23778, N23783, N23791, N23795, N23800, N23803, N23805, N23815, N23817, N23819, N23824, N23830, N23831, N23832, N23843, N23844, N23845, N23846, N23847, N23848, N23852, N23853, N23858, N23861, N23869, N23870, N23872, N23874, N23878, N23889, N23891, N23894, N23896, N23897, N23905, N23908, N23922, N23925, N23926, N23942, N23944, N23947, N23951, N23954, N23963, N23967, N23975, N23978, N23981, N23983, N23988, N23991, N23994, N24010, N24023, N24024, N24027, N24028, N24033, N24041, N24043, N24047, N24052, N24053, N24061, N24062, N24065, N24066, N24068, N24069, N24079, N24080, N24081, N24084, N24092, N24097, N24098, N24104, N24115, N24117, N24130, N24131, N24133, N24134, N24137, N24138, N24139, N24140, N24143, N24144, N24151, N24153, N24161, N24162, N24164, N24168, N24172, N24173, N24178, N24188, N24192, N24196, N24214, N24221, N24222, N24230, N24234, N24238, N24241, N24244, N24246, N24249, N24254, N24259, N24266, N24273, N24274, N24277, N24279, N24283, N24286, N24290, N24295, N24297, N24298, N24299, N24302, N24305, N24309, N24312, N24314, N24315, N24325, N24327, N24342, N24347, N24352, N24360, N24362, N24372, N24374, N24380, N24381, N24393, N24399, N24403, N24404, N24407, N24420, N24426, N24436, N24440, N24443, N24445, N24446, N24454, N24457, N24466, N24468, N24472, N24483, N24486, N24489, N24493, N24506, N24512, N24515, N24516, N24519, N24527, N24530, N24531, N24534, N24535, N24539, N24544, N24552, N24555, N24557, N24574, N24578, N24582, N24584, N24590, N24592, N24593, N24598, N24599, N24603, N24607, N24609, N24613, N24615, N24619, N24621, N24622, N24624, N24628, N24633, N24638, N24642, N24644, N24646, N24647, N24650, N24651, N24657, N24663, N24675, N24696, N24706, N24711, N24715, N24717, N24724, N24732, N24736, N24739, N24742, N24747, N24749, N24752, N24757, N24761, N24775, N24776, N24777, N24782, N24783, N24784, N24785, N24807, N24813, N24814, N24815, N24823, N24824, N24826, N24829, N24830, N24832, N24840, N24844, N24847, N24848, N24855, N24856, N24858, N24859, N24864, N24869, N24870, N24871, N24872, N24877, N24884, N24885, N24887, N24890, N24894, N24895, N24896, N24903, N24917, N24922, N24927, N24929, N24933, N24937, N24938, N24939, N24941, N24943, N24945, N24946, N24950, N24954, N24956, N24964, N24968, N24969, N24973, N24975, N24978, N24979, N24983, N24990, N24992, N25003, N25006, N25012, N25016, N25017, N25021, N25033, N25042, N25045, N25054, N25057, N25062, N25064, N25066, N25067, N25069, N25079, N25080, N25088, N25091, N25092, N25113, N25114, N25115, N25118, N25120, N25121, N25122, N25123, N25132, N25135, N25136, N25143, N25144, N25157, N25158, N25165, N25170, N25171, N25172, N25179, N25181, N25186, N25190, N25192, N25193, N25199, N25200, N25207, N25210, N25229, N25233, N25235, N25237, N25238, N25239, N25240, N25247, N25256, N25257, N25260, N25265, N25266, N25267, N25268, N25272, N25278, N25281, N25282, N25285, N25288, N25295, N25296, N25309, N25310, N25313, N25316, N25318, N25319, N25324, N25330, N25337, N25339, N25340, N25345, N25347, N25350, N25356, N25358, N25359, N25368, N25373, N25375, N25376, N25380, N25381, N25390, N25396, N25397, N25399, N25400, N25401, N25407, N25412, N25420, N25425, N25426, N25429, N25430, N25431, N25434, N25437, N25439, N25443, N25448, N25451, N25452, N25456, N25458, N25461, N25464, N25468, N25470, N25472, N25473, N25480, N25483, N25489, N25491, N25500, N25501, N25505, N25506, N25512, N25514, N25520, N25521, N25523, N25527, N25530, N25535, N25538, N25540, N25541, N25542, N25543, N25545, N25549, N25552, N25554, N25556, N25558, N25559, N25560, N25575, N25576, N25577, N25578, N25585, N25587, N25589, N25595, N25596, N25599, N25606, N25609, N25610, N25611, N25612, N25616, N25617, N25618, N25620, N25622, N25623, N25628, N25629, N25634, N25637, N25643, N25645, N25646, N25647, N25648, N25652, N25655, N25659, N25666, N25667, N25670, N25673, N25674, N25675, N25678, N25682, N25684, N25686, N25687, N25688, N25690, N25695, N25705, N25709, N25711, N25713, N25714, N25715, N25722, N25724, N25726, N25727, N25729, N25733, N25735, N25736, N25737, N25739, N25740, N25742, N25744, N25746, N25749, N25752, N25755, N25757, N25761, N25762, N25763, N25767, N25769, N25770, N25772, N25779, N25780, N25781, N25791, N25793, N25797, N25798, N25807, N25809, N25811, N25812, N25818, N25828, N25835, N25838, N25840, N25843, N25848, N25851, N25853, N25854, N25855, N25859, N25861, N25867, N25870, N25888, N25892, N25896, N25907, N25908, N25910, N25913, N25914, N25918, N25923, N25928, N25935, N25936, N25944, N25946, N25948, N25958, N25959, N25960, N25968, N25970, N25971, N25972, N25976, N25978, N25988, N26000, N26002, N26005, N26006, N26009, N26010, N26020, N26023, N26024, N26028, N26029, N26032, N26034, N26039, N26042, N26048, N26050, N26052, N26053, N26055, N26056, N26058, N26062, N26065, N26072, N26073, N26076, N26077, N26078, N26079, N26080, N26091, N26094, N26096, N26097, N26100, N26103, N26104, N26106, N26112, N26113, N26116, N26118, N26120, N26123, N26124, N26131, N26132, N26134, N26137, N26138, N26139, N26141, N26146, N26152, N26153, N26154, N26161, N26162, N26163, N26166, N26170, N26171, N26181, N26183, N26188, N26189, N26191, N26192, N26197, N26199, N26200, N26201, N26204, N26206, N26208, N26214, N26215, N26219, N26221, N26223, N26227, N26228, N26230, N26231, N26234, N26235, N26236, N26237, N26238, N26244, N26246, N26247, N26249, N26251, N26254, N26259, N26261, N26264, N26273, N26274, N26276, N26277, N26279, N26284, N26285, N26286, N26288, N26289, N26298, N26304, N26317, N26322, N26326, N26329, N26337, N26339, N26346, N26347, N26349, N26351, N26353, N26354, N26358, N26359, N26361, N26363, N26365, N26367, N26369, N26372, N26374, N26375, N26378, N26384, N26385, N26386, N26387, N26397, N26399, N26400, N26402, N26403, N26406, N26408, N26409, N26410, N26413, N26429, N26432, N26434, N26435, N26436, N26440, N26442, N26446, N26452, N26453, N26454, N26461, N26467, N26470, N26475, N26477, N26478, N26480, N26483, N26490, N26492, N26494, N26496, N26499, N26500, N26503, N26505, N26514, N26515, N26518, N26521, N26522, N26523, N26524, N26528, N26529, N26531, N26534, N26535, N26537, N26540, N26541, N26551, N26553, N26558, N26562, N26563, N26570, N26571, N26573, N26574, N26575, N26577, N26592, N26593, N26594, N26603, N26609, N26611, N26620, N26625, N26629, N26630, N26631, N26637, N26640, N26644, N26649, N26656, N26659, N26660, N26662, N26668, N26672, N26681, N26692, N26698, N26699, N26701, N26702, N26705, N26706, N26710, N26712, N26714, N26717, N26718, N26721, N26726, N26728, N26736, N26739, N26741, N26743, N26745, N26747, N26757, N26760, N26765, N26766, N26771, N26776, N26777, N26781, N26784, N26785, N26787, N26789, N26790, N26794, N26798, N26799, N26800, N26803, N26809, N26816, N26820, N26821, N26822, N26823, N26825, N26828, N26830, N26832, N26837, N26844, N26845, N26851, N26854, N26855, N26857, N26864, N26865, N26880, N26885, N26886, N26895, N26896, N26899, N26903, N26904, N26905, N26907, N26909, N26912, N26913, N26921, N26923, N26924, N26930, N26931, N26939, N26940, N26942, N26945, N26950, N26954, N26955, N26957, N26961, N26964, N26971, N26973, N26984, N26986, N26987, N26988, N26989, N26991, N26992, N26993, N26997, N26999, N27001, N27002, N27004, N27010, N27013, N27014, N27016, N27021, N27023, N27024, N27025, N27027, N27034, N27035, N27036, N27038, N27040, N27041, N27042, N27045, N27046, N27047, N27048, N27058, N27061, N27063, N27065, N27071, N27073, N27074, N27075, N27078, N27079, N27088, N27090, N27091, N27094, N27106, N27114, N27118, N27120, N27128, N27129, N27130, N27133, N27134, N27135, N27136, N27142, N27148, N27150, N27158, N27159, N27166, N27169, N27172, N27180, N27187, N27188, N27189, N27192, N27193, N27194, N27195, N27198, N27200, N27202, N27203, N27204, N27208, N27212, N27216, N27222, N27224, N27227, N27228, N27230, N27233, N27238, N27242, N27243, N27244, N27246, N27248, N27251, N27253, N27254, N27258, N27263, N27273, N27277, N27284, N27292, N27295, N27299, N27302, N27306, N27307, N27311, N27312, N27313, N27315, N27322, N27323, N27326, N27330, N27333, N27335, N27338, N27341, N27343, N27344, N27345, N27348, N27350, N27351, N27352, N27356, N27359, N27363, N27364, N27367, N27371, N27372, N27375, N27381, N27383, N27385, N27386, N27388, N27390, N27395, N27398, N27400, N27409, N27410, N27414, N27415, N27418, N27424, N27430, N27432, N27435, N27437, N27441, N27443, N27446, N27447, N27450, N27451, N27457, N27458, N27460, N27461, N27466, N27468, N27469, N27470, N27471, N27475, N27476, N27481, N27485, N27487, N27490, N27491, N27493, N27494, N27495, N27497, N27502, N27504, N27505, N27529, N27530, N27531, N27539, N27542, N27548, N27550, N27551, N27555, N27559, N27563, N27568, N27569, N27570, N27576, N27579, N27580, N27586, N27587, N27590, N27591, N27603, N27611, N27612, N27613, N27614, N27618, N27622, N27626, N27627, N27628, N27629, N27630, N27632, N27633, N27635, N27636, N27646, N27647, N27648, N27649, N27650, N27653, N27654, N27655, N27660, N27662, N27664, N27665, N27671, N27672, N27675, N27676, N27681, N27682, N27685, N27686, N27689, N27693, N27699, N27701, N27704, N27708, N27711, N27713, N27716, N27719, N27720, N27721, N27722, N27728, N27729, N27731, N27733, N27735, N27738, N27744, N27748, N27751, N27752, N27756, N27757, N27762, N27764, N27769, N27770, N27775, N27778, N27780, N27783, N27786, N27787, N27788, N27789, N27790, N27792, N27794, N27798, N27804, N27805, N27807, N27809, N27811, N27813, N27818, N27828, N27829, N27830, N27833, N27835, N27837, N27841, N27842, N27844, N27848, N27849, N27850, N27854, N27856, N27861, N27868, N27873, N27879, N27883, N27886, N27887, N27890, N27894, N27896, N27900, N27903, N27906, N27907, N27915, N27918, N27922, N27931, N27932, N27935, N27941, N27942, N27944, N27947, N27949, N27954, N27955, N27958, N27959, N27965, N27967, N27974, N27976, N27977, N27984, N27986, N27988, N27990, N27994, N28000, N28001, N28003, N28005, N28007, N28012, N28026, N28030, N28032, N28033, N28035, N28038, N28039, N28040, N28048, N28051, N28054, N28059, N28062, N28065, N28067, N28068, N28071, N28073, N28074, N28075, N28080, N28084, N28085, N28099, N28100, N28108, N28117, N28119, N28120, N28123, N28128, N28129, N28130, N28131, N28134, N28140, N28145, N28149, N28152, N28153, N28155, N28157, N28166, N28167, N28168, N28173, N28175, N28180, N28181, N28184, N28187, N28188, N28189, N28196, N28200, N28207, N28209, N28210, N28212, N28213, N28216, N28221, N28223, N28224, N28225, N28228, N28230, N28231, N28236, N28239, N28240, N28243, N28247, N28249, N28251, N28255, N28259, N28261, N28262, N28263, N28266, N28268, N28274, N28275, N28278, N28280, N28281, N28283, N28285, N28286, N28288, N28291, N28292, N28293, N28296, N28300, N28306, N28315, N28316, N28319, N28322, N28323, N28327, N28330, N28331, N28332, N28333, N28337, N28338, N28340, N28341, N28343, N28351, N28355, N28357, N28360, N28362, N28366, N28367, N28369, N28370, N28373, N28376, N28377, N28378, N28383, N28388, N28391, N28394, N28395, N28398, N28400, N28402, N28407, N28413, N28414, N28415, N28416, N28420, N28424, N28425, N28428, N28433, N28438, N28442, N28447, N28449, N28453, N28454, N28462, N28464, N28468, N28470, N28473, N28474, N28480, N28482, N28484, N28489, N28492, N28502, N28504, N28505, N28509, N28517, N28518, N28519, N28524, N28525, N28527, N28530, N28533, N28534, N28535, N28536, N28539, N28541, N28542, N28543, N28549, N28550, N28552, N28558, N28562, N28563, N28573, N28576, N28579, N28580, N28583, N28584, N28591, N28592, N28593, N28595, N28597, N28598, N28604, N28605, N28607, N28608, N28609, N28612, N28613, N28621, N28623, N28624, N28626, N28632, N28638, N28641, N28647, N28648, N28658, N28661, N28666, N28670, N28671, N28672, N28676, N28683, N28694, N28696, N28700, N28707, N28713, N28715, N28722, N28723, N28725, N28728, N28733, N28734, N28735, N28736, N28745, N28748, N28751, N28752, N28755, N28759, N28765, N28775, N28778, N28780, N28784, N28790, N28791, N28792, N28799, N28800, N28802, N28806, N28811, N28812, N28814, N28816, N28818, N28824, N28826, N28827, N28829, N28830, N28834, N28835, N28849, N28851, N28852, N28853, N28858, N28862, N28863, N28866, N28869, N28872, N28875, N28879, N28881, N28883, N28887, N28890, N28898, N28899, N28900, N28902, N28903, N28917, N28918, N28924, N28926, N28928, N28929, N28931, N28932, N28934, N28935, N28936, N28940, N28941, N28947, N28955, N28961, N28967, N28971, N28972, N28976, N28985, N28992, N28994, N29001, N29002, N29003, N29017, N29020, N29023, N29029, N29034, N29042, N29045, N29053, N29054, N29056, N29057, N29059, N29060, N29062, N29067, N29068, N29070, N29073, N29074, N29076, N29077, N29080, N29081, N29086, N29092, N29095, N29096, N29103, N29111, N29112, N29115, N29121, N29123, N29124, N29126, N29127, N29128, N29137, N29138, N29140, N29141, N29142, N29143, N29145, N29152, N29155, N29161, N29166, N29171, N29177, N29178, N29184, N29187, N29189, N29192, N29194, N29199, N29200, N29202, N29203, N29204, N29206, N29209, N29213, N29215, N29218, N29220, N29224, N29229, N29234, N29237, N29252, N29256, N29258, N29261, N29267, N29268, N29269, N29273, N29277, N29283, N29288, N29290, N29291, N29297, N29301, N29302, N29303, N29306, N29307, N29312, N29328, N29334, N29336, N29338, N29341, N29342, N29345, N29348, N29349, N29350, N29356, N29357, N29360, N29361, N29362, N29368, N29369, N29370, N29373, N29378, N29379, N29380, N29381, N29387, N29390, N29395, N29396, N29404, N29411, N29414, N29415, N29417, N29421, N29426, N29427, N29429, N29439, N29447, N29448, N29452, N29461, N29462, N29466, N29469, N29471, N29473, N29476, N29478, N29482, N29488, N29493, N29497, N29498, N29499, N29501, N29507, N29520, N29527, N29529, N29530, N29533, N29534, N29537, N29538, N29539, N29543, N29549, N29550, N29552, N29554, N29558, N29562, N29563, N29568, N29570, N29571, N29572, N29573, N29576, N29579, N29581, N29584, N29585, N29588, N29590, N29594, N29601, N29605, N29606, N29610, N29614, N29620, N29624, N29627, N29628, N29631, N29632, N29633, N29640, N29641, N29643, N29645, N29646, N29648, N29649, N29651, N29652, N29654, N29655, N29657, N29658, N29659, N29662, N29663, N29666, N29668, N29669, N29670, N29676, N29679, N29682, N29686, N29690, N29691, N29693, N29699, N29700, N29703, N29711, N29712, N29713, N29724, N29726, N29727, N29729, N29731, N29734, N29742, N29746, N29747, N29748, N29750, N29751, N29760, N29764, N29765, N29767, N29768, N29779, N29785, N29786, N29787, N29789, N29794, N29795, N29796, N29798, N29802, N29804, N29808, N29811, N29812, N29813, N29816, N29817, N29820, N29822, N29825, N29829, N29833, N29836, N29837, N29840, N29843, N29845, N29846, N29849, N29850, N29852, N29853, N29855, N29857, N29863, N29866, N29873, N29874, N29875, N29876, N29878, N29879, N29885, N29886, N29894, N29899, N29901, N29907, N29913, N29918, N29923, N29925, N29926, N29927, N29928, N29931, N29934, N29935, N29942, N29944, N29946, N29947, N29948, N29952, N29953, N29955, N29956, N29957, N29959, N29960, N29965, N29966, N29969, N29972, N29975, N29976, N29980, N29981, N29984, N29987, N29988, N30007, N30008, N30009, N30012, N30015, N30027, N30031, N30034, N30035, N30036, N30042, N30044, N30045, N30046, N30050, N30057, N30059, N30060, N30064, N30066, N30070, N30077, N30079, N30080, N30084, N30085, N30091, N30093, N30096, N30097, N30098, N30102, N30104, N30105, N30108, N30109, N30110, N30111, N30116, N30118, N30119, N30123, N30124, N30127, N30135, N30137, N30138, N30139, N30140, N30141, N30142, N30143, N30144, N30146, N30148, N30149, N30150, N30155, N30157, N30158, N30161, N30162, N30163, N30164, N30165, N30169, N30170, N30171, N30174, N30176, N30177, N30178, N30179, N30180, N30181, N30183, N30184, N30186, N30187, N30188, N30189, N30190, N30191, N30192, N30193, N30194, N30195, N30196, N30197, N30198, N30199, N30201, N30203, N30205, N30206, N30208, N30210, N30212, N30213, N30214, N30215, N30216, N30217, N30218, N30219, N30221, N30222, N30223, N30224, N30225, N30226, N30227, N30228, N30230, N30233, N30236, N30237, N30239, N30241, N30242, N30243, N30245, N30247, N30248, N30249, N30252, N30253, N30255, N30256, N30258, N30259, N30260, N30262, N30263, N30264, N30265, N30266, N30267, N30268, N30270, N30272, N30273, N30275, N30278, N30279, N30280, N30281, N30283, N30284, N30286, N30288, N30292, N30293, N30295, N30296, N30297, N30298, N30301, N30303, N30305, N30307, N30309, N30313, N30314, N30316, N30317, N30319, N30321, N30322, N30323, N30325, N30326, N30330, N30331, N30333, N30334, N30336, N30337, N30338, N30339, N30341, N30343, N30344, N30345, N30347, N30348, N30350, N30352, N30354, N30357, N30358, N30359, N30361, N30363, N30364, N30365, N30366, N30367, N30369, N30370, N30372, N30373, N30374, N30375, N30376, N30377, N30378, N30381, N30382, N30383, N30386, N30389, N30391, N30393, N30395, N30396, N30398, N30401, N30404, N30405, N30406, N30407, N30411, N30412, N30413, N30414, N30415, N30416, N30418, N30419, N30420, N30421, N30424, N30426, N30427, N30428, N30432, N30434, N30435, N30437, N30438, N30440, N30442, N30443, N30444, N30446, N30447, N30448, N30449, N30452, N30453, N30454, N30455, N30456, N30457, N30458, N30459, N30460, N30461, N30462, N30463, N30466, N30467, N30468, N30469, N30470, N30471, N30474, N30476, N30477, N30479, N30480, N30481, N30484, N30485, N30487, N30488, N30491, N30493, N30495, N30496, N30497, N30498, N30499, N30500, N30502, N30503, N30504, N30505, N30506, N30507, N30508, N30509, N30510, N30514, N30515, N30517, N30519, N30520, N30521, N30522, N30523, N30524, N30527, N30528, N30529, N30530, N30531, N30532, N30533, N30534, N30536, N30537, N30539, N30540, N30544, N30545, N30546, N30551, N30553, N30554, N30557, N30559, N30560, N30561, N30564, N30572, N30575, N30577, N30578, N30579, N30580, N30582, N30584, N30585, N30586, N30588, N30589, N30590, N30591, N30592, N30593, N30595, N30596, N30597, N30598, N30601, N30602, N30603, N30605, N30608, N30609, N30611, N30612, N30613, N30615, N30616, N30617, N30618, N30620, N30621, N30622, N30623, N30625, N30627, N30628, N30631, N30633, N30634, N30635, N30636, N30638, N30639, N30641, N30642, N30643, N30644, N30649, N30650, N30651, N30652, N30654, N30655, N30656, N30658, N30659, N30660, N30662, N30663, N30664, N30665, N30666, N30667, N30668, N30669, N30670, N30671, N30672, N30673, N30674, N30675, N30676, N30677, N30678, N30679, N30681, N30682, N30683, N30685, N30687, N30688, N30689, N30691, N30692, N30693, N30694, N30696, N30699, N30703, N30704, N30705, N30706, N30710, N30712, N30713, N30714, N30716, N30717, N30718, N30719, N30721, N30724, N30725, N30726, N30727, N30730, N30731, N30732, N30735, N30737, N30739, N30741, N30742, N30743, N30744, N30747, N30749, N30750, N30751, N30753, N30755, N30756, N30758, N30759, N30761, N30763, N30766, N30767, N30768, N30769, N30772, N30773, N30774, N30777, N30779, N30780, N30781, N30782, N30784, N30785, N30786, N30787, N30789, N30790, N30791, N30792, N30793, N30794, N30795, N30796, N30801, N30803, N30804, N30806, N30808, N30809, N30810, N30813, N30815, N30816, N30817, N30818, N30819, N30822, N30823, N30824, N30826, N30827, N30828, N30829, N30832, N30833, N30834, N30836, N30837, N30838, N30839, N30840, N30842, N30843, N30845, N30846, N30847, N30849, N30850, N30851, N30852, N30853, N30855, N30856, N30858, N30861, N30862, N30863, N30864, N30865, N30866, N30869, N30871, N30872, N30873, N30875, N30876, N30877, N30879, N30880, N30881, N30882, N30883, N30885, N30886, N30887, N30888, N30890, N30893, N30895, N30896, N30898, N30900, N30901, N30902, N30903, N30904, N30905, N30907, N30908, N30912, N30913, N30914, N30915, N30916, N30917, N30918, N30919, N30921, N30922, N30923, N30925, N30926, N30930, N30933, N30934, N30935, N30936, N30937, N30939, N30942, N30944, N30945, N30946, N30947, N30948, N30949, N30950, N30952, N30953, N30957, N30959, N30960, N30962, N30963, N30964, N30965, N30966, N30968, N30970, N30971, N30972, N30974, N30975, N30976, N30977, N30979, N30981, N30982, N30983, N30986, N30987, N30988, N30991, N30992, N30993, N30994, N30998, N30999, N31000, N31003, N31004, N31005, N31006, N31007, N31009, N31010, N31016, N31017, N31018, N31019, N31020, N31021, N31022, N31023, N31028, N31029, N31032, N31033, N31035, N31036, N31037, N31038, N31039, N31041, N31043, N31045, N31047, N31048, N31050, N31051, N31052, N31053, N31054, N31056, N31057, N31058, N31059, N31061, N31062, N31064, N31065, N31068, N31069, N31071, N31072, N31077, N31078, N31080, N31081, N31082, N31083, N31085, N31088, N31089, N31093, N31094, N31096, N31097, N31098, N31101, N31103, N31105, N31107, N31108, N31110, N31111, N31112, N31113, N31115, N31116, N31117, N31118, N31123, N31125, N31127, N31128, N31129, N31131, N31133, N31134, N31137, N31138, N31141, N31145, N31148, N31149, N31152, N31153, N31155, N31157, N31158, N31159, N31160, N31163, N31164, N31165, N31166, N31167, N31169, N31171, N31172, N31174, N31176, N31178, N31180, N31182, N31184, N31185, N31186, N31188, N31189, N31192, N31193, N31194, N31196, N31197, N31199, N31200, N31202, N31203, N31204, N31205, N31206, N31207, N31210, N31211, N31212, N31213, N31218, N31219, N31220, N31221, N31223, N31224, N31225, N31227, N31229, N31230, N31231, N31232, N31233, N31235, N31236, N31240, N31241, N31243, N31246, N31248, N31251, N31252, N31253, N31255, N31258, N31259, N31260, N31262, N31263, N31266, N31269, N31270, N31271, N31272, N31273, N31274, N31275, N31277, N31280, N31282, N31283, N31284, N31285, N31286, N31287, N31290, N31291, N31293, N31294, N31295, N31297, N31299, N31301, N31308, N31309, N31310, N31312, N31313, N31315, N31317, N31319, N31320, N31321, N31324, N31325, N31326, N31328, N31329, N31332, N31333, N31335, N31336, N31337, N31338, N31339, N31340, N31341, N31342, N31343, N31346, N31350, N31352, N31355, N31356, N31357, N31361, N31362, N31364, N31365, N31367, N31368, N31370, N31371, N31372, N31374, N31375, N31376, N31377, N31378, N31379, N31382, N31383, N31385, N31386, N31387, N31388, N31389, N31390, N31391, N31392, N31393, N31395, N31396, N31397, N31398, N31401, N31402, N31403, N31404, N31405, N31406, N31407, N31408, N31409, N31412, N31414, N31415, N31416, N31417, N31418, N31420, N31421, N31422, N31424, N31425, N31428, N31430, N31431, N31432, N31433, N31434, N31438, N31439, N31441, N31443, N31447, N31448, N31450, N31451, N31452, N31453, N31459, N31463, N31464, N31465, N31466, N31467, N31469, N31471, N31472, N31473, N31474, N31475, N31477, N31478, N31479, N31481, N31482, N31483, N31484, N31485, N31488, N31489, N31490, N31491, N31492, N31495, N31496, N31497, N31498, N31499, N31501, N31502, N31505, N31506, N31507, N31508, N31511, N31512, N31513, N31514, N31516, N31517, N31518, N31519, N31520, N31521, N31522, N31524, N31525, N31527, N31528, N31529, N31532, N31533, N31535, N31536, N31537, N31538, N31540, N31541, N31542, N31543, N31544, N31546, N31548, N31550, N31551, N31553, N31554, N31556, N31557, N31560, N31561, N31562, N31563, N31565, N31566, N31567, N31568, N31570, N31571, N31573, N31574, N31575, N31576, N31579, N31580, N31581, N31582, N31583, N31584, N31586, N31587, N31588, N31589, N31591, N31593, N31594, N31595, N31596, N31597, N31598, N31600, N31603, N31605, N31606, N31608, N31610, N31614, N31615, N31617, N31618, N31619, N31620, N31621, N31622, N31624, N31627, N31628, N31629, N31630, N31632, N31637, N31638, N31642, N31643, N31645, N31647, N31648, N31649, N31651, N31652, N31653, N31654, N31655, N31656, N31657, N31658, N31659, N31660, N31664, N31665, N31666, N31667, N31668, N31670, N31672, N31673, N31674, N31677, N31679, N31681, N31682, N31684, N31685, N31686, N31687, N31688, N31689, N31691, N31692, N31693, N31694, N31695, N31696, N31697, N31698, N31699, N31700, N31701, N31703, N31704, N31705, N31706, N31707, N31708, N31710, N31711, N31712, N31714, N31715, N31717, N31718, N31719, N31720, N31724, N31725, N31728, N31731, N31734, N31736, N31737, N31738, N31740, N31742, N31744, N31745, N31746, N31749, N31752, N31753, N31754, N31757, N31759, N31760, N31761, N31762, N31763, N31764, N31765, N31766, N31767, N31768, N31771, N31772, N31773, N31775, N31776, N31777, N31778, N31781, N31783, N31785, N31787, N31788, N31789, N31790, N31791, N31793, N31794, N31797, N31801, N31802, N31803, N31805, N31806, N31807, N31808, N31810, N31811, N31812, N31813, N31814, N31815, N31817, N31818, N31819, N31820, N31821, N31822, N31823, N31824, N31825, N31826, N31827, N31828, N31829, N31830, N31831, N31833, N31834, N31836, N31837, N31840, N31841, N31842, N31843, N31845, N31846, N31848, N31849, N31850, N31851, N31852, N31854, N31855, N31857, N31858, N31859, N31860, N31865, N31867, N31868, N31870, N31871, N31872, N31873, N31875, N31876, N31880, N31881, N31882, N31883, N31884, N31885, N31887, N31888, N31890, N31891, N31892, N31895, N31896, N31899, N31900, N31903, N31904, N31906, N31907, N31908, N31910, N31911, N31912, N31913, N31915, N31916, N31918, N31920, N31922, N31924, N31925, N31928, N31929, N31930, N31932, N31933, N31937, N31939, N31940, N31941, N31942, N31944, N31945, N31946, N31947, N31948, N31949, N31950, N31953, N31954, N31956, N31957, N31959, N31960, N31962, N31963, N31964, N31965, N31966, N31967, N31969, N31971, N31973, N31974, N31976, N31977, N31979, N31981, N31982, N31983, N31984, N31985, N31988, N31989, N31990, N31991, N31992, N31994, N31996, N31998, N31999, N32000, N32001, N32002, N32004, N32007, N32010, N32012, N32013, N32014, N32015, N32017, N32018, N32019, N32020, N32021, N32026, N32027, N32028, N32030, N32032, N32034, N32036, N32037, N32038, N32040, N32041, N32042, N32045, N32047, N32048, N32050, N32051, N32053, N32054, N32055, N32056, N32057, N32058, N32059, N32062, N32064, N32065, N32066, N32068, N32069, N32070, N32073, N32075, N32076, N32077, N32078, N32079, N32080, N32081, N32082, N32083, N32084, N32087, N32088, N32089, N32090, N32092, N32093, N32097, N32098, N32099, N32101, N32104, N32105, N32106, N32108, N32109, N32110, N32111, N32114, N32117, N32118, N32119, N32121, N32124, N32127, N32129, N32130, N32134, N32135, N32136, N32137, N32138, N32141, N32143, N32144, N32145, N32146, N32147, N32148, N32150, N32151, N32152, N32153, N32154, N32155, N32160, N32161, N32162, N32164, N32165, N32167, N32171, N32173, N32174, N32175, N32176, N32177, N32179, N32182, N32183, N32184, N32186, N32187, N32189, N32190, N32192, N32193, N32195, N32199, N32200, N32201, N32203, N32209, N32210, N32212, N32214, N32216, N32218, N32219, N32222, N32223, N32224, N32225, N32226, N32228, N32229, N32230, N32232, N32233, N32234, N32235, N32236, N32237, N32238, N32240, N32243, N32244, N32246, N32247, N32249, N32250, N32251, N32252, N32253, N32255, N32257, N32259, N32260, N32262, N32263, N32264, N32265, N32266, N32267, N32269, N32272, N32273, N32274, N32275, N32276, N32277, N32278, N32279, N32280, N32282, N32283, N32287, N32288, N32290, N32291, N32292, N32293, N32294, N32295, N32296, N32298, N32301, N32302, N32303, N32304, N32305, N32308, N32309, N32310, N32311, N32312, N32313, N32314, N32315, N32316, N32317, N32318, N32319, N32320, N32321, N32325, N32327, N32328, N32329, N32330, N32333, N32336, N32337, N32339, N32340, N32341, N32342, N32343, N32345, N32346, N32347, N32348, N32349, N32350, N32351, N32352, N32353, N32354, N32355, N32356, N32357, N32359, N32361, N32362, N32363, N32365, N32367, N32369, N32370, N32372, N32373, N32374, N32377, N32378, N32379, N32380, N32382, N32383, N32384, N32385, N32386, N32387, N32388, N32389, N32392, N32393, N32394, N32396, N32397, N32399, N32400, N32401, N32404, N32405, N32406, N32407, N32408, N32409, N32410, N32411, N32412, N32416, N32418, N32419, N32420, N32421, N32422, N32424, N32425, N32426, N32427, N32428, N32429, N32430, N32431, N32432, N32433, N32434, N32435, N32437, N32438, N32439, N32440, N32441, N32442, N32444, N32445, N32446, N32447, N32448, N32449, N32451, N32454, N32455, N32456, N32459, N32460, N32461, N32464, N32465, N32466, N32469, N32471, N32472, N32473, N32474, N32475, N32476, N32480, N32481, N32482, N32483, N32489, N32490, N32491, N32492, N32494, N32496, N32498, N32500, N32501, N32502, N32505, N32506, N32507, N32508, N32511, N32513, N32514, N32517, N32519, N32521, N32522, N32525, N32526, N32527, N32528, N32531, N32532, N32535, N32539, N32540, N32542, N32543, N32544, N32547, N32548, N32550, N32552, N32553, N32554, N32557, N32558, N32559, N32560, N32562, N32563, N32564, N32565, N32567, N32568, N32570, N32573, N32575, N32576, N32577, N32579, N32581, N32582, N32583, N32584, N32585, N32586, N32587, N32589, N32590, N32592, N32593, N32595, N32597, N32598, N32599, N32600, N32602, N32603, N32604, N32606, N32607, N32608, N32610, N32613, N32615, N32616, N32617, N32618, N32619, N32621, N32622, N32623, N32624, N32625, N32626, N32628, N32629, N32631, N32633, N32634, N32635, N32637, N32638, N32639, N32640, N32641, N32642, N32643, N32644, N32645, N32650, N32652, N32653, N32654, N32655, N32656, N32657, N32658, N32661, N32662, N32663, N32665, N32666, N32667, N32668, N32669, N32670, N32671, N32673, N32674, N32676, N32677, N32678, N32679, N32682, N32685, N32686, N32689, N32690, N32691, N32693, N32694, N32695, N32696, N32698, N32700, N32702, N32703, N32704, N32705, N32706, N32707, N32709, N32710, N32712, N32713, N32714, N32716, N32718, N32719, N32720, N32722, N32723, N32725, N32726, N32728, N32730, N32731, N32732, N32733, N32735, N32736, N32737, N32738, N32740, N32741, N32742, N32743, N32744, N32745, N32747, N32748, N32749, N32750, N32752, N32754, N32755, N32756, N32758, N32759, N32760, N32762, N32763, N32764, N32765, N32769, N32770, N32771, N32772, N32773, N32774, N32777, N32778, N32779, N32781, N32782, N32784, N32785, N32786, N32787, N32788, N32789, N32790, N32792, N32793, N32794, N32795, N32796, N32797, N32798, N32799, N32800, N32801, N32802, N32804, N32807, N32809, N32810, N32811, N32812, N32813, N32814, N32817, N32818, N32819, N32820, N32821, N32822, N32823, N32824, N32825, N32828, N32829, N32830, N32832, N32833, N32834, N32837, N32838, N32841, N32842, N32846, N32848, N32849, N32850, N32851, N32852, N32853, N32854, N32858, N32859, N32860, N32862, N32863, N32866, N32867, N32868, N32869, N32871, N32872, N32873, N32874, N32875, N32876, N32877, N32878, N32879, N32880, N32881, N32882, N32883, N32884, N32885, N32886, N32887, N32888, N32890, N32892, N32893, N32896, N32899, N32900, N32901, N32905, N32906, N32907, N32908, N32909, N32911, N32912, N32916, N32917, N32918, N32920, N32923, N32924, N32926, N32930, N32931, N32935, N32936, N32937, N32939, N32940, N32942, N32943, N32944, N32946, N32947, N32948, N32949, N32950, N32952, N32953, N32956, N32957, N32958, N32960, N32965, N32966, N32968, N32969, N32970, N32971, N32972, N32973, N32977, N32978, N32979, N32980, N32982, N32983, N32985, N32986, N32987, N32988, N32990, N32991, N32993, N32994, N32995, N32998, N32999, N33000, N33001, N33002, N33005, N33006, N33007, N33009, N33010, N33012, N33013, N33016, N33018, N33020, N33021, N33022, N33024, N33025, N33026, N33027, N33028, N33029, N33031, N33032, N33034, N33035, N33036, N33037, N33038, N33040, N33044, N33045, N33046, N33047, N33049, N33054, N33055, N33056, N33057, N33058, N33061, N33063, N33064, N33068, N33072, N33073, N33075, N33077, N33078, N33079, N33082, N33083, N33084, N33085, N33087, N33088, N33091, N33092, N33093, N33096, N33098, N33099, N33101, N33105, N33107, N33108, N33109, N33110, N33111, N33112, N33113, N33114, N33115, N33116, N33117, N33119, N33120, N33122, N33124, N33125, N33126, N33127, N33129, N33131, N33132, N33133, N33136, N33138, N33141, N33142, N33143, N33144, N33145, N33146, N33149, N33150, N33151, N33152, N33156, N33157, N33158, N33159, N33160, N33162, N33163, N33164, N33165, N33167, N33168, N33170, N33171, N33173, N33174, N33175, N33177, N33178, N33179, N33180, N33181, N33182, N33183, N33185, N33186, N33188, N33189, N33190, N33191, N33192, N33193, N33194, N33195, N33196, N33197, N33198, N33202, N33203, N33206, N33208, N33209, N33211, N33215, N33216, N33217, N33220, N33221, N33223, N33224, N33226, N33227, N33229, N33231, N33232, N33233, N33234, N33236, N33238, N33240, N33241, N33242, N33244, N33245, N33247, N33248, N33249, N33250, N33253, N33254, N33256, N33257, N33259, N33262, N33263, N33264, N33265, N33266, N33267, N33269, N33274, N33277, N33279, N33282, N33284, N33285, N33287, N33288, N33289, N33291, N33292, N33293, N33294, N33295, N33297, N33299, N33300, N33301, N33302, N33304, N33305, N33306, N33307, N33309, N33310, N33311, N33313, N33315, N33316, N33317, N33318, N33319, N33320, N33321, N33324, N33325, N33327, N33329, N33330, N33331, N33332, N33335, N33336, N33337, N33338, N33339, N33340, N33341, N33342, N33343, N33344, N33345, N33346, N33347, N33348, N33349, N33351, N33352, N33353, N33354, N33355, N33356, N33358, N33359, N33360, N33361, N33362, N33363, N33364, N33365, N33366, N33367, N33368, N33369, N33372, N33373, N33374, N33377, N33378, N33379, N33380, N33384, N33385, N33386, N33387, N33388, N33392, N33396, N33398, N33400, N33401, N33404, N33405, N33406, N33407, N33408, N33410, N33411, N33413, N33414, N33415, N33416, N33418, N33419, N33422, N33423, N33424, N33427, N33431, N33432, N33433, N33434, N33436, N33437, N33441, N33442, N33443, N33446, N33447, N33448, N33450, N33451, N33452, N33453, N33455, N33457, N33458, N33462, N33463, N33464, N33466, N33467, N33468, N33469, N33474, N33476, N33477, N33479, N33481, N33485, N33486, N33487, N33489, N33490, N33491, N33492, N33493, N33496, N33497, N33500, N33501, N33502, N33503, N33504, N33506, N33508, N33509, N33510, N33511, N33513, N33514, N33515, N33516, N33517, N33518, N33519, N33521, N33522, N33524, N33526, N33527, N33528, N33529, N33530, N33531, N33532, N33534, N33536, N33537, N33538, N33539, N33540, N33543, N33546, N33547, N33548, N33550, N33551, N33552, N33553, N33554, N33555, N33556, N33557, N33559, N33560, N33561, N33562, N33563, N33564, N33565, N33568, N33570, N33573, N33574, N33576, N33577, N33578, N33579, N33583, N33584, N33586, N33587, N33588, N33590, N33593, N33594, N33599, N33606, N33609, N33610, N33611, N33613, N33614, N33616, N33618, N33619, N33620, N33621, N33622, N33623, N33625, N33626, N33627, N33628, N33629, N33630, N33631, N33635, N33637, N33639, N33640, N33641, N33642, N33643, N33646, N33647, N33650, N33651, N33652, N33653, N33654, N33655, N33656, N33657, N33658, N33659, N33660, N33661, N33663, N33670, N33672, N33673, N33674, N33675, N33677, N33678, N33679, N33680, N33681, N33683, N33684, N33685, N33687, N33689, N33691, N33692, N33693, N33694, N33695, N33697, N33700, N33701, N33703, N33705, N33706, N33707, N33708, N33709, N33710, N33711, N33712, N33713, N33714, N33718, N33720, N33721, N33722, N33723, N33724, N33725, N33726, N33727, N33729, N33730, N33731, N33733, N33734, N33735, N33738, N33740, N33741, N33742, N33743, N33745, N33746, N33747, N33749, N33750, N33751, N33752, N33753, N33754, N33755, N33757, N33758, N33759, N33761, N33763, N33764, N33765, N33766, N33767, N33769, N33772, N33773, N33774, N33775, N33776, N33777, N33778, N33779, N33780, N33782, N33783, N33784, N33785, N33786, N33787, N33788, N33789, N33792, N33793, N33794, N33795, N33796, N33797, N33798, N33799, N33800, N33801, N33802, N33803, N33804, N33805, N33807, N33809, N33811, N33812, N33813, N33814, N33815, N33818, N33820, N33821, N33822, N33824, N33825, N33826, N33827, N33828, N33829, N33830, N33832, N33833, N33835, N33836, N33837, N33839, N33841, N33842, N33844, N33846, N33848, N33849, N33850, N33851, N33852, N33853, N33854, N33856, N33858, N33859, N33861, N33862, N33863, N33864, N33866, N33867, N33869, N33870, N33871, N33872, N33873, N33875, N33876, N33877, N33878, N33879, N33880, N33881, N33882, N33884, N33888, N33889, N33890, N33891, N33892, N33896, N33897, N33898, N33899, N33900, N33901, N33903, N33904, N33905, N33906, N33907, N33908, N33909, N33911, N33914, N33915, N33916, N33917, N33919, N33921, N33922, N33925, N33927, N33928, N33929, N33930, N33933, N33934, N33935, N33936, N33937, N33940, N33943, N33944, N33945, N33946, N33947, N33948, N33949, N33950, N33951, N33952, N33953, N33955, N33956, N33960, N33961, N33963, N33965, N33966, N33967, N33968, N33969, N33970, N33971, N33972, N33973, N33974, N33975, N33976, N33977, N33978, N33979, N33980, N33983, N33984, N33985, N33986, N33987, N33990, N33992, N33993, N33994, N33995, N33996, N33997, N33998, N34000, N34001, N34002, N34003, N34004, N34005, N34006, N34008, N34009, N34010, N34011, N34016, N34019, N34020, N34021, N34023, N34024, N34025, N34026, N34028, N34031, N34032, N34033, N34035, N34036, N34037, N34039, N34040, N34042, N34043, N34044, N34045, N34046, N34047, N34049, N34050, N34052, N34053, N34054, N34055, N34057, N34058, N34059, N34060, N34061, N34062, N34063, N34065, N34066, N34067, N34068, N34070, N34072, N34073, N34074, N34076, N34077, N34081, N34082, N34084, N34085, N34088, N34090, N34092, N34093, N34095, N34096, N34097, N34098, N34100, N34102, N34103, N34105, N34106, N34107, N34108, N34109, N34110, N34112, N34114, N34115, N34116, N34117, N34118, N34119, N34120, N34121, N34122, N34123, N34124, N34125, N34127, N34128, N34129, N34130, N34131, N34132, N34133, N34135, N34136, N34137, N34141, N34142, N34143, N34145, N34146, N34147, N34148, N34149, N34150, N34151, N34153, N34155, N34156, N34158, N34160, N34161, N34163, N34165, N34166, N34170, N34171, N34174, N34177, N34178, N34179, N34180, N34181, N34183, N34184, N34185, N34186, N34187, N34188, N34189, N34193, N34195, N34196, N34197, N34198, N34199, N34201, N34202, N34205, N34206, N34209, N34210, N34212, N34214, N34217, N34218, N34221, N34223, N34225, N34228, N34229, N34231, N34232, N34233, N34235, N34236, N34237, N34239, N34240, N34242, N34243, N34244, N34245, N34246, N34247, N34248, N34250, N34251, N34252, N34253, N34257, N34259, N34260, N34261, N34263, N34265, N34266, N34267, N34270, N34271, N34274, N34276, N34277, N34278, N34279, N34281, N34282, N34284, N34285, N34287, N34289, N34290, N34292, N34293, N34294, N34295, N34296, N34298, N34299, N34300, N34301, N34302, N34303, N34305, N34306, N34307, N34309, N34310, N34312, N34313, N34314, N34316, N34318, N34319, N34321, N34322, N34323, N34324, N34325, N34330, N34331, N34334, N34336, N34337, N34338, N34341, N34343, N34344, N34345, N34346, N34347, N34350, N34351, N34352, N34355, N34356, N34358, N34359, N34361, N34363, N34364, N34365, N34369, N34371, N34372, N34373, N34374, N34375, N34376, N34378, N34379, N34380, N34384, N34386, N34388, N34389, N34390, N34392, N34393, N34396, N34397, N34399, N34400, N34401, N34403, N34405, N34406, N34409, N34410, N34411, N34412, N34413, N34414, N34416, N34417, N34418, N34419, N34420, N34421, N34422, N34424, N34425, N34426, N34427, N34430, N34432, N34433, N34435, N34436, N34437, N34439, N34440, N34442, N34445, N34446, N34447, N34448, N34449, N34450, N34451, N34454, N34455, N34456, N34457, N34458, N34459, N34460, N34461, N34462, N34463, N34466, N34467, N34468, N34469, N34470, N34471, N34473, N34478, N34480, N34481, N34484, N34487, N34488, N34490, N34493, N34494, N34495, N34496, N34497, N34498, N34499, N34500, N34501, N34502, N34503, N34505, N34508, N34512, N34514, N34517, N34519, N34521, N34522, N34523, N34525, N34526, N34527, N34528, N34531, N34532, N34533, N34534, N34535, N34536, N34537, N34539, N34540, N34541, N34542, N34544, N34545, N34546, N34547, N34548, N34549, N34552, N34554, N34555, N34556, N34557, N34558, N34560, N34561, N34563, N34564, N34565, N34566, N34567, N34568, N34569, N34570, N34571, N34572, N34574, N34576, N34577, N34578, N34579, N34580, N34581, N34583, N34585, N34586, N34587, N34589, N34590, N34591, N34593, N34594, N34595, N34596, N34597, N34598, N34599, N34600, N34602, N34604, N34605, N34606, N34608, N34612, N34613, N34614, N34616, N34618, N34619, N34622, N34623, N34624, N34625, N34626, N34627, N34628, N34629, N34630, N34631, N34633, N34636, N34637, N34638, N34640, N34641, N34642, N34643, N34644, N34646, N34647, N34648, N34649, N34650, N34653, N34655, N34657, N34659, N34660, N34662, N34663, N34665, N34667, N34670, N34671, N34672, N34673, N34674, N34675, N34677, N34678, N34679, N34680, N34681, N34682, N34683, N34685, N34686, N34687, N34688, N34689, N34693, N34697, N34698, N34699, N34701, N34703, N34704, N34705, N34707, N34708, N34711, N34712, N34713, N34719, N34720, N34722, N34724, N34725, N34726, N34727, N34728, N34729, N34730, N34731, N34732, N34735, N34738, N34741, N34742, N34743, N34744, N34745, N34746, N34748, N34749, N34750, N34751, N34752, N34753, N34754, N34756, N34758, N34763, N34764, N34766, N34767, N34769, N34771, N34772, N34773, N34774, N34775, N34777, N34778, N34780, N34781, N34787, N34788, N34789, N34794, N34795, N34796, N34797, N34799, N34800, N34804, N34806, N34807, N34808, N34809, N34810, N34811, N34814, N34815, N34818, N34821, N34822, N34823, N34826, N34827, N34829, N34830, N34831, N34832, N34833, N34836, N34837, N34839, N34840, N34841, N34842, N34844, N34845, N34847, N34848, N34850, N34851, N34853, N34854, N34855, N34856, N34857, N34861, N34863, N34865, N34867, N34868, N34869, N34870, N34871, N34874, N34877, N34878, N34879, N34881, N34882, N34883, N34885, N34886, N34889, N34891, N34893, N34895, N34896, N34897, N34898, N34899, N34900, N34901, N34903, N34904, N34906, N34907, N34908, N34909, N34910, N34911, N34912, N34913, N34914, N34915, N34917, N34918, N34919, N34920, N34921, N34922, N34923, N34925, N34926, N34928, N34929, N34932, N34933, N34934, N34937, N34938, N34939, N34940, N34944, N34945, N34946, N34948, N34951, N34953, N34954, N34956, N34957, N34958, N34959, N34960, N34961, N34962, N34963, N34965, N34967, N34968, N34970, N34977, N34978, N34979, N34982, N34983, N34984, N34985, N34986, N34987, N34988, N34990, N34992, N34993, N34994, N34995, N34996, N34999, N35000, N35001, N35002, N35005, N35006, N35007, N35009, N35013, N35015, N35017, N35018, N35019, N35020, N35021, N35022, N35024, N35025, N35026, N35027, N35028, N35029, N35030, N35032, N35033, N35034, N35035, N35036, N35039, N35042, N35043, N35045, N35046, N35048, N35049, N35050, N35052, N35053, N35054, N35055, N35056, N35057, N35058, N35059, N35060, N35062, N35063, N35064, N35065, N35066, N35067, N35069, N35070, N35071, N35073, N35074, N35077, N35078, N35082, N35083, N35085, N35086, N35087, N35088, N35089, N35091, N35092, N35093, N35095, N35096, N35097, N35098, N35099, N35100, N35101, N35103, N35104, N35107, N35108, N35109, N35110, N35111, N35113, N35115, N35117, N35118, N35119, N35120, N35123, N35125, N35126, N35128, N35129, N35131, N35132, N35133, N35134, N35135, N35136, N35139, N35140, N35143, N35144, N35145, N35146, N35147, N35148, N35149, N35150, N35151, N35152, N35153, N35154, N35155, N35156, N35159, N35160, N35161, N35163, N35166, N35167, N35168, N35169, N35171, N35172, N35173, N35174, N35175, N35176, N35177, N35178, N35179, N35180, N35181, N35185, N35186, N35187, N35188, N35189, N35190, N35191, N35192, N35193, N35196, N35197, N35198, N35199, N35200, N35203, N35204, N35206, N35207, N35208, N35209, N35210, N35211, N35212, N35215, N35217, N35218, N35220, N35221, N35222, N35224, N35225, N35227, N35228, N35230, N35232, N35234, N35236, N35237, N35239, N35240, N35241, N35242, N35244, N35246, N35247, N35248, N35249, N35252, N35253, N35254, N35256, N35257, N35258, N35259, N35260, N35261, N35262, N35263, N35264, N35265, N35266, N35267, N35268, N35269, N35275, N35278, N35279, N35280, N35281, N35282, N35283, N35284, N35286, N35288, N35289, N35290, N35291, N35295, N35296, N35298, N35299, N35300, N35301, N35302, N35304, N35305, N35308, N35309, N35310, N35311, N35313, N35314, N35315, N35318, N35319, N35321, N35322, N35323, N35324, N35326, N35327, N35328, N35330, N35331, N35332, N35333, N35334, N35337, N35338, N35340, N35342, N35343, N35344, N35345, N35346, N35349, N35350, N35351, N35352, N35353, N35354, N35355, N35356, N35357, N35358, N35359, N35362, N35363, N35366, N35368, N35370, N35371, N35373, N35374, N35375, N35376, N35377, N35378, N35379, N35380, N35381, N35383, N35384, N35385, N35386, N35387, N35388, N35389, N35391, N35392, N35394, N35395, N35396, N35398, N35399, N35400, N35401, N35402, N35403, N35406, N35407, N35408, N35409, N35411, N35413, N35414, N35415, N35416, N35417, N35418, N35419, N35422, N35423, N35424, N35425, N35427, N35428, N35429, N35431, N35433, N35435, N35436, N35438, N35439, N35440, N35441, N35442, N35443, N35444, N35445, N35446, N35448, N35449, N35453, N35456, N35457, N35458, N35459, N35460, N35463, N35464, N35467, N35468, N35469, N35470, N35471, N35472, N35474, N35476, N35477, N35479, N35481, N35482, N35485, N35486, N35488, N35490, N35492, N35495, N35496, N35497, N35498, N35499, N35500, N35501, N35502, N35503, N35504, N35507, N35508, N35511, N35512, N35513, N35514, N35516, N35517, N35519, N35521, N35522, N35524, N35525, N35526, N35527, N35529, N35530, N35531, N35532, N35533, N35534, N35536, N35538, N35542, N35544, N35545, N35547, N35548, N35549, N35550, N35551, N35553, N35554, N35555, N35557, N35558, N35560, N35561, N35563, N35564, N35565, N35567, N35569, N35570, N35571, N35573, N35574, N35575, N35576, N35577, N35578, N35579, N35582, N35583, N35584, N35585, N35586, N35587, N35588, N35589, N35591, N35592, N35593, N35594, N35595, N35596, N35598, N35600, N35601, N35603, N35604, N35605, N35606, N35608, N35609, N35611, N35612, N35613, N35615, N35618, N35619, N35620, N35621, N35623, N35624, N35625, N35626, N35627, N35629, N35630, N35631, N35632, N35633, N35635, N35637, N35642, N35643, N35645, N35647, N35649, N35650, N35652, N35653, N35655, N35659, N35661, N35663, N35665, N35666, N35668, N35669, N35670, N35672, N35674, N35675, N35676, N35677, N35678, N35680, N35681, N35682, N35684, N35687, N35690, N35691, N35692, N35694, N35695, N35697, N35698, N35700, N35701, N35702, N35703, N35704, N35705, N35707, N35710, N35711, N35715, N35716, N35718, N35720, N35721, N35722, N35723, N35724, N35725, N35726, N35728, N35731, N35732, N35734, N35735, N35737, N35739, N35740, N35743, N35745, N35747, N35749, N35751, N35752, N35754, N35755, N35756, N35757, N35758, N35759, N35760, N35762, N35764, N35766, N35767, N35768, N35769, N35770, N35771, N35776, N35777, N35779, N35781, N35782, N35785, N35786, N35791, N35793, N35795, N35796, N35797, N35798, N35799, N35800, N35801, N35802, N35803, N35804, N35805, N35806, N35807, N35808, N35811, N35814, N35815, N35816, N35818, N35820, N35821, N35822, N35823, N35828, N35831, N35832, N35833, N35835, N35836, N35837, N35838, N35840, N35841, N35842, N35843, N35844, N35845, N35846, N35847, N35848, N35849, N35851, N35852, N35853, N35855, N35856, N35858, N35860, N35861, N35862, N35863, N35864, N35865, N35868, N35869, N35870, N35872, N35875, N35876, N35878, N35880, N35884, N35885, N35889, N35891, N35892, N35893, N35894, N35895, N35896, N35897, N35898, N35899, N35900, N35901, N35903, N35905, N35906, N35907, N35908, N35910, N35911, N35913, N35914, N35917, N35918, N35919, N35921, N35923, N35924, N35926, N35927, N35929, N35931, N35932, N35933, N35934, N35935, N35936, N35938, N35940, N35941, N35943, N35944, N35947, N35948, N35949, N35950, N35952, N35953, N35954, N35955, N35957, N35958, N35959, N35961, N35962, N35965, N35966, N35971, N35972, N35973, N35974, N35975, N35977, N35979, N35980, N35981, N35982, N35983, N35984, N35986, N35987, N35988, N35989, N35992, N35994, N35995, N35996, N35998, N36000, N36001, N36002, N36003, N36004, N36005, N36006, N36008, N36011, N36013, N36016, N36017, N36019, N36020, N36022, N36024, N36025, N36026, N36027, N36029, N36030, N36031, N36035, N36036, N36037, N36038, N36041, N36042, N36043, N36044, N36047, N36048, N36050, N36051, N36052, N36053, N36055, N36057, N36058, N36059, N36060, N36061, N36063, N36065, N36066, N36068, N36069, N36070, N36072, N36073, N36074, N36076, N36077, N36080, N36081, N36083, N36086, N36087, N36089, N36091, N36092, N36093, N36094, N36097, N36098, N36100, N36102, N36103, N36105, N36106, N36107, N36108, N36109, N36111, N36112, N36113, N36114, N36115, N36116, N36117, N36118, N36121, N36122, N36123, N36124, N36125, N36127, N36130, N36131, N36133, N36134, N36135, N36138, N36139, N36140, N36141, N36143, N36145, N36146, N36148, N36150, N36151, N36153, N36154, N36155, N36158, N36159, N36160, N36161, N36163, N36164, N36169, N36170, N36172, N36174, N36175, N36176, N36177, N36178, N36180, N36181, N36182, N36186, N36187, N36188, N36189, N36191, N36192, N36193, N36194, N36195, N36196, N36197, N36198, N36201, N36202, N36205, N36206, N36209, N36210, N36212, N36214, N36215, N36216, N36219, N36222, N36224, N36225, N36226, N36227, N36228, N36229, N36230, N36231, N36232, N36233, N36234, N36235, N36236, N36238, N36239, N36241, N36242, N36246, N36247, N36249, N36250, N36251, N36252, N36256, N36257, N36259, N36260, N36261, N36262, N36263, N36264, N36265, N36266, N36267, N36271, N36272, N36273, N36274, N36275, N36276, N36277, N36278, N36279, N36281, N36282, N36284, N36285, N36286, N36288, N36289, N36293, N36294, N36295, N36296, N36298, N36300, N36301, N36304, N36307, N36308, N36309, N36313, N36315, N36317, N36318, N36319, N36322, N36325, N36326, N36328, N36329, N36330, N36331, N36333, N36336, N36337, N36338, N36339, N36341, N36342, N36344, N36345, N36346, N36347, N36348, N36351, N36353, N36354, N36355, N36356, N36358, N36362, N36363, N36364, N36365, N36366, N36367, N36368, N36371, N36372, N36373, N36374, N36376, N36378, N36380, N36381, N36383, N36385, N36387, N36388, N36390, N36391, N36393, N36394, N36395, N36396, N36398, N36400, N36401, N36403, N36404, N36406, N36408, N36410, N36412, N36413, N36415, N36416, N36419, N36420, N36421, N36422, N36423, N36424, N36425, N36426, N36427, N36428, N36429, N36430, N36431, N36432, N36433, N36434, N36435, N36436, N36437, N36439, N36442, N36443, N36448, N36451, N36452, N36453, N36455, N36456, N36457, N36458, N36463, N36464, N36465, N36466, N36467, N36468, N36469, N36470, N36471, N36472, N36473, N36474, N36475, N36477, N36478, N36480, N36481, N36482, N36483, N36484, N36488, N36489, N36490, N36491, N36492, N36493, N36497, N36498, N36499, N36500, N36501, N36502, N36503, N36505, N36506, N36507, N36512, N36515, N36516, N36518, N36519, N36521, N36522, N36524, N36525, N36526, N36527, N36528, N36529, N36531, N36532, N36534, N36536, N36537, N36539, N36540, N36542, N36543, N36545, N36546, N36548, N36549, N36552, N36553, N36554, N36556, N36557, N36558, N36560, N36561, N36562, N36563, N36564, N36565, N36566, N36567, N36569, N36570, N36571, N36575, N36576, N36577, N36578, N36580, N36583, N36584, N36585, N36587, N36588, N36592, N36594, N36595, N36596, N36597, N36598, N36599, N36600, N36601, N36602, N36603, N36604, N36605, N36607, N36608, N36609, N36610, N36611, N36613, N36615, N36617, N36618, N36619, N36621, N36622, N36623, N36624, N36625, N36626, N36627, N36629, N36630, N36633, N36634, N36635, N36636, N36638, N36639, N36640, N36642, N36644, N36645, N36646, N36647, N36649, N36650, N36651, N36653, N36654, N36655, N36656, N36657, N36661, N36662, N36663, N36664, N36665, N36666, N36667, N36668, N36669, N36671, N36672, N36673, N36674, N36675, N36677, N36678, N36679, N36680, N36682, N36683, N36684, N36686, N36687, N36688, N36689, N36691, N36695, N36697, N36699, N36701, N36702, N36703, N36705, N36706, N36707, N36709, N36711, N36713, N36715, N36716, N36717, N36718, N36719, N36720, N36721, N36722, N36723, N36724, N36725, N36727, N36729, N36730, N36733, N36734, N36735, N36737, N36738, N36740, N36742, N36743, N36744, N36746, N36747, N36748, N36749, N36752, N36754, N36755, N36756, N36758, N36760, N36764, N36765, N36767, N36768, N36769, N36770, N36771, N36773, N36774, N36777, N36778, N36779, N36780, N36782, N36783, N36784, N36785, N36786, N36787, N36788, N36789, N36791, N36793, N36795, N36797, N36798, N36799, N36803, N36804, N36805, N36806, N36807, N36808, N36809, N36810, N36811, N36812, N36813, N36816, N36817, N36818, N36820, N36821, N36822, N36823, N36824, N36825, N36828, N36829, N36831, N36834, N36835, N36839, N36840, N36842, N36845, N36846, N36848, N36850, N36851, N36852, N36853, N36854, N36855, N36858, N36859, N36861, N36862, N36863, N36864, N36865, N36866, N36867, N36869, N36870, N36871, N36872, N36873, N36874, N36879, N36880, N36881, N36882, N36886, N36887, N36888, N36889, N36890, N36891, N36892, N36893, N36896, N36897, N36898, N36900, N36902, N36906, N36907, N36908, N36909, N36910, N36911, N36912, N36915, N36916, N36917, N36918, N36920, N36921, N36922, N36923, N36925, N36926, N36928, N36929, N36930, N36931, N36932, N36933, N36934, N36936, N36937, N36938, N36939, N36946, N36948, N36949, N36950, N36951, N36952, N36954, N36955, N36956, N36958, N36959, N36960, N36961, N36962, N36964, N36967, N36970, N36972, N36977, N36978, N36980, N36981, N36982, N36985, N36990, N36991, N36992, N36995, N36998, N36999, N37000, N37001, N37002, N37003, N37004, N37006, N37011, N37013, N37014, N37016, N37017, N37018, N37019, N37020, N37021, N37023, N37024, N37025, N37026, N37028, N37029, N37031, N37032, N37035, N37037, N37038, N37039, N37042, N37043, N37044, N37046, N37048, N37052, N37053, N37054, N37055, N37059, N37061, N37063, N37065, N37066, N37067, N37068, N37070, N37071, N37075, N37079, N37083, N37084, N37085, N37087, N37088, N37089, N37090, N37091, N37092, N37093, N37094, N37097, N37099, N37100, N37103, N37108, N37109, N37111, N37113, N37115, N37117, N37120, N37121, N37123, N37124, N37125, N37128, N37131, N37137, N37139, N37140, N37141, N37142, N37144, N37145, N37148, N37149, N37150, N37152, N37153, N37154, N37155, N37156, N37157, N37158, N37159, N37161, N37162, N37163, N37164, N37165, N37166, N37167, N37169, N37170, N37171, N37173, N37176, N37177, N37179, N37180, N37181, N37182, N37185, N37186, N37187, N37192, N37193, N37194, N37195, N37196, N37197, N37198, N37199, N37200, N37201, N37202, N37204, N37205, N37206, N37211, N37212, N37213, N37214, N37215, N37216, N37218, N37220, N37222, N37226, N37228, N37230, N37231, N37232, N37234, N37235, N37237, N37238, N37239, N37242, N37243, N37244, N37245, N37247, N37248, N37249, N37251, N37252, N37253, N37254, N37256, N37260, N37264, N37265, N37266, N37267, N37269, N37271, N37272, N37273, N37274, N37275, N37276, N37277, N37278, N37279, N37280, N37282, N37284, N37285, N37286, N37288, N37289, N37290, N37294, N37297, N37299, N37300, N37302, N37304, N37305, N37306, N37307, N37308, N37309, N37310, N37311, N37312, N37313, N37316, N37319, N37320, N37321, N37322, N37324, N37325, N37326, N37327, N37328, N37331, N37334, N37335, N37336, N37338, N37339, N37341, N37342, N37343, N37345, N37346, N37347, N37348, N37349, N37350, N37351, N37352, N37353, N37354, N37355, N37358, N37359, N37360, N37363, N37365, N37366, N37368, N37371, N37373, N37374, N37375, N37376, N37377, N37378, N37379, N37380, N37381, N37382, N37383, N37386, N37387, N37388, N37389, N37390, N37391, N37392, N37393, N37394, N37399, N37401, N37402, N37403, N37404, N37405, N37407, N37408, N37409, N37410, N37411, N37414, N37415, N37417, N37418, N37419, N37420, N37421, N37424, N37425, N37426, N37427, N37428, N37430, N37432, N37433, N37434, N37435, N37437, N37438, N37439, N37440, N37442, N37443, N37444, N37445, N37446, N37448, N37450, N37453, N37454, N37455, N37457, N37460, N37463, N37464, N37466, N37467, N37469, N37470, N37475, N37477, N37479, N37480, N37481, N37482, N37483, N37485, N37486, N37488, N37490, N37492, N37496, N37497, N37498, N37500, N37501, N37502, N37503, N37504, N37505, N37506, N37508, N37509, N37512, N37513, N37514, N37515, N37517, N37518, N37519, N37520, N37521, N37523, N37524, N37526, N37527, N37528, N37529, N37531, N37532, N37533, N37534, N37535, N37536, N37537, N37538, N37540, N37542, N37543, N37545, N37546, N37547, N37548, N37549, N37550, N37551, N37552, N37553, N37554, N37556, N37557, N37558, N37559, N37563, N37564, N37565, N37566, N37571, N37572, N37573, N37574, N37575, N37576, N37578, N37579, N37580, N37581, N37582, N37583, N37584, N37585, N37586, N37588, N37590, N37591, N37592, N37593, N37595, N37596, N37598, N37600, N37601, N37602, N37603, N37604, N37605, N37607, N37608, N37609, N37610, N37611, N37612, N37613, N37614, N37616, N37617, N37618, N37620, N37621, N37622, N37623, N37624, N37625, N37628, N37629, N37630, N37631, N37632, N37633, N37635, N37636, N37638, N37639, N37643, N37644, N37645, N37646, N37647, N37648, N37649, N37650, N37651, N37654, N37655, N37656, N37658, N37659, N37660, N37661, N37663, N37664, N37666, N37668, N37670, N37671, N37672, N37673, N37674, N37677, N37678, N37680, N37684, N37687, N37688, N37690, N37691, N37692, N37693, N37695, N37696, N37697, N37701, N37705, N37707, N37708, N37709, N37710, N37711, N37712, N37713, N37714, N37715, N37716, N37717, N37720, N37723, N37724, N37726, N37727, N37728, N37729, N37730, N37731, N37734, N37736, N37737, N37738, N37739, N37740, N37742, N37743, N37745, N37746, N37747, N37748, N37749, N37750, N37751, N37752, N37753, N37754, N37756, N37757, N37759, N37761, N37763, N37764, N37766, N37768, N37769, N37770, N37772, N37773, N37774, N37775, N37776, N37777, N37778, N37779, N37780, N37781, N37782, N37783, N37786, N37788, N37789, N37790, N37791, N37792, N37793, N37795, N37796, N37797, N37798, N37803, N37804, N37806, N37807, N37808, N37809, N37811, N37813, N37814, N37816, N37819, N37820, N37826, N37827, N37828, N37830, N37831, N37832, N37833, N37837, N37838, N37840, N37841, N37844, N37846, N37847, N37851, N37852, N37853, N37854, N37855, N37857, N37858, N37859, N37860, N37861, N37862, N37863, N37864, N37865, N37866, N37867, N37868, N37869, N37871, N37872, N37874, N37875, N37876, N37877, N37878, N37879, N37882, N37884, N37885, N37887, N37888, N37889, N37890, N37891, N37892, N37893, N37894, N37895, N37896, N37898, N37900, N37903, N37904, N37905, N37907, N37908, N37909, N37911, N37912, N37913, N37914, N37915, N37917, N37918, N37919, N37920, N37921, N37922, N37923, N37924, N37927, N37928, N37929, N37930, N37932, N37933, N37934, N37935, N37937, N37938, N37939, N37940, N37941, N37943, N37944, N37945, N37946, N37948, N37949, N37950, N37952, N37953, N37957, N37959, N37960, N37961, N37964, N37965, N37966, N37967, N37968, N37969, N37970, N37971, N37972, N37973, N37977, N37979, N37980, N37981, N37982, N37983, N37986, N37987, N37988, N37989, N37990, N37994, N37998, N37999, N38000, N38003, N38005, N38006, N38009, N38010, N38011, N38012, N38015, N38016, N38017, N38019, N38022, N38023, N38024, N38025, N38026, N38027, N38029, N38030, N38031, N38032, N38033, N38034, N38035, N38040, N38041, N38043, N38045, N38046, N38047, N38048, N38049, N38050, N38051, N38052, N38053, N38054, N38055, N38056, N38057, N38059, N38062, N38063, N38064, N38065, N38066, N38067, N38069, N38071, N38074, N38075, N38077, N38078, N38080, N38082, N38083, N38084, N38088, N38090, N38091, N38092, N38093, N38094, N38095, N38096, N38097, N38098, N38099, N38100, N38103, N38104, N38105, N38108, N38109, N38111, N38113, N38114, N38116, N38117, N38118, N38119, N38121, N38122, N38124, N38125, N38126, N38127, N38128, N38129, N38132, N38133, N38134, N38135, N38136, N38137, N38139, N38141, N38142, N38143, N38144, N38145, N38146, N38147, N38148, N38149, N38150, N38151, N38152, N38153, N38154, N38155, N38157, N38159, N38160, N38161, N38163, N38164, N38166, N38168, N38171, N38175, N38177, N38178, N38179, N38182, N38183, N38186, N38187, N38188, N38189, N38190, N38191, N38192, N38193, N38194, N38196, N38197, N38199, N38202, N38204, N38205, N38206, N38207, N38209, N38210, N38212, N38213, N38217, N38218, N38220, N38221, N38222, N38224, N38225, N38226, N38227, N38228, N38230, N38232, N38233, N38234, N38235, N38237, N38238, N38240, N38243, N38245, N38246, N38247, N38248, N38249, N38250, N38255, N38259, N38260, N38261, N38262, N38263, N38264, N38267, N38268, N38270, N38271, N38275, N38276, N38277, N38278, N38279, N38281, N38283, N38284, N38285, N38287, N38288, N38289, N38290, N38293, N38294, N38296, N38297, N38299, N38302, N38304, N38305, N38307, N38308, N38309, N38312, N38313, N38314, N38315, N38316, N38318, N38319, N38321, N38322, N38324, N38325, N38326, N38328, N38329, N38331, N38332, N38335, N38336, N38337, N38338, N38339, N38340, N38341, N38342, N38345, N38346, N38349, N38350, N38351, N38353, N38354, N38359, N38360, N38362, N38365, N38368, N38369, N38371, N38372, N38374, N38375, N38376, N38378, N38379, N38380, N38381, N38384, N38385, N38386, N38387, N38388, N38389, N38391, N38392, N38393, N38394, N38396, N38397, N38398, N38399, N38400, N38402, N38403, N38404, N38405, N38407, N38408, N38409, N38410, N38411, N38412, N38413, N38415, N38416, N38418, N38419, N38421, N38422, N38423, N38424, N38426, N38427, N38428, N38429, N38430, N38431, N38433, N38434, N38435, N38436, N38437, N38438, N38439, N38440, N38443, N38444, N38445, N38446, N38447, N38448, N38449, N38452, N38453, N38454, N38455, N38458, N38459, N38460, N38461, N38462, N38464, N38465, N38467, N38468, N38469, N38470, N38471, N38472, N38473, N38474, N38476, N38478, N38479, N38480, N38482, N38483, N38486, N38487, N38488, N38489, N38493, N38494, N38495, N38496, N38497, N38498, N38501, N38504, N38505, N38506, N38507, N38508, N38509, N38510, N38511, N38512, N38515, N38517, N38518, N38520, N38521, N38522, N38524, N38525, N38527, N38528, N38530, N38531, N38533, N38535, N38536, N38538, N38539, N38540, N38541, N38542, N38544, N38545, N38546, N38547, N38548, N38549, N38550, N38551, N38552, N38553, N38555, N38556, N38557, N38558, N38559, N38561, N38562, N38563, N38567, N38569, N38570, N38571, N38572, N38573, N38574, N38575, N38576, N38577, N38579, N38580, N38582, N38583, N38585, N38586, N38587, N38588, N38589, N38591, N38596, N38597, N38598, N38599, N38602, N38604, N38608, N38609, N38614, N38615, N38616, N38618, N38619, N38620, N38622, N38623, N38627, N38628, N38629, N38630, N38631, N38632, N38633, N38634, N38636, N38637, N38638, N38639, N38643, N38646, N38648, N38650, N38652, N38653, N38654, N38655, N38656, N38657, N38658, N38659, N38660, N38662, N38663, N38664, N38665, N38667, N38668, N38669, N38670, N38671, N38672, N38674, N38675, N38676, N38679, N38680, N38682, N38684, N38686, N38687, N38688, N38689, N38695, N38696, N38697, N38699, N38700, N38704, N38705, N38707, N38708, N38710, N38712, N38713, N38714, N38715, N38717, N38718, N38719, N38720, N38721, N38722, N38723, N38725, N38726, N38728, N38730, N38731, N38733, N38734, N38736, N38737, N38739, N38740, N38741, N38744, N38746, N38747, N38749, N38750, N38751, N38753, N38755, N38756, N38757, N38758, N38759, N38761, N38762, N38764, N38765, N38766, N38767, N38768, N38769, N38770, N38771, N38772, N38775, N38776, N38778, N38779, N38780, N38781, N38782, N38784, N38785, N38786, N38788, N38791, N38792, N38793, N38794, N38795, N38796, N38798, N38801, N38802, N38803, N38805, N38806, N38808, N38812, N38813, N38815, N38817, N38819, N38821, N38823, N38826, N38827, N38829, N38830, N38832, N38834, N38835, N38836, N38838, N38840, N38841, N38842, N38844, N38845, N38849, N38850, N38851, N38853, N38856, N38857, N38858, N38859, N38862, N38865, N38867, N38868, N38869, N38870, N38874, N38876, N38877, N38880, N38882, N38883, N38884, N38885, N38886, N38887, N38888, N38889, N38890, N38891, N38892, N38893, N38895, N38897, N38898, N38901, N38903, N38904, N38905, N38906, N38907, N38910, N38911, N38913, N38914, N38915, N38916, N38917, N38918, N38919, N38920, N38921, N38922, N38923, N38924, N38925, N38926, N38928, N38931, N38932, N38933, N38934, N38937, N38938, N38939, N38940, N38941, N38944, N38946, N38947, N38949, N38950, N38951, N38952, N38953, N38954, N38956, N38957, N38960, N38961, N38962, N38964, N38966, N38967, N38968, N38970, N38971, N38972, N38974, N38976, N38977, N38980, N38984, N38986, N38987, N38990, N38993, N38994, N38999, N39000, N39001, N39002, N39003, N39005, N39007, N39008, N39010, N39011, N39014, N39016, N39017, N39019, N39020, N39021, N39023, N39024, N39025, N39026, N39028, N39029, N39030, N39031, N39033, N39034, N39035, N39036, N39037, N39038, N39041, N39042, N39043, N39044, N39045, N39046, N39047, N39048, N39049, N39050, N39051, N39053, N39054, N39055, N39057, N39059, N39060, N39061, N39062, N39063, N39064, N39065, N39066, N39068, N39069, N39070, N39071, N39073, N39074, N39076, N39077, N39078, N39079, N39081, N39082, N39084, N39086, N39089, N39090, N39091, N39092, N39093, N39097, N39098, N39101, N39102, N39103, N39104, N39105, N39106, N39107, N39108, N39109, N39110, N39111, N39112, N39117, N39119, N39122, N39123, N39124, N39125, N39126, N39128, N39129, N39131, N39132, N39133, N39134, N39135, N39136, N39137, N39139, N39142, N39143, N39144, N39148, N39149, N39151, N39153, N39154, N39155, N39156, N39157, N39160, N39161, N39163, N39164, N39165, N39166, N39168, N39169, N39170, N39171, N39172, N39173, N39175, N39176, N39177, N39178, N39181, N39182, N39184, N39185, N39186, N39187, N39188, N39190, N39194, N39195, N39196, N39197, N39200, N39201, N39203, N39204, N39206, N39208, N39209, N39211, N39213, N39214, N39216, N39217, N39218, N39219, N39220, N39222, N39223, N39224, N39225, N39227, N39228, N39229, N39230, N39233, N39234, N39236, N39238, N39241, N39242, N39243, N39244, N39247, N39248, N39249, N39250, N39251, N39252, N39253, N39255, N39257, N39258, N39260, N39261, N39262, N39267, N39268, N39270, N39271, N39272, N39273, N39274, N39277, N39278, N39281, N39283, N39284, N39285, N39286, N39287, N39289, N39290, N39291, N39293, N39294, N39295, N39297, N39298, N39299, N39301, N39303, N39304, N39305, N39306, N39308, N39310, N39311, N39316, N39318, N39320, N39321, N39322, N39324, N39325, N39327, N39328, N39329, N39330, N39331, N39332, N39334, N39335, N39336, N39337, N39338, N39339, N39340, N39342, N39345, N39347, N39348, N39351, N39352, N39353, N39354, N39357, N39358, N39359, N39360, N39361, N39366, N39368, N39369, N39372, N39373, N39375, N39376, N39378, N39379, N39380, N39383, N39384, N39388, N39389, N39390, N39391, N39393, N39394, N39395, N39396, N39398, N39401, N39403, N39404, N39406, N39407, N39409, N39410, N39411, N39413, N39414, N39417, N39418, N39419, N39420, N39421, N39422, N39423, N39425, N39429, N39431, N39432, N39433, N39436, N39437, N39438, N39439, N39440, N39441, N39442, N39443, N39444, N39445, N39450, N39451, N39452, N39453, N39456, N39459, N39461, N39463, N39465, N39467, N39468, N39472, N39473, N39475, N39477, N39480, N39482, N39484, N39485, N39486, N39487, N39488, N39489, N39490, N39491, N39494, N39496, N39497, N39499, N39500, N39501, N39502, N39503, N39506, N39507, N39508, N39509, N39511, N39512, N39516, N39517, N39519, N39521, N39522, N39524, N39526, N39527, N39528, N39530, N39531, N39533, N39534, N39535, N39536, N39537, N39539, N39540, N39543, N39544, N39545, N39547, N39548, N39551, N39552, N39553, N39554, N39555, N39556, N39557, N39558, N39560, N39561, N39563, N39564, N39565, N39566, N39567, N39568, N39569, N39570, N39571, N39572, N39573, N39574, N39575, N39576, N39578, N39579, N39581, N39582, N39584, N39586, N39587, N39588, N39589, N39591, N39592, N39593, N39595, N39596, N39598, N39602, N39603, N39606, N39608, N39609, N39610, N39611, N39613, N39615, N39616, N39617, N39618, N39621, N39622, N39623, N39624, N39625, N39626, N39627, N39628, N39629, N39631, N39633, N39634, N39635, N39636, N39637, N39638, N39642, N39643, N39645, N39646, N39647, N39649, N39653, N39654, N39656, N39658, N39661, N39662, N39663, N39664, N39666, N39669, N39672, N39674, N39679, N39680, N39681, N39682, N39685, N39686, N39687, N39692, N39695, N39697, N39698, N39699, N39700, N39701, N39702, N39703, N39704, N39706, N39707, N39708, N39709, N39711, N39713, N39714, N39715, N39717, N39718, N39720, N39721, N39722, N39724, N39725, N39726, N39727, N39729, N39730, N39731, N39733, N39734, N39736, N39737, N39740, N39741, N39743, N39745, N39748, N39751, N39754, N39755, N39756, N39757, N39758, N39759, N39760, N39761, N39763, N39765, N39766, N39768, N39770, N39771, N39773, N39776, N39778, N39779, N39781, N39782, N39783, N39786, N39787, N39788, N39789, N39790, N39791, N39792, N39793, N39794, N39795, N39797, N39798, N39800, N39801, N39803, N39804, N39805, N39806, N39808, N39809, N39810, N39811, N39813, N39814, N39815, N39816, N39817, N39818, N39820, N39821, N39822, N39823, N39825, N39827, N39828, N39830, N39831, N39833, N39834, N39837, N39838, N39839, N39841, N39842, N39843, N39846, N39847, N39848, N39849, N39850, N39851, N39852, N39853, N39854, N39855, N39856, N39860, N39862, N39863, N39864, N39865, N39866, N39867, N39868, N39870, N39871, N39872, N39875, N39876, N39877, N39879, N39880, N39882, N39883, N39884, N39885, N39886, N39889, N39890, N39892, N39894, N39895, N39896, N39897, N39899, N39901, N39902, N39904, N39905, N39906, N39907, N39910, N39912, N39913, N39914, N39915, N39917, N39918, N39920, N39921, N39922, N39923, N39924, N39925, N39926, N39927, N39928, N39929, N39930, N39931, N39933, N39935, N39936, N39939, N39940, N39942, N39944, N39946, N39948, N39950, N39951, N39952, N39954, N39955, N39956, N39957, N39959, N39960, N39961, N39962, N39963, N39965, N39966, N39968, N39969, N39972, N39973, N39974, N39975, N39976, N39977, N39978, N39980, N39982, N39984, N39985, N39987, N39988, N39990, N39991, N39992, N39993, N39994, N39995, N39996, N39999, N40001, N40003, N40005, N40006, N40007, N40008, N40009, N40011, N40013, N40014, N40016, N40017, N40019, N40023, N40024, N40027, N40028, N40031, N40032, N40036, N40037, N40038, N40039, N40044, N40046, N40047, N40048, N40051, N40052, N40053, N40054, N40055, N40056, N40057, N40058, N40061, N40062, N40063, N40064, N40066, N40068, N40069, N40070, N40071, N40073, N40074, N40076, N40077, N40078, N40080, N40081, N40082, N40083, N40084, N40085, N40088, N40089, N40090, N40091, N40092, N40094, N40096, N40099, N40101, N40102, N40103, N40104, N40106, N40107, N40108, N40109, N40111, N40112, N40114, N40115, N40116, N40118, N40119, N40120, N40121, N40124, N40125, N40126, N40127, N40128, N40129, N40133, N40134, N40136, N40137, N40138, N40139, N40142, N40143, N40144, N40145, N40147, N40148, N40152, N40153, N40154, N40155, N40156, N40157, N40158, N40159, N40160, N40161, N40164, N40166, N40168, N40169, N40170, N40171, N40172, N40173, N40174, N40176, N40177, N40178, N40179, N40180, N40181, N40188, N40191, N40192, N40196, N40199, N40200, N40201, N40202, N40204, N40205, N40206, N40207, N40208, N40209, N40210, N40211, N40212, N40213, N40214, N40216, N40217, N40218, N40220, N40221, N40222, N40223, N40225, N40227, N40229, N40230, N40231, N40232, N40233, N40234, N40236, N40237, N40238, N40239, N40240, N40242, N40244, N40245, N40247, N40248, N40249, N40250, N40252, N40253, N40254, N40258, N40259, N40260, N40261, N40263, N40267, N40268, N40270, N40272, N40274, N40275, N40276, N40278, N40279, N40280, N40281, N40282, N40284, N40287, N40288, N40289, N40291, N40294, N40296, N40299, N40300, N40301, N40302, N40303, N40306, N40307, N40308, N40309, N40311, N40313, N40314, N40315, N40316, N40318, N40319, N40320, N40321, N40322, N40324, N40325, N40326, N40329, N40330, N40331, N40332, N40333, N40334, N40335, N40336, N40338, N40339, N40341, N40342, N40344, N40345, N40346, N40347, N40348, N40349, N40350, N40351, N40352, N40353, N40354, N40355, N40357, N40358, N40360, N40361, N40362, N40363, N40364, N40365, N40367, N40369, N40370, N40371, N40372, N40373, N40375, N40376, N40377, N40379, N40381, N40382, N40384, N40385, N40386, N40389, N40390, N40392, N40393, N40394, N40396, N40397, N40398, N40399, N40400, N40404, N40405, N40406, N40408, N40409, N40410, N40412, N40413, N40415, N40416, N40417, N40418, N40420, N40421, N40422, N40423, N40424, N40425, N40427, N40428, N40433, N40434, N40435, N40436, N40437, N40438, N40439, N40441, N40443, N40444, N40445, N40446, N40447, N40450, N40452, N40454, N40455, N40456, N40457, N40458, N40459, N40461, N40462, N40464, N40465, N40466, N40467, N40468, N40469, N40470, N40472, N40474, N40477, N40478, N40479, N40481, N40483, N40484, N40486, N40488, N40489, N40490, N40491, N40492, N40493, N40494, N40495, N40497, N40498, N40499, N40500, N40502, N40505, N40506, N40507, N40509, N40510, N40511, N40513, N40514, N40516, N40517, N40518, N40522, N40523, N40525, N40526, N40527, N40528, N40530, N40531, N40533, N40535, N40537, N40542, N40544, N40545, N40546, N40547, N40549, N40550, N40551, N40552, N40553, N40554, N40557, N40558, N40560, N40561, N40562, N40563, N40564, N40565, N40566, N40567, N40568, N40571, N40573, N40574, N40575, N40577, N40578, N40579, N40583, N40585, N40587, N40589, N40590, N40591, N40592, N40594, N40595, N40596, N40598, N40599, N40601, N40602, N40604, N40605, N40607, N40608, N40610, N40612, N40613, N40614, N40615, N40616, N40617, N40618, N40619, N40620, N40621, N40626, N40627, N40630, N40631, N40632, N40633, N40634, N40636, N40637, N40640, N40642, N40645, N40647, N40648, N40649, N40650, N40654, N40655, N40657, N40658, N40659, N40661, N40662, N40664, N40665, N40668, N40670, N40671, N40673, N40675, N40676, N40677, N40678, N40680, N40681, N40682, N40683, N40684, N40685, N40686, N40687, N40688, N40691, N40693, N40694, N40695, N40696, N40697, N40698, N40699, N40700, N40701, N40702, N40708, N40709, N40710, N40711, N40712, N40713, N40714, N40715, N40716, N40719, N40720, N40721, N40722, N40723, N40724, N40728, N40729, N40731, N40732, N40733, N40735, N40736, N40738, N40739, N40740, N40742, N40744, N40746, N40747, N40748, N40749, N40750, N40756, N40757, N40758, N40760, N40761, N40762, N40763, N40766, N40767, N40768, N40769, N40770, N40771, N40772, N40773, N40775, N40776, N40778, N40779, N40780, N40786, N40787, N40788, N40789, N40790, N40791, N40793, N40794, N40795, N40797, N40798, N40801, N40804, N40805, N40809, N40810, N40811, N40813, N40816, N40822, N40823, N40826, N40827, N40828, N40829, N40830, N40831, N40832, N40833, N40834, N40836, N40837, N40838, N40839, N40840, N40841, N40843, N40844, N40845, N40846, N40849, N40850, N40852, N40854, N40855, N40856, N40857, N40858, N40859, N40860, N40861, N40862, N40863, N40865, N40866, N40868, N40869, N40870, N40871, N40872, N40875, N40876, N40878, N40879, N40880, N40886, N40888, N40892, N40893, N40896, N40899, N40902, N40903, N40904, N40905, N40906, N40907, N40908, N40909, N40910, N40911, N40913, N40915, N40917, N40919, N40920, N40922, N40923, N40924, N40926, N40929, N40930, N40931, N40933, N40934, N40935, N40936, N40937, N40939, N40940, N40942, N40944, N40945, N40946, N40947, N40949, N40950, N40954, N40955, N40956, N40957, N40959, N40960, N40961, N40962, N40963, N40965, N40969, N40971, N40973, N40974, N40978, N40979, N40981, N40983, N40984, N40986, N40987, N40989, N40990, N40991, N40993, N40994, N40995, N40997, N40998, N40999, N41000, N41003, N41006, N41008, N41010, N41012, N41013, N41017, N41018, N41020, N41021, N41022, N41023, N41024, N41026, N41027, N41028, N41029, N41031, N41032, N41033, N41034, N41035, N41036, N41037, N41038, N41039, N41041, N41043, N41045, N41046, N41047, N41048, N41049, N41050, N41052, N41053, N41054, N41055, N41057, N41059, N41060, N41062, N41063, N41064, N41065, N41066, N41067, N41068, N41069, N41070, N41071, N41072, N41073, N41074, N41075, N41076, N41078, N41079, N41080, N41081, N41083, N41084, N41085, N41088, N41093, N41094, N41095, N41096, N41097, N41098, N41100, N41101, N41103, N41104, N41105, N41106, N41107, N41108, N41110, N41111, N41114, N41115, N41117, N41119, N41120, N41121, N41122, N41123, N41124, N41127, N41128, N41129, N41130, N41131, N41132, N41134, N41135, N41136, N41138, N41139, N41144, N41145, N41146, N41147, N41148, N41149, N41150, N41151, N41152, N41153, N41154, N41159, N41160, N41161, N41162, N41165, N41166, N41167, N41168, N41170, N41171, N41172, N41173, N41174, N41176, N41178, N41179, N41181, N41182, N41183, N41184, N41185, N41186, N41187, N41189, N41190, N41193, N41194, N41195, N41196, N41199, N41200, N41201, N41202, N41204, N41208, N41209, N41210, N41211, N41212, N41213, N41214, N41215, N41216, N41219, N41220, N41223, N41224, N41225, N41226, N41227, N41228, N41229, N41232, N41234, N41235, N41236, N41237, N41239, N41240, N41242, N41244, N41246, N41247, N41248, N41249, N41250, N41252, N41253, N41255, N41256, N41257, N41259, N41260, N41262, N41263, N41265, N41266, N41267, N41271, N41273, N41276, N41278, N41279, N41280, N41282, N41283, N41284, N41285, N41286, N41287, N41289, N41290, N41293, N41294, N41295, N41296, N41297, N41299, N41300, N41302, N41303, N41304, N41305, N41306, N41309, N41310, N41311, N41312, N41313, N41315, N41316, N41318, N41319, N41321, N41322, N41323, N41324, N41325, N41329, N41330, N41331, N41333, N41334, N41336, N41337, N41339, N41341, N41342, N41343, N41344, N41348, N41349, N41350, N41352, N41353, N41354, N41355, N41356, N41357, N41359, N41360, N41362, N41363, N41364, N41367, N41368, N41369, N41371, N41372, N41373, N41374, N41375, N41376, N41377, N41378, N41379, N41380, N41381, N41382, N41384, N41386, N41387, N41388, N41389, N41390, N41391, N41392, N41393, N41394, N41395, N41397, N41399, N41400, N41401, N41403, N41404, N41405, N41406, N41407, N41409, N41410, N41412, N41414, N41415, N41417, N41418, N41419, N41421, N41424, N41425, N41426, N41428, N41430, N41431, N41432, N41433, N41434, N41435, N41437, N41438, N41439, N41440, N41441, N41443, N41445, N41446, N41450, N41452, N41453, N41456, N41457, N41458, N41459, N41460, N41461, N41462, N41464, N41466, N41467, N41470, N41471, N41473, N41474, N41476, N41479, N41481, N41483, N41484, N41486, N41489, N41490, N41491, N41493, N41494, N41495, N41496, N41497, N41499, N41500, N41504, N41505, N41506, N41511, N41512, N41513, N41514, N41515, N41518, N41519, N41520, N41521, N41522, N41525, N41526, N41527, N41528, N41529, N41530, N41531, N41532, N41536, N41537, N41540, N41541, N41542, N41543, N41544, N41545, N41547, N41549, N41550, N41551, N41552, N41553, N41554, N41555, N41556, N41558, N41559, N41560, N41561, N41562, N41564, N41565, N41566, N41567, N41568, N41569, N41570, N41571, N41572, N41573, N41574, N41575, N41576, N41577, N41578, N41579, N41580, N41582, N41583, N41584, N41586, N41587, N41588, N41589, N41590, N41591, N41593, N41595, N41596, N41597, N41598, N41600, N41601, N41603, N41604, N41606, N41607, N41608, N41609, N41612, N41613, N41616, N41619, N41621, N41622, N41623, N41628, N41632, N41633, N41636, N41638, N41639, N41640, N41642, N41643, N41645, N41646, N41649, N41650, N41651, N41652, N41654, N41655, N41657, N41658, N41659, N41660, N41661, N41662, N41664, N41665, N41666, N41667, N41668, N41669, N41670, N41671, N41673, N41674, N41675, N41679, N41680, N41681, N41685, N41687, N41692, N41695, N41697, N41698, N41699, N41700, N41701, N41707, N41708, N41709, N41710, N41712, N41714, N41715, N41716, N41717, N41720, N41724, N41725, N41726, N41727, N41728, N41731, N41732, N41733, N41736, N41737, N41741, N41743, N41745, N41749, N41750, N41751, N41752, N41753, N41754, N41758, N41759, N41760, N41761, N41763, N41764, N41765, N41766, N41767, N41768, N41769, N41770, N41775, N41776, N41777, N41778, N41781, N41783, N41786, N41787, N41788, N41792, N41793, N41795, N41796, N41797, N41798, N41800, N41802, N41803, N41804, N41805, N41806, N41807, N41810, N41811, N41812, N41813, N41814, N41815, N41818, N41820, N41822, N41823, N41827, N41829, N41830, N41831, N41832, N41833, N41835, N41836, N41837, N41838, N41839, N41840, N41842, N41843, N41844, N41845, N41846, N41848, N41849, N41851, N41856, N41859, N41860, N41861, N41862, N41865, N41866, N41867, N41869, N41871, N41873, N41874, N41875, N41876, N41877, N41878, N41880, N41881, N41882, N41883, N41885, N41887, N41888, N41889, N41890, N41891, N41892, N41893, N41894, N41895, N41896, N41897, N41898, N41899, N41900, N41901, N41902, N41903, N41904, N41906, N41907, N41908, N41910, N41911, N41912, N41915, N41916, N41917, N41918, N41919, N41920, N41921, N41923, N41924, N41927, N41929, N41931, N41932, N41933, N41935, N41936, N41937, N41938, N41941, N41942, N41943, N41944, N41945, N41947, N41948, N41950, N41951, N41952, N41953, N41956, N41957, N41958, N41959, N41960, N41962, N41964, N41965, N41966, N41968, N41969, N41970, N41972, N41973, N41975, N41977, N41979, N41980, N41982, N41983, N41984, N41985, N41986, N41988, N41990, N41991, N41992, N41993, N41994, N41995, N41996, N41998, N42000, N42001, N42002, N42003, N42004, N42005, N42006, N42008, N42011, N42012, N42013, N42014, N42015, N42016, N42018, N42019, N42020, N42022, N42024, N42025, N42026, N42028, N42029, N42030, N42031, N42033, N42035, N42039, N42040, N42041, N42045, N42047, N42051, N42054, N42055, N42056, N42059, N42061, N42062, N42064, N42066, N42068, N42069, N42070, N42071, N42072, N42074, N42076, N42078, N42080, N42082, N42084, N42085, N42086, N42087, N42088, N42089, N42091, N42092, N42094, N42095, N42096, N42097, N42100, N42101, N42103, N42104, N42105, N42106, N42107, N42108, N42109, N42110, N42113, N42114, N42115, N42116, N42118, N42125, N42127, N42128, N42129, N42131, N42132, N42133, N42136, N42138, N42140, N42141, N42142, N42144, N42145, N42146, N42149, N42150, N42151, N42152, N42153, N42154, N42156, N42158, N42160, N42162, N42164, N42168, N42169, N42170, N42174, N42175, N42176, N42177, N42178, N42180, N42181, N42182, N42185, N42186, N42187, N42188, N42189, N42191, N42192, N42194, N42195, N42197, N42198, N42199, N42200, N42201, N42203, N42204, N42206, N42207, N42208, N42209, N42210, N42211, N42212, N42213, N42214, N42217, N42218, N42219, N42220, N42221, N42222, N42224, N42225, N42227, N42229, N42230, N42232, N42233, N42234, N42235, N42237, N42238, N42240, N42241, N42242, N42243, N42245, N42246, N42247, N42248, N42249, N42250, N42252, N42254, N42255, N42256, N42257, N42258, N42259, N42260, N42262, N42263, N42264, N42265, N42267, N42269, N42270, N42271, N42272, N42273, N42276, N42279, N42280, N42281, N42283, N42284, N42286, N42287, N42288, N42290, N42292, N42294, N42295, N42296, N42297, N42299, N42300, N42301, N42302, N42303, N42304, N42305, N42306, N42308, N42310, N42311, N42313, N42315, N42317, N42318, N42320, N42322, N42323, N42326, N42327, N42328, N42330, N42331, N42332, N42336, N42337, N42342, N42343, N42344, N42345, N42350, N42351, N42352, N42353, N42354, N42355, N42356, N42357, N42360, N42362, N42363, N42364, N42365, N42367, N42368, N42369, N42370, N42376, N42378, N42381, N42382, N42384, N42385, N42386, N42388, N42389, N42390, N42392, N42393, N42395, N42397, N42398, N42399, N42400, N42404, N42406, N42407, N42410, N42411, N42412, N42413, N42414, N42415, N42417, N42418, N42420, N42421, N42422, N42423, N42426, N42427, N42428, N42430, N42431, N42432, N42433, N42434, N42436, N42438, N42439, N42440, N42441, N42446, N42448, N42449, N42450, N42451, N42453, N42457, N42458, N42459, N42460, N42461, N42462, N42463, N42464, N42465, N42466, N42468, N42469, N42470, N42471, N42472, N42473, N42475, N42476, N42477, N42480, N42482, N42483, N42484, N42487, N42488, N42491, N42492, N42493, N42494, N42496, N42498, N42499, N42500, N42502, N42503, N42505, N42508, N42512, N42513, N42515, N42516, N42517, N42519, N42522, N42523, N42524, N42527, N42528, N42529, N42531, N42532, N42534, N42535, N42541, N42542, N42545, N42547, N42548, N42549, N42551, N42552, N42553, N42554, N42556, N42559, N42561, N42562, N42563, N42564, N42565, N42569, N42571, N42572, N42573, N42575, N42577, N42578, N42579, N42581, N42582, N42584, N42585, N42586, N42587, N42588, N42589, N42590, N42591, N42592, N42596, N42599, N42601, N42602, N42603, N42605, N42606, N42607, N42609, N42610, N42611, N42612, N42614, N42615, N42616, N42619, N42620, N42622, N42624, N42628, N42629, N42630, N42631, N42632, N42635, N42636, N42638, N42639, N42642, N42645, N42646, N42649, N42650, N42651, N42653, N42655, N42657, N42659, N42662, N42664, N42665, N42667, N42671, N42672, N42673, N42679, N42681, N42682, N42683, N42684, N42685, N42686, N42687, N42688, N42691, N42693, N42698, N42699, N42700, N42701, N42702, N42703, N42704, N42708, N42710, N42711, N42713, N42714, N42717, N42718, N42719, N42721, N42723, N42724, N42725, N42726, N42727, N42729, N42730, N42731, N42732, N42733, N42734, N42737, N42739, N42740, N42741, N42742, N42745, N42746, N42747, N42748, N42753, N42754, N42755, N42756, N42757, N42758, N42760, N42763, N42764, N42765, N42766, N42768, N42769, N42771, N42773, N42774, N42775, N42776, N42777, N42778, N42779, N42780, N42781, N42782, N42784, N42785, N42786, N42787, N42789, N42791, N42794, N42795, N42796, N42797, N42799, N42801, N42802, N42803, N42804, N42805, N42808, N42809, N42810, N42811, N42813, N42814, N42815, N42816, N42817, N42818, N42820, N42821, N42822, N42823, N42824, N42825, N42826, N42830, N42831, N42833, N42837, N42838, N42842, N42843, N42845, N42846, N42847, N42848, N42849, N42850, N42852, N42853, N42854, N42855, N42857, N42859, N42860, N42863, N42864, N42866, N42868, N42869, N42871, N42872, N42874, N42875, N42876, N42880, N42882, N42884, N42885, N42887, N42888, N42889, N42892, N42893, N42894, N42896, N42897, N42898, N42900, N42902, N42903, N42904, N42905, N42906, N42908, N42909, N42910, N42911, N42912, N42913, N42914, N42915, N42917, N42918, N42919, N42920, N42921, N42922, N42923, N42924, N42925, N42926, N42927, N42928, N42929, N42932, N42936, N42938, N42939, N42940, N42941, N42942, N42944, N42946, N42947, N42949, N42950, N42951, N42952, N42953, N42956, N42957, N42958, N42959, N42963, N42964, N42965, N42966, N42969, N42971, N42972, N42973, N42974, N42977, N42979, N42983, N42984, N42985, N42986, N42987, N42988, N42989, N42990, N42991, N42993, N42994, N42995, N42996, N42997, N42999, N43001, N43002, N43003, N43004, N43005, N43006, N43008, N43009, N43010, N43011, N43012, N43013, N43014, N43016, N43018, N43019, N43020, N43021, N43022, N43024, N43026, N43027, N43028, N43029, N43030, N43031, N43033, N43034, N43035, N43036, N43037, N43038, N43039, N43040, N43041, N43042, N43043, N43044, N43047, N43048, N43049, N43050, N43051, N43052, N43054, N43057, N43058, N43059, N43060, N43061, N43062, N43063, N43064, N43065, N43066, N43068, N43069, N43070, N43071, N43072, N43075, N43079, N43080, N43081, N43082, N43083, N43084, N43088, N43089, N43091, N43093, N43094, N43095, N43098, N43105, N43106, N43107, N43108, N43110, N43111, N43112, N43113, N43114, N43115, N43116, N43117, N43118, N43119, N43121, N43122, N43123, N43124, N43125, N43126, N43127, N43130, N43131, N43132, N43134, N43135, N43137, N43139, N43140, N43141, N43142, N43143, N43144, N43145, N43146, N43147, N43148, N43150, N43151, N43152, N43153, N43154, N43156, N43157, N43158, N43159, N43161, N43162, N43163, N43164, N43165, N43166, N43168, N43169, N43170, N43173, N43174, N43175, N43179, N43180, N43181, N43183, N43187, N43188, N43189, N43190, N43191, N43192, N43193, N43194, N43196, N43197, N43200, N43203, N43204, N43206, N43207, N43210, N43211, N43212, N43214, N43215, N43216, N43219, N43222, N43223, N43225, N43226, N43230, N43232, N43233, N43234, N43236, N43237, N43238, N43240, N43241, N43242, N43243, N43244, N43245, N43246, N43247, N43248, N43250, N43252, N43253, N43255, N43256, N43258, N43259, N43260, N43262, N43263, N43266, N43267, N43270, N43274, N43275, N43277, N43279, N43280, N43281, N43283, N43284, N43285, N43287, N43288, N43289, N43290, N43294, N43295, N43297, N43298, N43299, N43300, N43301, N43302, N43305, N43306, N43307, N43308, N43310, N43313, N43316, N43317, N43318, N43319, N43320, N43321, N43322, N43323, N43328, N43332, N43334, N43335, N43336, N43337, N43338, N43339, N43340, N43341, N43342, N43343, N43345, N43348, N43349, N43350, N43351, N43352, N43353, N43354, N43355, N43356, N43357, N43361, N43362, N43364, N43365, N43368, N43369, N43372, N43373, N43374, N43376, N43377, N43378, N43379, N43380, N43381, N43382, N43383, N43384, N43386, N43387, N43388, N43390, N43391, N43392, N43393, N43394, N43397, N43399, N43400, N43401, N43402, N43403, N43404, N43407, N43409, N43411, N43412, N43413, N43414, N43416, N43417, N43418, N43420, N43421, N43422, N43423, N43424, N43425, N43426, N43428, N43430, N43431, N43432, N43433, N43434, N43437, N43438, N43439, N43440, N43442, N43443, N43444, N43446, N43447, N43448, N43449, N43450, N43452, N43455, N43456, N43457, N43458, N43459, N43460, N43461, N43462, N43463, N43465, N43466, N43467, N43468, N43469, N43470, N43472, N43473, N43474, N43476, N43477, N43478, N43479, N43480, N43481, N43482, N43483, N43484, N43485, N43486, N43487, N43488, N43489, N43490, N43491, N43492, N43493, N43494, N43495, N43496, N43497, N43498, N43499, N43500, N43501, N43502, N43503, N43504, N43505, N43506, N43507, N43508, N43509, N43510, N43511, N43512, N43513, N43514, N43515, N43516, N43517, N43518, N43519, N43520, N43521, N43522, N43524, N43525, N43526, N43527, N43528, N43529, N43530, N43531, N43532, N43533, N43535, N43536, N43537, N43538, N43540, N43541, N43542, N43544, N43545, N43546, N43547, N43548, N43549, N43550, N43551, N43552, N43553, N43555, N43556, N43558, N43560, N43562, N43563, N43565, N43566, N43567, N43568, N43569, N43570, N43571, N43572, N43573, N43574, N43576, N43577, N43578, N43579, N43580, N43581, N43583, N43584, N43586, N43587, N43588, N43589, N43590, N43591, N43592, N43594, N43595, N43596, N43597, N43598, N43599, N43600, N43601, N43602, N43603, N43604, N43605, N43606, N43607, N43608, N43609, N43610, N43611, N43612, N43613, N43614, N43615, N43616, N43617, N43618, N43619, N43621, N43622, N43623, N43624, N43625, N43626, N43628, N43629, N43630, N43632, N43634, N43635, N43636, N43637, N43638, N43639, N43640, N43641, N43642, N43644, N43645, N43646, N43647, N43648, N43649, N43650, N43651, N43652, N43653, N43654, N43655, N43656, N43657, N43658, N43659, N43660, N43661, N43662, N43663, N43664, N43665, N43666, N43667, N43668, N43669, N43670, N43671, N43672, N43673, N43674, N43676, N43677, N43678, N43679, N43680, N43681, N43682, N43683, N43684, N43685, N43686, N43687, N43688, N43689, N43691, N43692, N43693, N43694, N43695, N43696, N43697, N43698, N43699, N43700, N43701, N43702, N43704, N43705, N43706, N43707, N43708, N43709, N43710, N43711, N43712, N43713, N43714, N43715, N43716, N43717, N43718, N43719, N43720, N43721, N43722, N43723, N43724, N43725, N43726, N43727, N43728, N43730, N43731, N43732, N43733, N43734, N43735, N43736, N43737, N43738, N43739, N43740, N43741, N43742, N43743, N43744, N43745, N43746, N43748, N43749, N43750, N43751, N43752, N43753, N43754, N43755, N43756, N43757, N43758, N43759, N43761, N43763, N43765, N43766, N43767, N43768, N43769, N43772, N43773, N43774, N43775, N43777, N43778, N43779, N43780, N43781, N43782, N43783, N43784, N43785, N43786, N43787, N43788, N43789, N43790, N43791, N43792, N43793, N43794, N43795, N43797, N43798, N43799, N43800, N43801, N43802, N43804, N43805, N43806, N43807, N43808, N43809, N43810, N43811, N43812, N43813, N43814, N43815, N43816, N43817, N43818, N43819, N43820, N43821, N43822, N43823, N43824, N43825, N43826, N43827, N43828, N43829, N43830, N43831, N43832, N43833, N43834, N43835, N43836, N43837, N43838, N43839, N43840, N43841, N43842, N43843, N43845, N43846, N43847, N43848, N43849, N43850, N43851, N43852, N43853, N43854, N43855, N43856, N43857, N43859, N43860, N43861, N43862, N43863, N43864, N43865, N43866, N43867, N43868, N43869, N43870, N43871, N43872, N43873, N43874, N43875, N43876, N43877, N43879, N43880, N43881, N43882, N43883, N43884, N43885, N43886, N43887, N43888, N43889, N43891, N43892, N43893, N43894, N43895, N43896, N43897, N43898, N43900, N43901, N43902, N43903, N43904, N43905, N43906, N43907, N43908, N43909, N43910, N43911, N43912, N43913, N43914, N43915, N43916, N43917, N43918, N43919, N43921, N43922, N43923, N43924, N43925, N43926, N43927, N43928, N43929, N43930, N43931, N43932, N43934, N43935, N43936, N43937, N43938, N43939, N43942, N43943, N43944, N43945, N43946, N43947, N43948, N43949, N43950, N43951, N43952, N43953, N43955, N43956, N43957, N43958, N43959, N43960, N43961, N43962, N43964, N43965, N43966, N43967, N43968, N43969, N43970, N43971, N43972, N43973, N43974, N43975, N43976, N43977, N43978, N43979, N43980, N43981, N43982, N43983, N43984, N43985, N43986, N43987, N43988, N43989, N43990, N43991, N43992, N43994, N43995, N43996, N43997, N43999, N44000, N44001, N44002, N44003, N44004, N44005, N44007, N44008, N44009, N44010, N44011, N44012, N44013, N44014, N44015, N44016, N44017, N44018, N44019, N44020, N44021, N44022, N44023, N44024, N44025, N44026, N44027, N44028, N44029, N44030, N44031, N44032, N44033, N44034, N44035, N44036, N44037, N44038, N44039, N44040, N44041, N44042, N44043, N44044, N44045, N44046, N44047, N44048, N44049, N44050, N44051, N44052, N44053, N44055, N44056, N44057, N44058, N44059, N44060, N44061, N44062, N44063, N44064, N44065, N44066, N44067, N44069, N44070, N44071, N44072, N44073, N44074, N44075, N44076, N44077, N44078, N44079, N44080, N44081, N44082, N44083, N44084, N44085, N44086, N44087, N44088, N44089, N44090, N44091, N44092, N44093, N44094, N44095, N44097, N44098, N44099, N44100, N44101, N44102, N44103, N44105, N44106, N44107, N44108, N44109, N44110, N44111, N44112, N44113, N44114, N44115, N44116, N44117, N44118, N44119, N44121, N44122, N44123, N44124, N44125, N44126, N44127, N44128, N44129, N44130, N44131, N44132, N44133, N44135, N44136, N44137, N44139, N44141, N44142, N44143, N44144, N44145, N44146, N44147, N44148, N44149, N44150, N44151, N44152, N44153, N44154, N44155, N44156, N44158, N44159, N44160, N44161, N44162, N44163, N44164, N44165, N44166, N44167, N44168, N44169, N44171, N44172, N44174, N44175, N44177, N44178, N44181, N44182, N44183, N44184, N44185, N44186, N44187, N44188, N44189, N44190, N44191, N44192, N44193, N44194, N44195, N44196, N44197, N44198, N44199, N44200, N44201, N44202, N44203, N44204, N44205, N44206, N44207, N44208, N44209, N44210, N44212, N44213, N44215, N44216, N44217, N44218, N44219, N44220, N44221, N44222, N44224, N44225, N44226, N44227, N44229, N44230, N44232, N44233, N44234, N44235, N44236, N44237, N44238, N44239, N44240, N44241, N44242, N44243, N44244, N44246, N44248, N44249, N44250, N44251, N44252, N44254, N44255, N44256, N44257, N44258, N44259, N44261, N44262, N44263, N44264, N44265, N44266, N44267, N44268, N44269, N44271, N44272, N44273, N44274, N44275, N44276, N44277, N44278, N44279, N44281, N44282, N44283, N44284, N44285, N44286, N44288, N44289, N44290, N44291, N44292, N44293, N44294, N44295, N44296, N44297, N44298, N44299, N44300, N44301, N44302, N44303, N44304, N44305, N44306, N44307, N44308, N44309, N44310, N44311, N44312, N44313, N44314, N44316, N44317, N44318, N44319, N44320, N44321, N44322, N44323, N44324, N44325, N44326, N44327, N44328, N44329, N44330, N44331, N44332, N44333, N44334, N44335, N44338, N44339, N44341, N44342, N44343, N44345, N44346, N44347, N44348, N44349, N44350, N44352, N44353, N44354, N44355, N44356, N44357, N44359, N44360, N44363, N44364, N44365, N44366, N44367, N44368, N44369, N44370, N44371, N44372, N44373, N44375, N44376, N44377, N44378, N44379, N44380, N44381, N44384, N44385, N44386, N44387, N44388, N44389, N44390, N44391, N44392, N44393, N44394, N44395, N44396, N44397, N44399, N44400, N44401, N44402, N44403, N44404, N44405, N44406, N44407, N44408, N44409, N44410, N44411, N44412, N44413, N44414, N44415, N44416, N44417, N44418, N44419, N44420, N44421, N44422, N44423, N44424, N44425, N44426, N44427, N44428, N44429, N44430, N44431, N44432, N44433, N44434, N44435, N44436, N44437, N44438, N44440, N44441, N44442, N44443, N44444, N44445, N44446, N44447, N44448, N44450, N44451, N44452, N44453, N44456, N44457, N44458, N44459, N44461, N44462, N44463, N44464, N44465, N44466, N44467, N44469, N44470, N44471, N44472, N44473, N44474, N44475, N44476, N44478, N44479, N44480, N44481, N44482, N44483, N44484, N44486, N44488, N44489, N44491, N44492, N44493, N44494, N44495, N44496, N44497, N44498, N44499, N44500, N44502, N44503, N44504, N44505, N44506, N44507, N44508, N44509, N44510, N44511, N44512, N44513, N44514, N44515, N44516, N44517, N44518, N44519, N44520, N44521, N44522, N44523, N44525, N44526, N44527, N44528, N44529, N44530, N44531, N44532, N44533, N44534, N44536, N44537, N44538, N44539, N44540, N44541, N44543, N44544, N44545, N44547, N44548, N44549, N44550, N44551, N44552, N44553, N44554, N44555, N44556, N44557, N44558, N44559, N44560, N44561, N44562, N44563, N44564, N44566, N44567, N44568, N44569, N44570, N44572, N44573, N44574, N44575, N44576, N44577, N44578, N44579, N44580, N44581, N44582, N44583, N44585, N44586, N44587, N44588, N44589, N44590, N44592, N44593, N44594, N44595, N44596, N44597, N44598, N44599, N44600, N44601, N44602, N44604, N44605, N44606, N44607, N44608, N44609, N44610, N44611, N44612, N44613, N44614, N44615, N44616, N44617, N44618, N44619, N44620, N44621, N44622, N44625, N44626, N44627, N44628, N44629, N44630, N44631, N44632, N44633, N44634, N44635, N44636, N44637, N44638, N44639, N44641, N44643, N44644, N44645, N44646, N44647, N44648, N44649, N44650, N44651, N44652, N44653, N44654, N44655, N44656, N44657, N44658, N44659, N44660, N44661, N44662, N44664, N44666, N44667, N44668, N44669, N44670, N44671, N44672, N44673, N44674, N44675, N44676, N44677, N44678, N44679, N44680, N44681, N44682, N44683, N44684, N44685, N44686, N44687, N44688, N44689, N44690, N44691, N44692, N44693, N44694, N44695, N44696, N44698, N44699, N44700, N44701, N44702, N44704, N44705, N44706, N44707, N44709, N44711, N44712, N44713, N44714, N44715, N44716, N44717, N44718, N44719, N44722, N44723, N44724, N44725, N44726, N44728, N44729, N44730, N44732, N44733, N44734, N44735, N44736, N44737, N44738, N44739, N44740, N44741, N44742, N44743, N44744, N44745, N44746, N44748, N44749, N44750, N44751, N44752, N44753, N44754, N44755, N44756, N44757, N44758, N44759, N44760, N44761, N44762, N44763, N44764, N44768, N44769, N44770, N44771, N44772, N44773, N44774, N44775, N44776, N44777, N44778, N44779, N44780, N44781, N44782, N44783, N44784, N44785, N44786, N44787, N44788, N44789, N44791, N44792, N44793, N44795, N44797, N44798, N44799, N44801, N44802, N44803, N44804, N44805, N44806, N44807, N44808, N44809, N44810, N44811, N44812, N44813, N44814, N44815, N44816, N44817, N44818, N44819, N44820, N44821, N44823, N44824, N44825, N44826, N44827, N44828, N44829, N44830, N44831, N44832, N44833, N44835, N44836, N44837, N44838, N44839, N44840, N44841, N44842, N44843, N44844, N44845, N44846, N44847, N44848, N44850, N44851, N44852, N44853, N44854, N44855, N44856, N44857, N44858, N44859, N44860, N44861, N44862, N44863, N44864, N44865, N44866, N44867, N44868, N44869, N44870, N44871, N44872, N44873, N44874, N44875, N44876, N44877, N44878, N44879, N44880, N44881, N44882, N44883, N44884, N44885, N44886, N44888, N44889, N44890, N44891, N44893, N44894, N44896, N44897, N44898, N44899, N44900, N44901, N44902, N44903, N44904, N44905, N44906, N44907, N44908, N44909, N44910, N44911, N44912, N44913, N44914, N44915, N44916, N44917, N44918, N44919, N44920, N44921, N44922, N44923, N44924, N44925, N44926, N44927, N44928, N44929, N44930, N44931, N44932, N44933, N44934, N44935, N44936, N44938, N44939, N44940, N44941, N44942, N44943, N44945, N44946, N44947, N44948, N44949, N44950, N44952, N44953, N44954, N44955, N44956, N44957, N44958, N44959, N44960, N44961, N44962, N44963, N44964, N44965, N44966, N44968, N44969, N44971, N44972, N44973, N44974, N44976, N44977, N44978, N44979, N44980, N44981, N44982, N44983, N44984, N44985, N44986, N44989, N44990, N44991, N44992, N44993, N44994, N44995, N44996, N44997, N44998, N44999, N45000, N45001, N45002, N45003, N45004, N45005, N45006, N45007, N45008, N45009, N45010, N45011, N45012, N45013, N45014, N45015, N45016, N45017, N45018, N45020, N45021, N45022, N45023, N45024, N45025, N45026, N45027, N45028, N45029, N45030, N45031, N45032, N45033, N45034, N45036, N45037, N45038, N45039, N45040, N45041, N45042, N45043, N45044, N45045, N45046, N45047, N45048, N45050, N45051, N45052, N45053, N45054, N45055, N45056, N45057, N45058, N45059, N45060, N45061, N45063, N45064, N45065, N45066, N45067, N45068, N45069, N45070, N45071, N45072, N45073, N45074, N45075, N45076, N45078, N45079, N45080, N45081, N45082, N45084, N45085, N45086, N45087, N45088, N45089, N45090, N45091, N45092, N45093, N45094, N45095, N45096, N45097, N45098, N45099, N45100, N45101, N45102, N45103, N45105, N45106, N45107, N45108, N45109, N45110, N45111, N45113, N45114, N45115, N45116, N45117, N45118, N45119, N45120, N45121, N45122, N45123, N45124, N45125, N45127, N45128, N45129, N45130, N45131, N45132, N45133, N45135, N45136, N45138, N45139, N45142, N45143, N45144, N45145, N45146, N45147, N45148, N45149, N45150, N45151, N45153, N45154, N45155, N45157, N45158, N45159, N45160, N45161, N45162, N45163, N45164, N45165, N45166, N45167, N45168, N45169, N45170, N45171, N45172, N45173, N45174, N45175, N45176, N45178, N45179, N45180, N45181, N45182, N45183, N45185, N45186, N45187, N45188, N45189, N45190, N45191, N45192, N45193, N45194, N45195, N45196, N45197, N45198, N45199, N45200, N45201, N45202, N45203, N45205, N45206, N45208, N45209, N45210, N45212, N45213, N45214, N45215, N45216, N45217, N45219, N45220, N45221, N45222, N45223, N45224, N45225, N45227, N45228, N45229, N45230, N45231, N45232, N45233, N45234, N45235, N45236, N45237, N45238, N45242, N45243, N45244, N45245, N45246, N45247, N45248, N45249, N45250, N45251, N45252, N45253, N45254, N45255, N45256, N45257, N45258, N45259, N45260, N45261, N45262, N45263, N45267, N45269, N45270, N45271, N45272, N45273, N45274, N45275, N45276, N45277, N45278, N45279, N45280, N45281, N45282, N45283, N45284, N45285, N45286, N45287, N45288, N45289, N45290, N45291, N45292, N45293, N45294, N45295, N45296, N45297, N45298, N45299, N45300, N45301, N45303, N45304, N45305, N45307, N45308, N45309, N45310, N45311, N45312, N45313, N45314, N45316, N45317, N45318, N45319, N45320, N45321, N45322, N45323, N45324, N45325, N45326, N45327, N45328, N45329, N45330, N45331, N45332, N45333, N45335, N45336, N45337, N45338, N45339, N45340, N45341, N45342, N45343, N45344, N45345, N45346, N45347, N45348, N45349, N45352, N45353, N45354, N45355, N45356, N45357, N45358, N45359, N45360, N45361, N45362, N45363, N45364, N45365, N45366, N45367, N45369, N45370, N45372, N45373, N45374, N45375, N45376, N45377, N45378, N45379, N45380, N45381, N45382, N45383, N45384, N45385, N45386, N45387, N45388, N45389, N45390, N45391, N45393, N45394, N45395, N45396, N45397, N45398, N45399, N45402, N45403, N45405, N45406, N45407, N45408, N45409, N45410, N45411, N45412, N45413, N45414, N45415, N45416, N45417, N45418, N45419, N45420, N45421, N45422, N45423, N45424, N45425, N45426, N45427, N45429, N45430, N45431, N45433, N45434, N45435, N45436, N45438, N45439, N45440, N45441, N45442, N45443, N45444, N45445, N45447, N45448, N45449, N45450, N45451, N45452, N45458, N45459, N45460, N45461, N45462, N45464, N45465, N45466, N45467, N45468, N45469, N45471, N45472, N45473, N45474, N45475, N45476, N45477, N45478, N45479, N45480, N45481, N45483, N45484, N45485, N45486, N45487, N45488, N45489, N45490, N45491, N45492, N45493, N45494, N45495, N45496, N45497, N45498, N45499, N45500, N45501, N45502, N45503, N45504, N45505, N45506, N45507, N45508, N45509, N45511, N45513, N45514, N45515, N45516, N45517, N45518, N45519, N45520, N45521, N45522, N45523, N45524, N45525, N45526, N45527, N45530, N45531, N45532, N45533, N45535, N45536, N45537, N45538, N45539, N45540, N45541, N45542, N45543, N45544, N45545, N45547, N45548, N45549, N45550, N45551, N45552, N45553, N45554, N45555, N45556, N45557, N45558, N45559, N45561, N45562, N45563, N45564, N45566, N45567, N45568, N45569, N45570, N45571, N45572, N45573, N45574, N45575, N45576, N45577, N45578, N45579, N45580, N45581, N45584, N45585, N45586, N45587, N45588, N45589, N45590, N45592, N45593, N45595, N45597, N45599, N45600, N45601, N45602, N45603, N45605, N45606, N45607, N45608, N45609, N45610, N45611, N45612, N45613, N45614, N45615, N45616, N45617, N45618, N45619, N45620, N45621, N45622, N45623, N45625, N45627, N45628, N45629, N45630, N45631, N45633, N45634, N45635, N45636, N45637, N45638, N45639, N45640, N45641, N45642, N45643, N45646, N45647, N45648, N45649, N45650, N45652, N45653, N45654, N45655, N45656, N45657, N45658, N45659, N45660, N45661, N45662, N45663, N45664, N45665, N45666, N45667, N45669, N45671, N45673, N45674, N45676, N45677, N45678, N45679, N45680, N45681, N45682, N45683, N45685, N45686, N45687, N45688, N45689, N45690, N45691, N45692, N45693, N45694, N45695, N45696, N45697, N45698, N45699, N45701, N45702, N45703, N45705, N45706, N45707, N45708, N45709, N45710, N45711, N45712, N45713, N45714, N45716, N45717, N45718, N45719, N45720, N45721, N45722, N45723, N45724, N45725, N45726, N45727, N45728, N45729, N45730, N45732, N45733, N45735, N45736, N45737, N45739, N45740, N45741, N45742, N45743, N45744, N45745, N45746, N45747, N45748, N45749, N45750, N45751, N45752, N45753, N45754, N45756, N45757, N45758, N45759, N45760, N45761, N45762, N45763, N45764, N45765, N45766, N45768, N45769, N45770, N45771, N45772, N45773, N45774, N45775, N45776, N45778, N45779, N45780, N45782, N45783, N45784, N45786, N45787, N45789, N45790, N45791, N45792, N45793, N45795, N45796, N45797, N45798, N45799, N45800, N45801, N45802, N45803, N45804, N45805, N45806, N45807, N45808, N45809, N45810, N45811, N45812, N45813, N45814, N45815, N45816, N45817, N45818, N45819, N45820, N45821, N45822, N45823, N45824, N45825, N45826, N45827, N45828, N45829, N45830, N45831, N45833, N45834, N45835, N45836, N45837, N45838, N45839, N45840, N45841, N45842, N45843, N45844, N45845, N45846, N45847, N45848, N45849, N45850, N45851, N45852, N45853, N45854, N45855, N45856, N45857, N45858, N45859, N45860, N45861, N45862, N45863, N45865, N45866, N45867, N45868, N45869, N45870, N45871, N45872, N45873, N45874, N45875, N45876, N45877, N45878, N45879, N45880, N45881, N45882, N45883, N45884, N45885, N45886, N45887, N45888, N45889, N45890, N45891, N45892, N45893, N45894, N45895, N45896, N45897, N45898, N45899, N45901, N45902, N45903, N45904, N45905, N45906, N45907, N45908, N45909, N45910, N45911, N45912, N45913, N45914, N45915, N45916, N45917, N45918, N45919, N45920, N45921, N45922, N45923, N45924, N45925, N45926, N45927, N45928, N45929, N45930, N45931, N45932, N45933, N45934, N45935, N45936, N45938, N45939, N45940, N45941, N45942, N45944, N45945, N45946, N45947, N45948, N45949, N45950, N45951, N45952, N45953, N45954, N45955, N45956, N45957, N45958, N45960, N45961, N45962, N45963, N45964, N45965, N45966, N45967, N45968, N45969, N45971, N45972, N45973, N45974, N45975, N45976, N45979, N45980, N45981, N45983, N45984, N45985, N45986, N45987, N45988, N45989, N45990, N45991, N45992, N45993, N45994, N45995, N45996, N45997, N45999, N46000, N46002, N46003, N46004, N46005, N46006, N46007, N46008, N46011, N46012, N46013, N46014, N46015, N46016, N46017, N46018, N46019, N46020, N46021, N46022, N46023, N46024, N46025, N46026, N46027, N46028, N46029, N46030, N46031, N46032, N46034, N46035, N46036, N46037, N46038, N46039, N46040, N46041, N46042, N46043, N46044, N46045, N46047, N46048, N46049, N46051, N46052, N46053, N46054, N46056, N46057, N46058, N46059, N46060, N46061, N46063, N46064, N46065, N46066, N46067, N46068, N46069, N46070, N46071, N46072, N46073, N46074, N46075, N46077, N46078, N46079, N46080, N46081, N46082, N46085, N46086, N46087, N46089, N46090, N46091, N46092, N46093, N46094, N46095, N46096, N46097, N46098, N46099, N46100, N46101, N46102, N46103, N46104, N46105, N46106, N46107, N46108, N46109, N46110, N46111, N46112, N46113, N46114, N46115, N46116, N46117, N46118, N46121, N46122, N46123, N46124, N46125, N46126, N46127, N46128, N46129, N46131, N46132, N46133, N46134, N46135, N46136, N46137, N46139, N46140, N46141, N46142, N46143, N46144, N46145, N46146, N46147, N46148, N46149, N46150, N46151, N46152, N46153, N46154, N46155, N46156, N46157, N46158, N46159, N46160, N46161, N46162, N46163, N46164, N46166, N46167, N46168, N46169, N46170, N46171, N46172, N46173, N46174, N46175, N46176, N46177, N46178, N46179, N46180, N46181, N46182, N46183, N46184, N46185, N46186, N46187, N46188, N46190, N46191, N46192, N46193, N46194, N46195, N46196, N46197, N46198, N46200, N46201, N46202, N46203, N46204, N46205, N46206, N46207, N46208, N46209, N46210, N46211, N46212, N46213, N46214, N46215, N46216, N46217, N46218, N46219, N46220, N46221, N46222, N46223, N46226, N46227, N46228, N46229, N46230, N46231, N46232, N46233, N46234, N46235, N46236, N46237, N46238, N46239, N46241, N46242, N46243, N46244, N46245, N46246, N46247, N46248, N46249, N46251, N46252, N46253, N46254, N46255, N46256, N46257, N46258, N46260, N46261, N46262, N46263, N46264, N46265, N46267, N46268, N46269, N46270, N46271, N46272, N46273, N46274, N46275, N46276, N46277, N46278, N46280, N46281, N46282, N46283, N46284, N46285, N46286, N46288, N46289, N46290, N46291, N46292, N46293, N46295, N46296, N46297, N46298, N46299, N46302, N46303, N46304, N46305, N46306, N46307, N46309, N46310, N46311, N46312, N46314, N46315, N46316, N46317, N46318, N46319, N46320, N46321, N46322, N46323, N46324, N46325, N46326, N46327, N46328, N46329, N46330, N46331, N46332, N46333, N46336, N46337, N46338, N46339, N46340, N46341, N46342, N46343, N46344, N46345, N46346, N46347, N46348, N46349, N46350, N46351, N46352, N46353, N46354, N46355, N46356, N46357, N46358, N46359, N46360, N46361, N46362, N46365, N46366, N46367, N46368, N46369, N46370, N46371, N46372, N46373, N46374, N46375, N46376, N46377, N46378, N46379, N46380, N46381, N46382, N46384, N46385, N46387, N46388, N46389, N46391, N46393, N46394, N46395, N46396, N46397, N46398, N46399, N46400, N46401, N46402, N46403, N46404, N46405, N46406, N46407, N46408, N46409, N46410, N46411, N46412, N46413, N46414, N46415, N46416, N46417, N46419, N46420, N46421, N46422, N46423, N46424, N46425, N46426, N46428, N46429, N46430, N46431, N46432, N46433, N46434, N46435, N46436, N46437, N46438, N46439, N46440, N46441, N46442, N46443, N46444, N46445, N46446, N46447, N46448, N46449, N46450, N46451, N46452, N46453, N46454, N46455, N46456, N46457, N46459, N46460, N46461, N46462, N46463, N46464, N46465, N46466, N46467, N46468, N46469, N46470, N46471, N46472, N46473, N46474, N46475, N46476, N46477, N46478, N46479, N46480, N46481, N46483, N46484, N46485, N46486, N46487, N46489, N46490, N46491, N46492, N46493, N46494, N46495, N46496, N46497, N46498, N46499, N46500, N46501, N46503, N46505, N46506, N46507, N46508, N46509, N46510, N46511, N46512, N46513, N46514, N46515, N46517, N46518, N46519, N46520, N46521, N46523, N46524, N46525, N46526, N46527, N46528, N46529, N46530, N46531, N46532, N46533, N46534, N46536, N46537, N46538, N46539, N46540, N46541, N46542, N46543, N46544, N46545, N46546, N46547, N46548, N46549, N46550, N46551, N46552, N46553, N46554, N46555, N46556, N46557, N46558, N46559, N46560, N46561, N46562, N46563, N46564, N46565, N46566, N46567, N46568, N46569, N46570, N46571, N46572, N46573, N46574, N46575, N46576, N46577, N46578, N46579, N46580, N46581, N46582, N46583, N46584, N46585, N46586, N46587, N46588, N46589, N46590, N46591, N46592, N46593, N46594, N46596, N46597, N46598, N46599, N46601, N46602, N46603, N46604, N46605, N46606, N46608, N46609, N46610, N46611, N46612, N46613, N46614, N46615, N46616, N46617, N46618, N46619, N46620, N46621, N46622, N46623, N46624, N46625, N46626, N46627, N46628, N46629, N46631, N46632, N46633, N46634, N46635, N46636, N46637, N46638, N46639, N46640, N46641, N46642, N46643, N46644, N46645, N46646, N46647, N46648, N46649, N46650, N46651, N46653, N46654, N46655, N46656, N46657, N46658, N46659, N46660, N46661, N46662, N46664, N46665, N46666, N46667, N46668, N46669, N46671, N46672, N46673, N46674, N46675, N46676, N46677, N46678, N46679, N46680, N46681, N46682, N46683, N46684, N46685, N46686, N46687, N46688, N46689, N46690, N46691, N46692, N46693, N46694, N46695, N46696, N46697, N46699, N46700, N46701, N46702, N46703, N46704, N46705, N46707, N46708, N46709, N46710, N46712, N46713, N46714, N46715, N46716, N46717, N46718, N46719, N46720, N46721, N46722, N46723, N46725, N46726, N46727, N46728, N46729, N46730, N46731, N46732, N46733, N46734, N46735, N46736, N46737, N46738, N46740, N46741, N46742, N46743, N46744, N46745, N46746, N46747, N46748, N46749, N46750, N46751, N46752, N46753, N46754, N46756, N46757, N46758, N46759, N46760, N46761, N46762, N46763, N46764, N46765, N46766, N46767, N46768, N46769, N46772, N46773, N46774, N46775, N46776, N46777, N46778, N46779, N46780, N46781, N46782, N46783, N46784, N46785, N46786, N46787, N46788, N46790, N46791, N46792, N46793, N46794, N46795, N46796, N46797, N46798, N46799, N46800, N46801, N46802, N46803, N46804, N46805, N46806, N46807, N46808, N46809, N46810, N46812, N46813, N46814, N46815, N46816, N46817, N46818, N46819, N46820, N46821, N46822, N46823, N46824, N46825, N46826, N46827, N46828, N46829, N46830, N46832, N46833, N46834, N46835, N46836, N46837, N46838, N46839, N46840, N46841, N46843, N46844, N46845, N46846, N46847, N46848, N46850, N46851, N46852, N46853, N46854, N46855, N46856, N46857, N46859, N46860, N46862, N46863, N46864, N46865, N46866, N46867, N46868, N46869, N46870, N46871, N46872, N46873, N46874, N46875, N46876, N46877, N46878, N46879, N46880, N46881, N46882, N46883, N46884, N46885, N46886, N46887, N46888, N46889, N46890, N46891, N46892, N46893, N46894, N46895, N46896, N46897, N46898, N46899, N46900, N46902, N46903, N46904, N46905, N46906, N46907, N46908, N46909, N46910, N46911, N46912, N46913, N46914, N46915, N46916, N46917, N46918, N46919, N46920, N46921, N46922, N46923, N46924, N46925, N46926, N46928, N46929, N46931, N46932, N46933, N46934, N46935, N46936, N46937, N46939, N46940, N46941, N46942, N46945, N46946, N46947, N46948, N46949, N46950, N46951, N46952, N46953, N46954, N46955, N46956, N46957, N46958, N46959, N46960, N46961, N46962, N46963, N46964, N46965, N46966, N46967, N46968, N46969, N46970, N46971, N46972, N46973, N46975, N46976, N46977, N46978, N46979, N46980, N46981, N46982, N46983, N46984, N46985, N46987, N46988, N46989, N46990, N46991, N46992, N46993, N46994, N46995, N46997, N46998, N46999, N47001, N47002, N47003, N47004, N47005, N47006, N47007, N47008, N47009, N47010, N47011, N47012, N47013, N47014, N47015, N47016, N47017, N47018, N47019, N47020, N47021, N47023, N47024, N47025, N47026, N47027, N47028, N47029, N47030, N47031, N47032, N47034, N47035, N47036, N47037, N47038, N47039, N47040, N47041, N47042, N47043, N47044, N47045, N47046, N47047, N47048, N47049, N47050, N47051, N47052, N47053, N47054, N47055, N47056, N47058, N47059, N47060, N47061, N47062, N47063, N47064, N47065, N47066, N47067, N47068, N47069, N47070, N47071, N47072, N47073, N47074, N47075, N47076, N47077, N47078, N47079, N47080, N47081, N47082, N47083, N47084, N47086, N47087, N47088, N47089, N47090, N47091, N47092, N47093, N47094, N47095, N47096, N47097, N47098, N47099, N47100, N47101, N47102, N47103, N47104, N47105, N47106, N47107, N47108, N47109, N47110, N47111, N47112, N47113, N47115, N47116, N47118, N47119, N47120, N47121, N47122, N47123, N47124, N47125, N47127, N47128, N47129, N47130, N47131, N47133, N47134, N47135, N47136, N47137, N47138, N47139, N47141, N47142, N47143, N47145, N47146, N47147, N47148, N47149, N47150, N47151, N47152, N47153, N47155, N47156, N47157, N47158, N47159, N47160, N47161, N47162, N47163, N47164, N47165, N47166, N47167, N47168, N47170, N47171, N47172, N47173, N47174, N47175, N47176, N47177, N47178, N47179, N47180, N47181, N47182, N47184, N47185, N47186, N47187, N47188, N47189, N47190, N47191, N47192, N47193, N47196, N47197, N47198, N47199, N47200, N47201, N47202, N47203, N47204, N47205, N47206, N47207, N47208, N47209, N47210, N47211, N47212, N47213, N47214, N47215, N47216, N47217, N47219, N47220, N47221, N47222, N47223, N47224, N47225, N47226, N47227, N47228, N47229, N47230, N47231, N47232, N47234, N47235, N47236, N47237, N47238, N47239, N47240, N47241, N47242, N47243, N47244, N47246, N47247, N47248, N47249, N47250, N47251, N47252, N47253, N47254, N47255, N47256, N47257, N47258, N47259, N47260, N47261, N47262, N47263, N47264, N47266, N47267, N47268, N47269, N47270, N47271, N47272, N47273, N47274, N47275, N47276, N47277, N47278, N47279, N47280, N47281, N47282, N47283, N47284, N47285, N47286, N47287, N47288, N47289, N47290, N47291, N47292, N47293, N47294, N47295, N47296, N47297, N47298, N47299, N47300, N47301, N47302, N47303, N47304, N47305, N47306, N47307, N47308, N47309, N47310, N47311, N47312, N47313, N47314, N47315, N47316, N47317, N47318, N47319, N47320, N47321, N47322, N47323, N47324, N47325, N47326, N47327, N47328, N47329, N47330, N47331, N47332, N47335, N47336, N47337, N47338, N47339, N47340, N47341, N47342, N47343, N47344, N47345, N47346, N47347, N47348, N47349, N47350, N47351, N47352, N47353, N47354, N47355, N47356, N47357, N47358, N47359, N47360, N47361, N47362, N47363, N47364, N47365, N47366, N47367, N47368, N47369, N47370, N47371, N47372, N47373, N47374, N47376, N47378, N47379, N47380, N47381, N47382, N47383, N47384, N47385, N47386, N47387, N47388, N47389, N47390, N47391, N47392, N47393, N47394, N47395, N47396, N47397, N47398, N47399, N47400, N47401, N47402, N47403, N47404, N47405, N47406, N47407, N47408, N47409, N47410, N47411, N47412, N47413, N47414, N47415, N47416, N47417, N47418, N47420, N47421, N47422, N47423, N47424, N47425, N47426, N47427, N47428, N47429, N47430, N47432, N47433, N47434, N47435, N47436, N47437, N47438, N47439, N47440, N47441, N47442, N47443, N47444, N47445, N47446, N47447, N47448, N47449, N47450, N47452, N47453, N47455, N47456, N47457, N47458, N47459, N47460, N47461, N47462, N47463, N47464, N47465, N47466, N47467, N47468, N47469, N47470, N47472, N47473, N47474, N47476, N47477, N47478, N47479, N47480, N47481, N47482, N47483, N47484, N47485, N47486, N47487, N47488, N47489, N47490, N47491, N47492, N47493, N47494, N47496, N47497, N47498, N47500, N47501, N47502, N47503, N47504, N47505, N47506, N47507, N47508, N47510, N47511, N47512, N47513, N47515, N47517, N47518, N47519, N47520, N47521, N47522, N47523, N47524, N47525, N47526, N47527, N47528, N47529, N47530, N47531, N47532, N47533, N47534, N47536, N47537, N47538, N47539, N47540, N47541, N47542, N47543, N47544, N47545, N47547, N47548, N47549, N47550, N47551, N47552, N47553, N47554, N47555, N47556, N47557, N47558, N47559, N47560, N47561, N47562, N47563, N47564, N47565, N47566, N47567, N47568, N47569, N47570, N47571, N47572, N47573, N47574, N47575, N47576, N47577, N47578, N47579, N47580, N47581, N47582, N47583, N47584, N47585, N47586, N47587, N47588, N47589, N47590, N47591, N47592, N47593, N47594, N47595, N47596, N47597, N47598, N47599, N47600, N47601, N47602, N47603, N47604, N47605, N47606, N47607, N47608, N47609, N47610, N47612, N47613, N47614, N47615, N47616, N47617, N47618, N47619, N47620, N47622, N47623, N47624, N47625, N47626, N47627, N47628, N47630, N47631, N47632, N47633, N47634, N47636, N47639, N47641, N47642, N47643, N47644, N47646, N47647, N47648, N47649, N47650, N47651, N47652, N47653, N47654, N47655, N47656, N47657, N47658, N47659, N47660, N47662, N47664, N47665, N47666, N47667, N47668, N47670, N47671, N47672, N47674, N47675, N47676, N47677, N47678, N47679, N47680, N47681, N47682, N47683, N47684, N47685, N47686, N47687, N47688, N47689, N47690, N47691, N47692, N47693, N47694, N47695, N47696, N47697, N47698, N47699, N47700, N47701, N47702, N47703, N47704, N47705, N47706, N47707, N47708, N47709, N47710, N47711, N47712, N47713, N47714, N47716, N47718, N47719, N47720, N47721, N47722, N47723, N47724, N47725, N47726, N47728, N47729, N47730, N47731, N47732, N47733, N47734, N47735, N47736, N47737, N47738, N47739, N47741, N47742, N47743, N47744, N47745, N47746, N47747, N47748, N47749, N47750, N47751, N47753, N47754, N47755, N47756, N47757, N47759, N47760, N47761, N47762, N47763, N47764, N47765, N47766, N47767, N47768, N47769, N47770, N47772, N47773, N47774, N47775, N47776, N47777, N47778, N47779, N47780, N47781, N47782, N47783, N47784, N47785, N47786, N47787, N47788, N47789, N47790, N47791, N47792, N47793, N47794, N47795, N47796, N47797, N47798, N47799, N47800, N47801, N47802, N47803, N47804, N47805, N47806, N47807, N47808, N47810, N47811, N47812, N47813, N47814, N47815, N47816, N47817, N47818, N47819, N47820, N47821, N47822, N47823, N47824, N47825, N47826, N47827, N47828, N47829, N47830, N47831, N47832, N47833, N47834, N47835, N47836, N47837, N47839, N47840, N47841, N47842, N47843, N47845, N47846, N47847, N47848, N47849, N47850, N47851, N47852, N47853, N47854, N47855, N47856, N47857, N47858, N47859, N47860, N47861, N47862, N47863, N47864, N47865, N47866, N47867, N47868, N47869, N47870, N47871, N47872, N47874, N47875, N47876, N47877, N47878, N47880, N47881, N47882, N47883, N47884, N47885, N47886, N47887, N47888, N47889, N47890, N47891, N47892, N47893, N47894, N47895, N47896, N47897, N47898, N47899, N47900, N47901, N47903, N47904, N47905, N47906, N47907, N47908, N47909, N47910, N47911, N47912, N47913, N47914, N47915, N47916, N47917, N47918, N47919, N47920, N47922, N47923, N47925, N47926, N47927, N47928, N47929, N47930, N47931, N47932, N47933, N47934, N47935, N47936, N47937, N47938, N47939, N47940, N47941, N47942, N47943, N47944, N47945, N47946, N47948, N47949, N47950, N47951, N47952, N47953, N47954, N47955, N47957, N47958, N47959, N47960, N47961, N47962, N47963, N47964, N47965, N47966, N47967, N47968, N47969, N47970, N47971, N47972, N47973, N47974, N47975, N47976, N47977, N47978, N47979, N47980, N47981, N47982, N47983, N47984, N47985, N47986, N47987, N47988, N47989, N47990, N47991, N47992, N47993, N47994, N47995, N47996, N47997, N47998, N47999, N48000, N48001, N48002, N48003, N48004, N48005, N48006, N48007, N48008, N48009, N48010, N48011, N48012, N48013, N48014, N48015, N48016, N48017, N48018, N48019, N48020, N48021, N48022, N48023, N48024, N48025, N48026, N48027, N48029, N48030, N48031, N48032, N48033, N48034, N48035, N48036, N48037, N48038, N48040, N48041, N48042, N48043, N48044, N48045, N48046, N48047, N48049, N48050, N48051, N48052, N48053, N48054, N48055, N48056, N48058, N48059, N48061, N48062, N48063, N48064, N48065, N48066, N48067, N48068, N48069, N48070, N48071, N48072, N48073, N48074, N48075, N48076, N48077, N48078, N48079, N48080, N48081, N48082, N48083, N48084, N48085, N48087, N48088, N48089, N48090, N48091, N48092, N48093, N48094, N48095, N48096, N48097, N48098, N48099, N48100, N48102, N48103, N48104, N48105, N48106, N48107, N48108, N48109, N48110, N48111, N48113, N48115, N48116, N48117, N48118, N48119, N48120, N48121, N48122, N48123, N48124, N48125, N48126, N48127, N48129, N48130, N48131, N48132, N48133, N48135, N48137, N48138, N48139, N48140, N48141, N48142, N48143, N48145, N48147, N48148, N48149, N48150, N48152, N48153, N48154, N48155, N48156, N48157, N48158, N48159, N48160, N48161, N48162, N48164, N48165, N48167, N48168, N48169, N48170, N48171, N48172, N48173, N48174, N48175, N48176, N48177, N48178, N48179, N48180, N48181, N48182, N48183, N48184, N48185, N48187, N48188, N48189, N48190, N48191, N48192, N48193, N48194, N48195, N48196, N48197, N48198, N48199, N48200, N48201, N48202, N48203, N48204, N48205, N48206, N48207, N48208, N48210, N48211, N48212, N48213, N48214, N48216, N48217, N48219, N48220, N48221, N48222, N48223, N48224, N48225, N48226, N48227, N48228, N48229, N48230, N48231, N48233, N48234, N48235, N48236, N48237, N48238, N48240, N48241, N48242, N48243, N48244, N48245, N48246, N48248, N48249, N48250, N48251, N48252, N48253, N48254, N48255, N48256, N48257, N48258, N48259, N48260, N48262, N48263, N48264, N48265, N48267, N48268, N48269, N48270, N48271, N48272, N48273, N48274, N48275, N48277, N48278, N48279, N48280, N48281, N48282, N48283, N48284, N48286, N48287, N48288, N48289, N48290, N48291, N48292, N48293, N48294, N48295, N48296, N48297, N48298, N48299, N48300, N48302, N48303, N48306, N48307, N48308, N48309, N48311, N48312, N48313, N48314, N48315, N48316, N48317, N48318, N48319, N48320, N48321, N48323, N48325, N48326, N48327, N48328, N48329, N48331, N48332, N48333, N48334, N48335, N48336, N48337, N48338, N48339, N48340, N48341, N48342, N48343, N48344, N48345, N48346, N48347, N48349, N48350, N48351, N48352, N48353, N48354, N48356, N48357, N48358, N48359, N48360, N48362, N48363, N48364, N48365, N48366, N48367, N48368, N48369, N48370, N48371, N48372, N48374, N48375, N48377, N48379, N48380, N48382, N48383, N48384, N48385, N48386, N48387, N48388, N48389, N48390, N48391, N48392, N48393, N48394, N48395, N48396, N48397, N48398, N48399, N48400, N48401, N48404, N48405, N48406, N48407, N48408, N48409, N48410, N48411, N48412, N48413, N48414, N48415, N48416, N48417, N48418, N48419, N48420, N48421, N48422, N48423, N48424, N48425, N48426, N48427, N48428, N48429, N48430, N48431, N48432, N48433, N48435, N48436, N48437, N48438, N48439, N48440, N48441, N48442, N48443, N48444, N48445, N48446, N48447, N48448, N48449, N48450, N48451, N48452, N48454, N48455, N48456, N48457, N48459, N48461, N48462, N48463, N48464, N48465, N48466, N48468, N48469, N48470, N48471, N48472, N48473, N48474, N48475, N48476, N48477, N48478, N48479, N48480, N48481, N48482, N48483, N48484, N48485, N48486, N48488, N48489, N48490, N48491, N48492, N48493, N48494, N48495, N48496, N48497, N48498, N48499, N48500, N48501, N48502, N48503, N48504, N48505, N48506, N48507, N48508, N48511, N48512, N48513, N48515, N48516, N48517, N48518, N48519, N48521, N48523, N48524, N48525, N48526, N48527, N48528, N48529, N48530, N48531, N48532, N48533, N48534, N48535, N48536, N48537, N48538, N48539, N48540, N48541, N48542, N48543, N48545, N48546, N48547, N48549, N48550, N48551, N48552, N48553, N48555, N48557, N48558, N48559, N48560, N48561, N48562, N48563, N48564, N48565, N48566, N48567, N48568, N48569, N48570, N48571, N48572, N48573, N48574, N48575, N48576, N48578, N48579, N48581, N48582, N48583, N48584, N48585, N48586, N48587, N48588, N48589, N48590, N48591, N48592, N48593, N48594, N48595, N48596, N48597, N48598, N48600, N48601, N48602, N48603, N48604, N48605, N48606, N48607, N48609, N48610, N48611, N48612, N48613, N48614, N48615, N48616, N48617, N48618, N48619, N48620, N48621, N48622, N48623, N48624, N48625, N48626, N48627, N48628, N48629, N48630, N48631, N48632, N48633, N48634, N48635, N48636, N48637, N48638, N48639, N48641, N48642, N48643, N48644, N48645, N48646, N48647, N48649, N48650, N48651, N48652, N48653, N48654, N48655, N48656, N48657, N48658, N48659, N48660, N48661, N48662, N48663, N48664, N48665, N48666, N48667, N48668, N48669, N48670, N48671, N48672, N48673, N48674, N48675, N48676, N48677, N48679, N48680, N48681, N48682, N48683, N48684, N48685, N48686, N48687, N48688, N48689, N48690, N48691, N48692, N48693, N48694, N48695, N48696, N48697, N48698, N48699, N48700, N48701, N48702, N48704, N48705, N48706, N48707, N48708, N48709, N48710, N48711, N48712, N48713, N48714, N48715, N48716, N48718, N48720, N48721, N48722, N48723, N48724, N48725, N48726, N48727, N48728, N48729, N48730, N48731, N48732, N48734, N48735, N48736, N48737, N48738, N48739, N48740, N48741, N48742, N48744, N48745, N48746, N48747, N48748, N48749, N48750, N48751, N48752, N48753, N48754, N48755, N48756, N48757, N48758, N48759, N48760, N48762, N48763, N48764, N48765, N48766, N48767, N48768, N48769, N48770, N48771, N48772, N48773, N48774, N48775, N48776, N48777, N48778, N48779, N48780, N48781, N48782, N48783, N48784, N48785, N48786, N48787, N48788, N48789, N48790, N48791, N48792, N48793, N48794, N48795, N48796, N48797, N48798, N48799, N48800, N48801, N48802, N48803, N48804, N48805, N48806, N48807, N48808, N48809, N48810, N48811, N48812, N48813, N48814, N48815, N48817, N48818, N48819, N48820, N48821, N48822, N48823, N48824, N48825, N48826, N48828, N48829, N48830, N48832, N48833, N48835, N48836, N48837, N48838, N48839, N48840, N48841, N48842, N48843, N48844, N48845, N48846, N48847, N48848, N48849, N48850, N48851, N48852, N48853, N48854, N48855, N48856, N48857, N48858, N48859, N48860, N48861, N48862, N48863, N48864, N48865, N48866, N48867, N48868, N48869, N48870, N48871, N48872, N48873, N48874, N48875, N48876, N48877, N48878, N48879, N48880, N48881, N48882, N48883, N48884, N48885, N48886, N48887, N48888, N48889, N48890, N48892, N48894, N48895, N48897, N48898, N48899, N48900, N48901, N48902, N48903, N48904, N48905, N48906, N48907, N48909, N48910, N48911, N48912, N48913, N48914, N48915, N48916, N48917, N48918, N48919, N48920, N48921, N48922, N48923, N48924, N48925, N48926, N48927, N48928, N48929, N48930, N48932, N48933, N48934, N48935, N48936, N48937, N48938, N48939, N48940, N48941, N48943, N48944, N48945, N48946, N48947, N48948, N48949, N48950, N48951, N48952, N48954, N48955, N48956, N48957, N48958, N48959, N48960, N48961, N48962, N48963, N48964, N48965, N48966, N48967, N48969, N48971, N48972, N48973, N48974, N48975, N48977, N48978, N48979, N48980, N48981, N48982, N48983, N48984, N48985, N48986, N48988, N48989, N48990, N48991, N48992, N48994, N48995, N48996, N48997, N48998, N48999, N49000, N49001, N49002, N49003, N49004, N49005, N49006, N49007, N49008, N49009, N49011, N49012, N49013, N49014, N49015, N49016, N49017, N49018, N49019, N49020, N49021, N49022, N49023, N49024, N49025, N49026, N49028, N49030, N49033, N49034, N49035, N49036, N49037, N49038, N49039, N49040, N49041, N49042, N49043, N49044, N49045, N49046, N49048, N49049, N49050, N49051, N49052, N49053, N49054, N49055, N49056, N49057, N49058, N49059, N49060, N49061, N49062, N49063, N49064, N49065, N49066, N49068, N49069, N49070, N49071, N49072, N49073, N49074, N49075, N49076, N49077, N49078, N49079, N49080, N49081, N49082, N49083, N49084, N49085, N49086, N49087, N49088, N49090, N49091, N49092, N49093, N49094, N49095, N49097, N49098, N49099, N49100, N49101, N49102, N49103, N49104, N49105, N49107, N49108, N49109, N49110, N49111, N49112, N49113, N49114, N49115, N49118, N49119, N49120, N49121, N49123, N49124, N49125, N49126, N49127, N49128, N49130, N49131, N49132, N49133, N49135, N49136, N49137, N49138, N49139, N49140, N49141, N49142, N49143, N49144, N49145, N49146, N49147, N49148, N49149, N49150, N49151, N49153, N49154, N49155, N49156, N49157, N49158, N49159, N49160, N49161, N49162, N49163, N49164, N49165, N49166, N49167, N49168, N49169, N49170, N49171, N49172, N49173, N49174, N49175, N49176, N49177, N49178, N49180, N49181, N49182, N49183, N49185, N49186, N49187, N49188, N49189, N49190, N49191, N49192, N49193, N49195, N49196, N49197, N49198, N49199, N49200, N49201, N49202, N49204, N49205, N49206, N49207, N49208, N49209, N49210, N49211, N49212, N49213, N49214, N49215, N49216, N49217, N49218, N49220, N49222, N49223, N49224, N49225, N49226, N49227, N49228, N49229, N49230, N49231, N49232, N49233, N49234, N49235, N49236, N49237, N49239, N49240, N49241, N49242, N49243, N49244, N49245, N49246, N49247, N49248, N49249, N49250, N49251, N49252, N49253, N49254, N49255, N49256, N49257, N49258, N49259, N49260, N49261, N49262, N49263, N49265, N49266, N49267, N49268, N49269, N49270, N49271, N49272, N49274, N49275, N49276, N49277, N49279, N49280, N49281, N49282, N49284, N49285, N49286, N49287, N49288, N49289, N49290, N49291, N49292, N49293, N49294, N49295, N49296, N49297, N49298, N49300, N49301, N49302, N49303, N49304, N49305, N49306, N49308, N49309, N49310, N49311, N49312, N49313, N49314, N49315, N49317, N49318, N49319, N49320, N49321, N49322, N49323, N49324, N49325, N49326, N49327, N49328, N49330, N49331, N49333, N49334, N49335, N49336, N49338, N49339, N49340, N49341, N49342, N49343, N49344, N49345, N49346, N49347, N49348, N49349, N49350, N49351, N49352, N49353, N49354, N49355, N49356, N49357, N49358, N49359, N49360, N49363, N49364, N49366, N49367, N49368, N49369, N49370, N49371, N49372, N49373, N49374, N49375, N49377, N49378, N49380, N49381, N49382, N49383, N49384, N49385, N49386, N49387, N49388, N49389, N49390, N49391, N49392, N49393, N49394, N49395, N49396, N49397, N49398, N49399, N49400, N49401, N49402, N49403, N49404, N49405, N49406, N49407, N49408, N49409, N49410, N49411, N49412, N49413, N49414, N49415, N49416, N49417, N49418, N49419, N49420, N49422, N49423, N49424, N49425, N49426, N49428, N49429, N49430, N49431, N49432, N49433, N49434, N49435, N49436, N49437, N49438, N49439, N49441, N49442, N49443, N49444, N49445, N49446, N49447, N49448, N49449, N49450, N49451, N49452, N49453, N49454, N49456, N49457, N49459, N49460, N49461, N49462, N49463, N49464, N49465, N49467, N49468, N49469, N49470, N49471, N49473, N49474, N49475, N49476, N49477, N49478, N49479, N49480, N49481, N49483, N49484, N49485, N49486, N49487, N49488, N49489, N49490, N49491, N49492, N49493, N49494, N49495, N49496, N49497, N49498, N49499, N49500, N49501, N49502, N49503, N49504, N49506, N49507, N49508, N49509, N49510, N49511, N49512, N49513, N49514, N49515, N49516, N49517, N49518, N49519, N49520, N49521, N49522, N49523, N49524, N49525, N49526, N49527, N49528, N49529, N49530, N49531, N49532, N49533, N49534, N49535, N49536, N49537, N49538, N49539, N49540, N49541, N49542, N49543, N49544, N49545, N49546, N49547, N49548, N49549, N49550, N49551, N49552, N49555, N49556, N49557, N49558, N49559, N49560, N49562, N49563, N49564, N49565, N49566, N49567, N49568, N49569, N49570, N49571, N49572, N49573, N49574, N49575, N49576, N49577, N49578, N49579, N49580, N49581, N49582, N49583, N49584, N49585, N49586, N49587, N49589, N49590, N49591, N49592, N49593, N49594, N49595, N49596, N49597, N49598, N49599, N49600, N49601, N49602, N49603, N49604, N49605, N49606, N49607, N49608, N49609, N49610, N49611, N49612, N49613, N49614, N49616, N49617, N49618, N49619, N49620, N49622, N49624, N49625, N49626, N49628, N49629, N49630, N49631, N49632, N49633, N49634, N49635, N49636, N49637, N49638, N49639, N49640, N49641, N49643, N49644, N49645, N49646, N49647, N49648, N49649, N49650, N49651, N49652, N49653, N49655, N49656, N49657, N49658, N49660, N49661, N49662, N49663, N49664, N49665, N49666, N49667, N49668, N49669, N49670, N49672, N49673, N49674, N49675, N49676, N49677, N49678, N49679, N49680, N49681, N49682, N49683, N49684, N49685, N49687, N49688, N49689, N49690, N49691, N49692, N49693, N49694, N49695, N49696, N49697, N49698, N49699, N49700, N49701, N49702, N49703, N49705, N49706, N49707, N49708, N49709, N49710, N49711, N49712, N49713, N49714, N49715, N49716, N49717, N49718, N49719, N49720, N49721, N49722, N49723, N49724, N49725, N49726, N49727, N49728, N49729, N49730, N49731, N49732, N49733, N49734, N49735, N49736, N49737, N49739, N49740, N49741, N49742, N49743, N49744, N49745, N49746, N49747, N49748, N49749, N49750, N49751, N49752, N49753, N49754, N49755, N49756, N49757, N49758, N49759, N49760, N49761, N49763, N49765, N49767, N49768, N49769, N49770, N49771, N49772, N49773, N49774, N49776, N49777, N49778, N49779, N49780, N49781, N49782, N49783, N49784, N49785, N49787, N49788, N49789, N49790, N49791, N49792, N49794, N49795, N49796, N49797, N49798, N49799, N49800, N49801, N49802, N49803, N49804, N49805, N49806, N49807, N49808, N49809, N49810, N49811, N49812, N49813, N49814, N49815, N49816, N49817, N49818, N49819, N49820, N49821, N49822, N49823, N49824, N49825, N49826, N49827, N49828, N49829, N49830, N49831, N49832, N49835, N49836, N49837, N49838, N49839, N49840, N49841, N49842, N49843, N49844, N49845, N49846, N49847, N49848, N49849, N49850, N49851, N49852, N49853, N49854, N49855, N49856, N49857, N49858, N49860, N49861, N49862, N49863, N49864, N49865, N49866, N49867, N49868, N49869, N49870, N49871, N49872, N49873, N49874, N49875, N49876, N49877, N49878, N49879, N49880, N49881, N49882, N49883, N49884, N49885, N49886, N49887, N49888, N49889, N49890, N49891, N49892, N49894, N49895, N49896, N49898, N49899, N49901, N49903, N49904, N49905, N49906, N49907, N49908, N49909, N49910, N49911, N49912, N49913, N49914, N49915, N49917, N49918, N49919, N49920, N49921, N49923, N49924, N49925, N49926, N49927, N49928, N49929, N49930, N49931, N49932, N49933, N49934, N49935, N49936, N49937, N49938, N49939, N49940, N49941, N49942, N49943, N49944, N49945, N49946, N49947, N49948, N49949, N49950, N49951, N49952, N49953, N49954, N49955, N49956, N49957, N49958, N49959, N49960, N49961, N49962, N49963, N49964, N49965, N49966, N49967, N49969, N49970, N49972, N49973, N49974, N49975, N49976, N49977, N49979, N49980, N49981, N49982, N49983, N49985, N49986, N49987, N49988, N49989, N49991, N49992, N49993, N49994, N49995, N49996, N49997, N49998, N49999, N50000, N50001, N50003, N50004, N50005, N50006, N50007, N50008, N50009, N50010, N50011, N50012, N50013, N50014, N50015, N50016, N50017, N50018, N50019, N50020, N50021, N50022, N50023, N50024, N50025, N50026, N50027, N50028, N50030, N50031, N50032, N50033, N50034, N50035, N50036, N50037, N50038, N50039, N50040, N50041, N50042, N50043, N50044, N50045, N50046, N50047, N50048, N50049, N50050, N50051, N50053, N50054, N50055, N50056, N50057, N50058, N50059, N50060, N50061, N50062, N50063, N50064, N50065, N50066, N50067, N50068, N50069, N50070, N50071, N50072, N50073, N50074, N50075, N50076, N50077, N50078, N50079, N50080, N50081, N50082, N50084, N50085, N50086, N50087, N50089, N50090, N50091, N50092, N50093, N50094, N50095, N50096, N50098, N50099, N50100, N50101, N50102, N50103, N50104, N50105, N50106, N50108, N50109, N50110, N50111, N50113, N50115, N50116, N50117, N50119, N50120, N50121, N50122, N50123, N50124, N50125, N50126, N50129, N50130, N50131, N50132, N50133, N50134, N50135, N50136, N50137, N50138, N50139, N50140, N50142, N50143, N50144, N50145, N50146, N50147, N50148, N50149, N50150, N50151, N50152, N50153, N50154, N50157, N50158, N50159, N50160, N50161, N50162, N50163, N50164, N50165, N50166, N50167, N50168, N50169, N50170, N50171, N50172, N50173, N50174, N50175, N50177, N50179, N50180, N50181, N50182, N50183, N50185, N50186, N50187, N50188, N50189, N50190, N50191, N50192, N50193, N50194, N50195, N50196, N50197, N50200, N50201, N50203, N50204, N50205, N50206, N50208, N50209, N50210, N50211, N50212, N50213, N50214, N50215, N50216, N50217, N50218, N50220, N50221, N50222, N50223, N50224, N50225, N50226, N50227, N50229, N50230, N50231, N50232, N50234, N50235, N50236, N50237, N50238, N50239, N50240, N50241, N50242, N50243, N50244, N50246, N50247, N50248, N50249, N50250, N50251, N50252, N50253, N50254, N50255, N50256, N50258, N50259, N50260, N50262, N50263, N50264, N50265, N50266, N50267, N50268, N50270, N50272, N50273, N50274, N50276, N50277, N50278, N50279, N50280, N50281, N50282, N50283, N50284, N50285, N50286, N50287, N50288, N50289, N50290, N50291, N50292, N50293, N50294, N50295, N50296, N50297, N50298, N50299, N50300, N50301, N50302, N50303, N50304, N50305, N50306, N50307, N50308, N50309, N50310, N50312, N50313, N50315, N50316, N50317, N50318, N50319, N50320, N50321, N50323, N50324, N50325, N50326, N50327, N50328, N50329, N50330, N50331, N50332, N50333, N50334, N50335, N50336, N50337, N50338, N50339, N50340, N50341, N50342, N50343, N50344, N50345, N50346, N50347, N50349, N50350, N50351, N50352, N50353, N50354, N50355, N50356, N50357, N50358, N50359, N50360, N50361, N50362, N50363, N50364, N50366, N50367, N50368, N50369, N50370, N50371, N50372, N50373, N50374, N50375, N50376, N50377, N50378, N50379, N50380, N50381, N50382, N50383, N50384, N50385, N50386, N50387, N50388, N50389, N50390, N50391, N50392, N50393, N50396, N50397, N50398, N50399, N50400, N50401, N50402, N50403, N50404, N50405, N50406, N50407, N50408, N50409, N50410, N50411, N50412, N50413, N50414, N50415, N50416, N50417, N50418, N50419, N50420, N50421, N50422, N50424, N50425, N50426, N50427, N50428, N50429, N50430, N50432, N50433, N50434, N50435, N50436, N50437, N50438, N50439, N50440, N50441, N50442, N50443, N50444, N50445, N50446, N50447, N50448, N50449, N50450, N50451, N50452, N50453, N50454, N50456, N50457, N50458, N50459, N50461, N50462, N50463, N50464, N50465, N50466, N50467, N50468, N50469, N50470, N50471, N50472, N50473, N50474, N50475, N50476, N50477, N50478, N50479, N50480, N50481, N50482, N50483, N50484, N50485, N50486, N50487, N50488, N50489, N50490, N50491, N50492, N50493, N50494, N50495, N50496, N50497, N50498, N50499, N50500, N50501, N50502, N50503, N50504, N50506, N50507, N50508, N50509, N50510, N50512, N50513, N50514, N50515, N50516, N50517, N50518, N50519, N50520, N50521, N50522, N50523, N50524, N50525, N50526, N50527, N50528, N50529, N50530, N50531, N50532, N50533, N50535, N50536, N50537, N50538, N50539, N50540, N50541, N50542, N50543, N50544, N50545, N50546, N50547, N50548, N50549, N50550, N50551, N50552, N50553, N50554, N50555, N50556, N50557, N50558, N50559, N50560, N50561, N50562, N50563, N50564, N50565, N50566, N50567, N50569, N50570, N50571, N50572, N50573, N50574, N50575, N50576, N50577, N50578, N50579, N50580, N50581, N50582, N50583, N50584, N50585, N50586, N50588, N50589, N50590, N50592, N50593, N50596, N50598, N50599, N50600, N50601, N50603, N50604, N50605, N50606, N50607, N50608, N50609, N50610, N50611, N50612, N50613, N50614, N50615, N50616, N50617, N50618, N50619, N50620, N50621, N50622, N50623, N50624, N50625, N50627, N50628, N50629, N50630, N50631, N50632, N50633, N50635, N50636, N50637, N50638, N50639, N50640, N50641, N50642, N50643, N50644, N50645, N50646, N50648, N50649, N50650, N50651, N50652, N50653, N50654, N50655, N50656, N50657, N50658, N50659, N50660, N50661, N50662, N50663, N50664, N50665, N50667, N50668, N50669, N50670, N50671, N50672, N50673, N50674, N50675, N50676, N50677, N50678, N50679, N50680, N50681, N50682, N50683, N50684, N50685, N50687, N50688, N50689, N50690, N50691, N50693, N50694, N50695, N50696, N50697, N50698, N50699, N50700, N50701, N50702, N50703, N50705, N50706, N50707, N50708, N50709, N50710, N50711, N50712, N50713, N50714, N50715, N50716, N50717, N50718, N50719, N50720, N50721, N50722, N50723, N50724, N50725, N50726, N50728, N50729, N50730, N50731, N50732, N50733, N50734, N50735, N50736, N50737, N50738, N50739, N50741, N50742, N50743, N50744, N50745, N50746, N50747, N50748, N50749, N50750, N50751, N50752, N50753, N50754, N50755, N50756, N50757, N50758, N50759, N50760, N50761, N50762, N50763, N50764, N50765, N50766, N50767, N50768, N50769, N50770, N50771, N50772, N50773, N50774, N50775, N50776, N50777, N50778, N50779, N50780, N50781, N50782, N50783, N50784, N50785, N50786, N50787, N50788, N50789, N50790, N50791, N50792, N50793, N50794, N50795, N50796, N50797, N50798, N50799, N50800, N50801, N50802, N50803, N50804, N50805, N50806, N50807, N50808, N50809, N50810, N50811, N50812, N50813, N50814, N50815, N50816, N50817, N50818, N50819, N50820, N50821, N50822, N50824, N50825, N50826, N50827, N50828, N50829, N50830, N50831, N50832, N50833, N50834, N50835, N50836, N50837, N50838, N50839, N50840, N50841, N50842, N50843, N50844, N50845, N50846, N50847, N50848, N50849, N50850, N50851, N50852, N50853, N50855, N50856, N50857, N50858, N50859, N50860, N50862, N50864, N50865, N50866, N50867, N50868, N50869, N50870, N50871, N50872, N50873, N50874, N50875, N50876, N50878, N50879, N50880, N50881, N50882, N50883, N50884, N50885, N50886, N50887, N50888, N50891, N50892, N50893, N50894, N50895, N50896, N50898, N50899, N50900, N50901, N50902, N50903, N50904, N50905, N50906, N50908, N50910, N50911, N50912, N50913, N50914, N50915, N50916, N50918, N50919, N50920, N50921, N50922, N50923, N50924, N50925, N50926, N50927, N50928, N50929, N50930, N50932, N50933, N50934, N50936, N50937, N50939, N50941, N50942, N50944, N50945, N50946, N50949, N50950, N50952, N50953, N50954, N50955, N50956, N50957, N50958, N50959, N50960, N50961, N50962, N50963, N50964, N50965, N50966, N50968, N50969, N50970, N50971, N50972, N50973, N50975, N50976, N50978, N50979, N50980, N50981, N50982, N50983, N50984, N50985, N50986, N50988, N50989, N50990, N50991, N50992, N50993, N50994, N50995, N50996, N50997, N50998, N50999, N51000, N51001, N51002, N51003, N51004, N51005, N51006, N51007, N51008, N51009, N51010, N51011, N51012, N51013, N51014, N51015, N51016, N51017, N51018, N51019, N51020, N51021, N51022, N51023, N51026, N51027, N51028, N51029, N51030, N51031, N51032, N51033, N51034, N51036, N51037, N51039, N51040, N51041, N51043, N51044, N51045, N51047, N51048, N51049, N51050, N51052, N51053, N51054, N51055, N51056, N51057, N51058, N51059, N51060, N51061, N51062, N51064, N51065, N51066, N51067, N51068, N51069, N51070, N51071, N51072, N51073, N51074, N51075, N51076, N51077, N51078, N51079, N51080, N51081, N51082, N51083, N51084, N51085, N51086, N51087, N51089, N51090, N51091, N51093, N51094, N51095, N51096, N51097, N51098, N51101, N51102, N51103, N51105, N51106, N51107, N51108, N51110, N51111, N51112, N51113, N51114, N51115, N51116, N51117, N51118, N51119, N51120, N51121, N51122, N51123, N51124, N51125, N51126, N51127, N51128, N51129, N51130, N51131, N51132, N51133, N51134, N51135, N51136, N51137, N51139, N51140, N51141, N51142, N51143, N51144, N51145, N51146, N51147, N51148, N51150, N51151, N51152, N51153, N51154, N51155, N51156, N51157, N51159, N51160, N51161, N51162, N51163, N51164, N51165, N51166, N51167, N51168, N51169, N51170, N51171, N51172, N51173, N51174, N51175, N51176, N51177, N51178, N51179, N51180, N51181, N51182, N51183, N51184, N51185, N51186, N51187, N51188, N51189, N51190, N51191, N51193, N51194, N51195, N51197, N51198, N51200, N51201, N51202, N51203, N51204, N51205, N51206, N51207, N51208, N51209, N51210, N51211, N51212, N51213, N51214, N51215, N51216, N51217, N51219, N51220, N51221, N51222, N51223, N51224, N51225, N51226, N51228, N51229, N51230, N51231, N51232, N51233, N51234, N51235, N51236, N51237, N51238, N51239, N51240, N51242, N51244, N51245, N51246, N51248, N51249, N51250, N51251, N51252, N51253, N51254, N51255, N51256, N51257, N51258, N51259, N51260, N51261, N51262, N51263, N51265, N51266, N51267, N51268, N51269, N51270, N51271, N51272, N51273, N51274, N51276, N51277, N51278, N51279, N51280, N51281, N51282, N51283, N51284, N51285, N51286, N51287, N51288, N51289, N51290, N51291, N51292, N51294, N51295, N51296, N51297, N51298, N51299, N51300, N51301, N51302, N51303, N51304, N51305, N51306, N51308, N51309, N51310, N51311, N51312, N51313, N51314, N51315, N51316, N51317, N51318, N51319, N51320, N51321, N51322, N51324, N51325, N51326, N51327, N51328, N51329, N51331, N51332, N51333, N51334, N51335, N51336, N51338, N51340, N51341, N51342, N51343, N51344, N51345, N51346, N51347, N51348, N51349, N51350, N51351, N51352, N51353, N51355, N51357, N51358, N51359, N51360, N51361, N51362, N51363, N51364, N51365, N51366, N51367, N51368, N51369, N51371, N51372, N51374, N51375, N51376, N51377, N51378, N51379, N51381, N51382, N51383, N51384, N51385, N51386, N51387, N51388, N51389, N51390, N51392, N51394, N51395, N51396, N51397, N51398, N51399, N51400, N51401, N51402, N51403, N51405, N51406, N51407, N51408, N51409, N51410, N51411, N51412, N51413, N51414, N51415, N51416, N51417, N51418, N51419, N51420, N51421, N51422, N51423, N51424, N51425, N51426, N51427, N51428, N51430, N51431, N51432, N51433, N51434, N51435, N51436, N51437, N51438, N51439, N51440, N51441, N51442, N51443, N51444, N51445, N51446, N51447, N51448, N51449, N51450, N51452, N51453, N51454, N51455, N51456, N51457, N51458, N51459, N51460, N51461, N51463, N51464, N51465, N51466, N51467, N51468, N51469, N51470, N51471, N51473, N51474, N51475, N51476, N51477, N51478, N51479, N51480, N51481, N51482, N51483, N51484, N51485, N51486, N51487, N51488, N51489, N51490, N51491, N51492, N51493, N51494, N51495, N51496, N51497, N51499, N51500, N51502, N51504, N51505, N51506, N51507, N51508, N51509, N51510, N51511, N51512, N51513, N51514, N51515, N51517, N51518, N51519, N51520, N51522, N51523, N51524, N51525, N51526, N51527, N51528, N51529, N51530, N51531, N51533, N51534, N51537, N51538, N51539, N51541, N51542, N51543, N51544, N51545, N51546, N51547, N51548, N51550, N51551, N51552, N51553, N51554, N51555, N51556, N51557, N51558, N51559, N51560, N51561, N51562, N51563, N51564, N51565, N51566, N51567, N51568, N51569, N51570, N51572, N51573, N51574, N51575, N51576, N51577, N51578, N51579, N51580, N51581, N51582, N51583, N51584, N51586, N51587, N51588, N51589, N51590, N51591, N51592, N51593, N51594, N51595, N51596, N51597, N51598, N51599, N51600, N51601, N51602, N51603, N51604, N51605, N51606, N51607, N51608, N51609, N51610, N51612, N51613, N51614, N51615, N51616, N51617, N51618, N51619, N51620, N51621, N51622, N51623, N51624, N51625, N51626, N51627, N51628, N51629, N51630, N51631, N51632, N51633, N51634, N51635, N51636, N51637, N51638, N51639, N51640, N51641, N51642, N51643, N51644, N51645, N51646, N51647, N51648, N51649, N51650, N51651, N51652, N51653, N51654, N51655, N51656, N51657, N51658, N51659, N51660, N51661, N51662, N51663, N51664, N51665, N51666, N51667, N51668, N51669, N51670, N51671, N51672, N51673, N51674, N51675, N51676, N51677, N51678, N51679, N51680, N51681, N51682, N51683, N51684, N51685, N51686, N51687, N51688, N51689, N51690, N51691, N51692, N51693, N51694, N51695, N51696, N51697, N51698, N51699, N51700, N51701, N51702, N51703, N51704, N51705, N51706, N51707, N51708, N51709, N51710, N51711, N51712, N51713, N51714, N51715, N51716, N51717, N51718, N51719, N51720, N51721, N51722, N51723, N51724, N51725, N51726, N51727, N51728, N51729, N51730, N51731, N51732, N51733, N51735, N51736, N51737, N51738, N51739, N51740, N51741, N51742, N51743, N51745, N51746, N51747, N51748, N51749, N51750, N51751, N51752, N51754, N51755, N51756, N51757, N51758, N51759, N51760, N51761, N51762, N51763, N51764, N51765, N51766, N51767, N51768, N51769, N51770, N51771, N51772, N51773, N51774, N51775, N51776, N51777, N51778, N51779, N51780, N51781, N51782, N51783, N51784, N51785, N51786, N51787, N51788, N51789, N51790, N51791, N51792, N51793, N51794, N51795, N51796, N51797, N51798, N51799, N51800, N51801, N51802, N51803, N51804, N51805, N51806, N51807, N51808, N51809, N51810, N51811, N51812, N51813, N51814, N51815, N51816, N51817, N51818, N51819, N51820, N51821, N51822, N51823, N51824, N51825, N51826, N51827, N51828, N51829, N51830, N51831, N51832, N51833, N51834, N51835, N51836, N51837, N51838, N51839, N51840, N51841, N51842, N51844, N51845, N51846, N51847, N51848, N51849, N51850, N51851, N51852, N51853, N51854, N51855, N51856, N51857, N51858, N51859, N51860, N51861, N51862, N51863, N51864, N51865, N51867, N51868, N51869, N51870, N51871, N51872, N51873, N51874, N51875, N51876, N51877, N51878, N51879, N51880, N51881, N51882, N51883, N51884, N51885, N51886, N51887, N51888, N51889, N51890, N51891, N51892, N51893, N51894, N51896, N51897, N51898, N51899, N51900, N51901, N51902, N51903, N51904, N51905, N51906, N51907, N51908, N51909, N51910, N51911, N51912, N51913, N51914, N51915, N51916, N51917, N51918, N51919, N51920, N51921, N51922, N51923, N51924, N51926, N51927, N51928, N51929, N51930, N51931, N51932, N51933, N51934, N51935, N51937, N51938, N51939, N51940, N51941, N51942, N51943, N51944, N51945, N51946, N51947, N51948, N51949, N51950, N51951, N51952, N51953, N51954, N51955, N51956, N51957, N51958, N51959, N51960, N51961, N51962, N51963, N51964, N51965, N51966, N51967, N51968, N51969, N51970, N51971, N51973, N51974, N51975, N51976, N51977, N51978, N51979, N51980, N51981, N51982, N51983, N51984, N51985, N51986, N51987, N51988, N51989, N51990, N51991, N51992, N51993, N51994, N51995, N51996, N51997, N51998, N51999, N52000, N52001, N52002, N52003, N52004, N52005, N52006, N52007, N52008, N52009, N52011, N52012, N52013, N52014, N52015, N52016, N52017, N52018, N52019, N52020, N52021, N52022, N52023, N52025, N52026, N52027, N52028, N52029, N52030, N52031, N52032, N52033, N52034, N52035, N52036, N52037, N52038, N52039, N52040, N52041, N52042, N52043, N52044, N52045, N52046, N52047, N52048, N52049, N52050, N52051, N52052, N52053, N52054, N52055, N52056, N52057, N52058, N52059, N52060, N52061, N52062, N52063, N52064, N52065, N52066, N52067, N52069, N52070, N52071, N52072, N52073, N52074, N52075, N52076, N52077, N52078, N52079, N52080, N52081, N52082, N52083, N52085, N52086, N52087, N52089, N52090, N52091, N52092, N52094, N52095, N52096, N52097, N52098, N52099, N52100, N52101, N52102, N52103, N52105, N52106, N52107, N52108, N52109, N52110, N52111, N52112, N52113, N52114, N52115, N52116, N52117, N52118, N52119, N52120, N52121, N52122, N52123, N52124, N52125, N52126, N52127, N52128, N52129, N52130, N52131, N52132, N52133, N52134, N52135, N52136, N52137, N52138, N52139, N52140, N52141, N52142, N52143, N52144, N52145, N52146, N52147, N52148, N52149, N52150, N52151, N52152, N52153, N52154, N52155, N52156, N52157, N52158, N52159, N52160, N52161, N52162, N52163, N52164, N52165, N52166, N52167, N52168, N52169, N52170, N52171, N52172, N52173, N52174, N52175, N52176, N52177, N52178, N52179, N52180, N52182, N52183, N52184, N52185, N52186, N52187, N52188, N52189, N52190, N52191, N52192, N52193, N52194, N52195, N52196, N52197, N52198, N52199, N52200, N52201, N52202, N52203, N52204, N52205, N52207, N52208, N52209, N52210, N52211, N52212, N52213, N52214, N52215, N52216, N52217, N52218, N52219, N52220, N52221, N52222, N52223, N52224, N52225, N52226, N52227, N52228, N52229, N52230, N52231, N52232, N52233, N52234, N52235, N52236, N52237, N52239, N52240, N52241, N52242, N52243, N52244, N52245, N52246, N52247, N52248, N52249, N52250, N52251, N52252, N52253, N52254, N52255, N52256, N52257, N52258, N52259, N52260, N52261, N52262, N52263, N52264, N52265, N52266, N52267, N52268, N52269, N52270, N52271, N52272, N52273, N52274, N52275, N52276, N52277, N52278, N52279, N52280, N52281, N52282, N52283, N52284, N52285, N52286, N52287, N52288, N52289, N52290, N52291, N52292, N52293, N52294, N52295, N52296, N52297, N52298, N52299, N52300, N52301, N52302, N52303, N52304, N52305, N52306, N52307, N52308, N52309, N52310, N52311, N52312, N52313, N52314, N52315, N52316, N52317, N52318, N52319, N52320, N52321, N52322, N52323, N52324, N52325, N52327, N52329, N52330, N52331, N52332, N52333, N52334, N52335, N52336, N52337, N52338, N52339, N52340, N52341, N52342, N52343, N52344, N52345, N52346, N52347, N52348, N52349, N52350, N52351, N52352, N52353, N52354, N52355, N52356, N52357, N52358, N52359, N52360, N52361, N52362, N52363, N52364, N52365, N52366, N52367, N52368, N52369, N52370, N52371, N52372, N52373, N52374, N52375, N52376, N52377, N52378, N52379, N52380, N52381, N52382, N52383, N52384, N52385, N52386, N52387, N52388, N52389, N52390, N52391, N52392, N52393, N52394, N52395, N52396, N52397, N52398, N52399, N52400, N52401, N52402, N52403, N52404, N52405, N52406, N52407, N52408, N52409, N52410, N52411, N52412, N52413, N52414, N52415, N52416, N52417, N52418, N52419, N52420, N52421, N52422, N52423, N52424, N52425, N52426, N52427, N52428, N52429, N52431, N52432, N52433, N52434, N52435, N52436, N52437, N52438, N52439, N52440, N52441, N52442, N52443, N52444, N52445, N52446, N52447, N52448, N52449, N52450, N52451, N52452, N52453, N52455, N52456, N52457, N52458, N52459, N52460, N52461, N52462, N52463, N52464, N52465, N52466, N52467, N52468, N52469, N52470, N52471, N52472, N52473, N52474, N52475, N52476, N52477, N52478, N52479, N52480, N52481, N52482, N52483, N52484, N52485, N52486, N52487, N52488, N52489, N52490, N52491, N52492, N52493, N52494, N52495, N52496, N52497, N52498, N52499, N52500, N52501, N52502, N52503, N52504, N52505, N52506, N52507, N52508, N52509, N52510, N52511, N52512, N52513, N52514, N52515, N52516, N52517, N52519, N52520, N52521, N52522, N52523, N52524, N52525, N52526, N52527, N52528, N52529, N52530, N52531, N52532, N52533, N52534, N52535, N52536, N52537, N52538, N52539, N52540, N52541, N52542, N52543, N52544, N52546, N52547, N52548, N52549, N52550, N52551, N52552, N52553, N52554, N52555, N52556, N52557, N52558, N52559, N52560, N52561, N52562, N52563, N52564, N52565, N52566, N52567, N52568, N52569, N52570, N52571, N52572, N52573, N52574, N52575, N52576, N52578, N52579, N52580, N52581, N52582, N52583, N52584, N52585, N52586, N52587, N52588, N52589, N52590, N52591, N52592, N52593, N52594, N52595, N52596, N52597, N52598, N52599, N52600, N52601, N52602, N52603, N52604, N52606, N52608, N52609, N52610, N52611, N52613, N52614, N52615, N52616, N52617, N52618, N52619, N52620, N52621, N52622, N52623, N52624, N52625, N52626, N52627, N52628, N52629, N52630, N52631, N52632, N52633, N52634, N52636, N52637, N52638, N52639, N52640, N52641, N52642, N52643, N52644, N52645, N52646, N52647, N52648, N52649, N52650, N52651, N52652, N52653, N52654, N52655, N52656, N52657, N52658, N52659, N52661, N52662, N52663, N52664, N52665, N52666, N52667, N52668, N52669, N52670, N52671, N52672, N52673, N52674, N52675, N52676, N52677, N52678, N52679, N52680, N52681, N52682, N52683, N52684, N52685, N52686, N52687, N52688, N52689, N52690, N52691, N52692, N52693, N52694, N52695, N52696, N52697, N52698, N52699, N52700, N52701, N52702, N52703, N52704, N52705, N52706, N52707, N52708, N52709, N52710, N52711, N52712, N52713, N52714, N52715, N52716, N52717, N52718, N52719, N52720, N52721, N52722, N52723, N52724, N52725, N52726, N52727, N52728, N52729, N52730, N52731, N52732, N52733, N52734, N52735, N52736, N52737, N52738, N52739, N52740, N52741, N52742, N52743, N52744, N52745, N52746, N52747, N52748, N52749, N52750, N52751, N52752, N52753, N52754, N52755, N52756, N52757, N52758, N52759, N52760, N52761, N52762, N52763, N52764, N52765, N52766, N52767, N52768, N52769, N52770, N52771, N52772, N52773, N52774, N52775, N52776, N52777, N52778, N52779, N52780, N52781, N52782, N52783, N52784, N52785, N52786, N52787, N52788, N52789, N52790, N52791, N52792, N52793, N52794, N52795, N52796, N52797, N52798, N52800, N52801, N52802, N52803, N52804, N52805, N52806, N52807, N52808, N52809, N52810, N52811, N52812, N52814, N52815, N52816, N52817, N52818, N52819, N52820, N52821, N52822, N52823, N52824, N52825, N52826, N52827, N52828, N52829, N52830, N52831, N52832, N52833, N52834, N52835, N52836, N52838, N52839, N52840, N52841, N52842, N52843, N52844, N52845, N52846, N52847, N52848, N52849, N52850, N52851, N52852, N52853, N52854, N52855, N52856, N52857, N52858, N52859, N52860, N52861, N52862, N52863, N52864, N52865, N52866, N52867, N52868, N52869, N52870, N52871, N52872, N52873, N52874, N52875, N52876, N52877, N52878, N52879, N52880, N52882, N52883, N52884, N52885, N52886, N52887, N52888, N52889, N52890, N52891, N52892, N52893, N52894, N52895, N52896, N52897, N52898, N52899, N52900, N52901, N52902, N52903, N52904, N52905, N52906, N52907, N52908, N52909, N52910, N52911, N52912, N52913, N52914, N52915, N52916, N52917, N52918, N52919, N52920, N52921, N52922, N52923, N52924, N52925, N52926, N52927, N52928, N52929, N52930, N52931, N52932, N52933, N52934, N52935, N52936, N52937, N52938, N52940, N52941, N52942, N52943, N52944, N52945, N52946, N52947, N52948, N52949, N52950, N52951, N52952, N52953, N52954, N52955, N52956, N52957, N52958, N52959, N52960, N52961, N52962, N52963, N52964, N52965, N52967, N52968, N52969, N52970, N52971, N52972, N52973, N52974, N52975, N52976, N52977, N52978, N52979, N52980, N52981, N52982, N52983, N52984, N52985, N52986, N52987, N52988, N52989, N52990, N52991, N52992, N52993, N52994, N52995, N52996, N52997, N52998, N52999, N53000, N53001, N53002, N53003, N53004, N53005, N53006, N53007, N53008, N53009, N53010, N53011, N53012, N53013, N53014, N53015, N53016, N53017, N53018, N53019, N53020, N53021, N53022, N53024, N53025, N53026, N53028, N53029, N53030, N53031, N53032, N53033, N53034, N53035, N53036, N53037, N53038, N53039, N53040, N53041, N53042, N53043, N53044, N53045, N53046, N53047, N53048, N53049, N53050, N53051, N53052, N53053, N53054, N53055, N53056, N53057, N53058, N53059, N53060, N53061, N53062, N53063, N53064, N53066, N53067, N53068, N53069, N53070, N53071, N53072, N53073, N53074, N53075, N53077, N53078, N53079, N53080, N53081, N53082, N53083, N53084, N53085, N53086, N53087, N53088, N53089, N53090, N53091, N53092, N53093, N53094, N53095, N53096, N53097, N53098, N53099, N53100, N53101, N53102, N53103, N53104, N53105, N53106, N53107, N53108, N53109, N53110, N53111, N53112, N53113, N53114, N53115, N53116, N53117, N53118, N53119, N53120, N53121, N53122, N53123, N53124, N53125, N53126, N53127, N53128, N53129, N53130, N53131, N53132, N53133, N53134, N53135, N53136, N53137, N53138, N53139, N53140, N53141, N53142, N53143, N53144, N53145, N53146, N53147, N53148, N53149, N53150, N53151, N53152, N53153, N53154, N53155, N53156, N53157, N53158, N53159, N53160, N53161, N53162, N53163, N53164, N53165, N53166, N53167, N53168, N53169, N53170, N53171, N53172, N53173, N53174, N53175, N53176, N53177, N53178, N53179, N53180, N53181, N53182, N53183, N53184, N53185, N53186, N53187, N53188, N53189, N53190, N53191, N53192, N53193, N53194, N53195, N53196, N53197, N53198, N53199, N53200, N53201, N53202, N53204, N53205, N53206, N53207, N53208, N53209, N53210, N53211, N53212, N53213, N53214, N53215, N53216, N53217, N53218, N53219, N53220, N53221, N53222, N53223, N53224, N53225, N53226, N53227, N53228, N53229, N53230, N53231, N53233, N53234, N53235, N53236, N53237, N53238, N53239, N53240, N53241, N53242, N53243, N53244, N53245, N53246, N53247, N53248, N53249, N53250, N53251, N53252, N53253, N53254, N53255, N53256, N53257, N53258, N53259, N53260, N53261, N53262, N53263, N53264, N53265, N53266, N53267, N53268, N53269, N53270, N53271, N53272, N53273, N53274, N53275, N53276, N53277, N53278, N53279, N53280, N53281, N53282, N53283, N53284, N53285, N53286, N53287, N53288, N53289, N53290, N53291, N53292, N53293, N53294, N53295, N53296, N53297, N53298, N53299, N53300, N53301, N53302, N53303, N53304, N53305, N53306, N53307, N53308, N53309, N53310, N53311, N53312, N53313, N53314, N53315, N53316, N53317, N53318, N53319, N53320, N53321, N53322, N53323, N53325, N53326, N53327, N53328, N53329, N53330, N53331, N53332, N53333, N53334, N53335, N53336, N53337, N53338, N53339, N53340, N53341, N53342, N53343, N53344, N53345, N53346, N53347, N53348, N53349, N53350, N53351, N53353, N53354, N53355, N53356, N53357, N53358, N53359, N53360, N53361, N53363, N53364, N53366, N53367, N53368, N53369, N53370, N53371, N53372, N53373, N53374, N53375, N53376, N53377, N53378, N53379, N53380, N53381, N53382, N53383, N53384, N53385, N53386, N53387, N53388, N53389, N53390, N53391, N53393, N53394, N53395, N53396, N53397, N53398, N53399, N53400, N53401, N53402, N53403, N53404, N53405, N53406, N53407, N53408, N53409, N53410, N53411, N53412, N53413, N53414, N53415, N53416, N53417, N53418, N53419, N53420, N53421, N53422, N53423, N53424, N53425, N53426, N53427, N53428, N53429, N53430, N53431, N53432, N53433, N53434, N53435, N53436, N53437, N53438, N53439, N53440, N53441, N53442, N53443, N53444, N53445, N53446, N53447, N53448, N53449, N53450, N53451, N53452, N53454, N53455, N53456, N53457, N53458, N53459, N53460, N53461, N53462, N53463, N53464, N53465, N53466, N53467, N53468, N53469, N53470, N53471, N53472, N53473, N53474, N53475, N53476, N53477, N53478, N53479, N53480, N53481, N53482, N53483, N53484, N53485, N53486, N53487, N53488, N53489, N53490, N53491, N53492, N53493, N53494, N53495, N53496, N53497, N53498, N53499, N53500, N53501, N53502, N53503, N53504, N53505, N53506, N53507, N53508, N53509, N53510, N53511, N53512, N53513, N53514, N53515, N53516, N53517, N53518, N53519, N53520, N53521, N53522, N53523, N53524, N53525, N53526, N53527, N53528, N53529, N53530, N53531, N53532, N53533, N53534, N53535, N53536, N53537, N53538, N53539, N53540, N53541, N53542, N53543, N53544, N53545, N53546, N53547, N53548, N53549, N53550, N53551, N53552, N53553, N53554, N53555, N53556, N53557, N53558, N53559, N53560, N53561, N53562, N53563, N53564, N53565, N53566, N53567, N53568, N53569, N53570, N53571, N53572, N53573, N53574, N53575, N53576, N53577, N53578, N53579, N53580, N53581, N53582, N53583, N53584, N53585, N53586, N53587, N53588, N53589, N53590, N53591, N53592, N53593, N53594, N53595, N53596, N53597, N53598, N53599, N53601, N53602, N53603, N53604, N53605, N53606, N53607, N53608, N53609, N53610, N53611, N53612, N53613, N53614, N53615, N53616, N53617, N53618, N53619, N53620, N53621, N53622, N53623, N53624, N53625, N53626, N53627, N53628, N53629, N53630, N53632, N53633, N53634, N53635, N53636, N53637, N53638, N53639, N53640, N53641, N53642, N53643, N53644, N53645, N53646, N53647, N53648, N53649, N53650, N53651, N53652, N53653, N53654, N53655, N53656, N53657, N53658, N53659, N53660, N53661, N53662, N53663, N53664, N53665, N53666, N53667, N53668, N53669, N53670, N53671, N53672, N53673, N53674, N53675, N53676, N53677, N53678, N53679, N53680, N53681, N53682, N53683, N53684, N53685, N53686, N53687, N53688, N53689, N53690, N53691, N53692, N53693, N53694, N53695, N53696, N53697, N53698, N53699, N53700, N53701, N53702, N53703, N53704, N53705, N53706, N53707, N53708, N53709, N53710, N53711, N53712, N53713, N53714, N53715, N53716, N53717, N53718, N53719, N53720, N53721, N53722, N53723, N53724, N53725, N53726, N53727, N53728, N53729, N53730, N53731, N53732, N53733, N53734, N53735, N53736, N53737, N53738, N53739, N53740, N53741, N53742, N53743, N53744, N53745, N53746, N53747, N53748, N53749, N53750, N53751, N53752, N53753, N53754, N53755, N53756, N53757, N53758, N53759, N53760, N53761, N53762, N53763, N53764, N53765, N53766, N53767, N53768, N53769, N53770, N53771, N53772, N53773, N53774, N53775, N53776, N53777, N53778, N53779, N53780, N53781, N53782, N53783, N53784, N53785, N53786, N53787, N53788, N53789, N53790, N53791, N53792, N53793, N53794, N53795, N53796, N53797, N53798, N53800, N53801, N53802, N53803, N53804, N53805, N53806, N53807, N53808, N53809, N53810, N53811, N53812, N53813, N53814, N53815, N53816, N53817, N53818, N53819, N53820, N53821, N53822, N53823, N53824, N53825, N53826, N53827, N53828, N53829, N53830, N53831, N53832, N53833, N53834, N53835, N53836, N53837, N53838, N53839, N53840, N53841, N53842, N53843, N53844, N53845, N53846, N53847, N53848, N53849, N53850, N53851, N53852, N53853, N53854, N53855, N53856, N53857, N53858, N53859, N53860, N53861, N53863, N53864, N53865, N53866, N53867, N53868, N53869, N53870, N53871, N53872, N53873, N53874, N53875, N53876, N53877, N53878, N53879, N53880, N53881, N53882, N53883, N53884, N53885, N53886, N53887, N53888, N53889, N53890, N53891, N53892, N53893, N53894, N53895, N53896, N53897, N53898, N53899, N53900, N53901, N53902, N53903, N53904, N53905, N53906, N53907, N53908, N53909, N53910, N53911, N53912, N53913, N53914, N53915, N53916, N53917, N53918, N53919, N53920, N53921, N53922, N53923, N53924, N53925, N53926, N53927, N53928, N53929, N53930, N53931, N53932, N53933, N53934, N53935, N53936, N53937, N53938, N53939, N53940, N53941, N53942, N53943, N53944, N53945, N53946, N53947, N53948, N53949, N53950, N53951, N53952, N53953, N53954, N53955, N53956, N53957, N53958, N53959, N53960, N53961, N53962, N53963, N53964, N53965, N53966, N53967, N53968, N53969, N53970, N53971, N53972, N53973, N53974, N53975, N53976, N53977, N53978, N53979, N53980, N53981, N53982, N53983, N53984, N53985, N53986, N53987, N53988, N53989, N53990, N53991, N53992, N53993, N53994, N53996, N53997, N53998, N53999, N54000, N54001, N54002, N54003, N54004, N54005, N54006, N54007, N54008, N54009, N54010, N54011, N54012, N54013, N54014, N54015, N54016, N54017, N54018, N54019, N54020, N54021, N54022, N54023, N54024, N54025, N54026, N54027, N54028, N54029, N54030, N54031, N54032, N54033, N54034, N54035, N54036, N54037, N54038, N54039, N54040, N54041, N54042, N54043, N54044, N54045, N54046, N54047, N54048, N54049, N54050, N54051, N54052, N54053, N54054, N54055, N54056, N54057, N54058, N54059, N54060, N54061, N54062, N54063, N54064, N54065, N54066, N54067, N54068, N54069, N54071, N54072, N54073, N54074, N54075, N54076, N54077, N54078, N54079, N54080, N54081, N54082, N54083, N54084, N54085, N54086, N54087, N54088, N54089, N54090, N54091, N54092, N54093, N54094, N54095, N54096, N54097, N54098, N54099, N54100, N54101, N54102, N54103, N54104, N54105, N54106, N54107, N54108, N54109, N54110, N54111, N54112, N54113, N54114, N54115, N54116, N54117, N54118, N54119, N54120, N54121, N54122, N54123, N54124, N54125, N54126, N54127, N54128, N54129, N54130, N54131, N54132, N54133, N54134, N54135, N54136, N54137, N54138, N54139, N54140, N54141, N54142, N54143, N54144, N54145, N54146, N54147, N54148, N54149, N54150, N54151, N54152, N54153, N54154, N54155, N54156, N54157, N54158, N54159, N54160, N54161, N54162, N54163, N54164, N54165, N54166, N54167, N54168, N54169, N54170, N54171, N54172, N54173, N54174, N54175, N54176, N54177, N54178, N54179, N54180, N54181, N54182, N54183, N54184, N54185, N54186, N54187, N54188, N54189, N54190, N54191, N54192, N54193, N54194, N54195, N54196, N54197, N54198, N54199, N54200, N54201, N54202, N54203, N54204, N54205, N54206, N54207, N54208, N54209, N54210, N54211, N54212, N54213, N54214, N54215, N54216, N54217, N54218, N54219, N54220, N54221, N54222, N54223, N54224, N54225, N54226, N54227, N54228, N54229, N54230, N54231, N54232, N54233, N54234, N54235, N54236, N54237, N54238, N54239, N54240, N54241, N54242, N54243, N54244, N54245, N54246, N54247, N54248, N54249, N54250, N54251, N54252, N54253, N54254, N54255, N54256, N54257, N54258, N54259, N54260, N54261, N54262, N54263, N54264, N54265, N54266, N54267, N54268, N54269, N54270, N54271, N54272, N54273, N54274, N54275, N54276, N54277, N54278, N54279, N54280, N54281, N54282, N54283, N54284, N54285, N54286, N54287, N54288, N54289, N54290, N54291, N54292, N54293, N54294, N54295, N54296, N54297, N54298, N54299, N54300, N54301, N54302, N54303, N54304, N54305, N54306, N54307, N54308, N54309, N54310, N54311, N54312, N54313, N54314, N54315, N54316, N54317, N54318, N54319, N54320, N54321);
    input N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413, N1414, N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503, N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513, N1514, N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563, N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612, N1613, N1614, N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664, N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734, N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804, N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1823, N1824, N1825, N1826, N1827, N1828, N1829, N1830, N1831, N1832, N1833, N1834, N1835, N1836, N1837, N1838, N1839, N1840, N1841, N1842, N1843, N1844, N1845, N1846, N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854, N1855, N1856, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1885, N1886, N1887, N1888, N1889, N1890, N1891, N1892, N1893, N1894, N1895, N1896, N1897, N1898, N1899, N1900, N1901, N1902, N1903, N1904, N1905, N1906, N1907, N1908, N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918, N1919, N1920, N1921, N1922, N1923, N1924, N1925, N1926, N1927, N1928, N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1947, N1948, N1949, N1950, N1951, N1952, N1953, N1954, N1955, N1956, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1964, N1965, N1966, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976, N1977, N1978, N1979, N1980, N1981, N1982, N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, N1991, N1992, N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, N2001, N2002, N2003, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044, N2045, N2046, N2047, N2048, N2049, N2050, N2051, N2052, N2053, N2054, N2055, N2056, N2057, N2058, N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079, N2080, N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2089, N2090, N2091, N2092, N2093, N2094, N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102, N2103, N2104, N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112, N2113, N2114, N2115, N2116, N2117, N2118, N2119, N2120, N2121, N2122, N2123, N2124, N2125, N2126, N2127, N2128, N2129, N2130, N2131, N2132, N2133, N2134, N2135, N2136, N2137, N2138, N2139, N2140, N2141, N2142, N2143, N2144, N2145, N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153, N2154, N2155, N2156, N2157, N2158, N2159, N2160, N2161, N2162, N2163, N2164, N2165, N2166, N2167, N2168, N2169, N2170, N2171, N2172, N2173, N2174, N2175, N2176, N2177, N2178, N2179, N2180, N2181, N2182, N2183, N2184, N2185, N2186, N2187, N2188, N2189, N2190, N2191, N2192, N2193, N2194, N2195, N2196, N2197, N2198, N2199, N2200, N2201, N2202, N2203, N2204, N2205, N2206, N2207, N2208, N2209, N2210, N2211, N2212, N2213, N2214, N2215, N2216, N2217, N2218, N2219, N2220, N2221, N2222, N2223, N2224, N2225, N2226, N2227, N2228, N2229, N2230, N2231, N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259, N2260, N2261, N2262, N2263, N2264, N2265, N2266, N2267, N2268, N2269, N2270, N2271, N2272, N2273, N2274, N2275, N2276, N2277, N2278, N2279, N2280, N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2288, N2289, N2290, N2291, N2292, N2293, N2294, N2295, N2296, N2297, N2298, N2299, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2369, N2370, N2371, N2372, N2373, N2374, N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393, N2394, N2395, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414, N2415, N2416, N2417, N2418, N2419, N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435, N2436, N2437, N2438, N2439, N2440, N2441, N2442, N2443, N2444, N2445, N2446, N2447, N2448, N2449, N2450, N2451, N2452, N2453, N2454, N2455, N2456, N2457, N2458, N2459, N2460, N2461, N2462, N2463, N2464, N2465, N2466, N2467, N2468, N2469, N2470, N2471, N2472, N2473, N2474, N2475, N2476, N2477, N2478, N2479, N2480, N2481, N2482, N2483, N2484, N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494, N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504, N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514, N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, N2542, N2543, N2544, N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2554, N2555, N2556, N2557, N2558, N2559, N2560, N2561, N2562, N2563, N2564, N2565, N2566, N2567, N2568, N2569, N2570, N2571, N2572, N2573, N2574, N2575, N2576, N2577, N2578, N2579, N2580, N2581, N2582, N2583, N2584, N2585, N2586, N2587, N2588, N2589, N2590, N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2623, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2648, N2649, N2650, N2651, N2652, N2653, N2654, N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2682, N2683, N2684, N2685, N2686, N2687, N2688, N2689, N2690, N2691, N2692, N2693, N2694, N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2704, N2705, N2706, N2707, N2708, N2709, N2710, N2711, N2712, N2713, N2714, N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2723, N2724, N2725, N2726, N2727, N2728, N2729, N2730, N2731, N2732, N2733, N2734, N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744, N2745, N2746, N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754, N2755, N2756, N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764, N2765, N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2788, N2789, N2790, N2791, N2792, N2793, N2794, N2795, N2796, N2797, N2798, N2799, N2800, N2801, N2802, N2803, N2804, N2805, N2806, N2807, N2808, N2809, N2810, N2811, N2812, N2813, N2814, N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859, N2860, N2861, N2862, N2863, N2864, N2865, N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, N3165, N3166, N3167, N3168, N3169, N3170, N3171, N3172, N3173, N3174, N3175, N3176, N3177, N3178, N3179, N3180, N3181, N3182, N3183, N3184, N3185, N3186, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196, N3197, N3198, N3199, N3200, N3201, N3202, N3203, N3204, N3205, N3206, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266, N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, N3338, N3339, N3340, N3341, N3342, N3343, N3344, N3345, N3346, N3347, N3348, N3349, N3350, N3351, N3352, N3353, N3354, N3355, N3356, N3357, N3358, N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3376, N3377, N3378, N3379, N3380, N3381, N3382, N3383, N3384, N3385, N3386, N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394, N3395, N3396, N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3417, N3418, N3419, N3420, N3421, N3422, N3423, N3424, N3425, N3426, N3427, N3428, N3429, N3430, N3431, N3432, N3433, N3434, N3435, N3436, N3437, N3438, N3439, N3440, N3441, N3442, N3443, N3444, N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, N3457, N3458, N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3467, N3468, N3469, N3470, N3471, N3472, N3473, N3474, N3475, N3476, N3477, N3478, N3479, N3480, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494, N3495, N3496, N3497, N3498, N3499, N3500, N3501, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514, N3515, N3516, N3517, N3518, N3519, N3520, N3521, N3522, N3523, N3524, N3525, N3526, N3527, N3528, N3529, N3530, N3531, N3532, N3533, N3534, N3535, N3536, N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544, N3545, N3546, N3547, N3548, N3549, N3550, N3551, N3552, N3553, N3554, N3555, N3556, N3557, N3558, N3559, N3560, N3561, N3562, N3563, N3564, N3565, N3566, N3567, N3568, N3569, N3570, N3571, N3572, N3573, N3574, N3575, N3576, N3577, N3578, N3579, N3580, N3581, N3582, N3583, N3584, N3585, N3586, N3587, N3588, N3589, N3590, N3591, N3592, N3593, N3594, N3595, N3596, N3597, N3598, N3599, N3600, N3601, N3602, N3603, N3604, N3605, N3606, N3607, N3608, N3609, N3610, N3611, N3612, N3613, N3614, N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3687, N3688, N3689, N3690, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3698, N3699, N3700, N3701, N3702, N3703, N3704, N3705, N3706, N3707, N3708, N3709, N3710, N3711, N3712, N3713, N3714, N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3733, N3734, N3735, N3736, N3737, N3738, N3739, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3772, N3773, N3774, N3775, N3776, N3777, N3778, N3779, N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, N3790, N3791, N3792, N3793, N3794, N3795, N3796, N3797, N3798, N3799, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, N3808, N3809, N3810, N3811, N3812, N3813, N3814, N3815, N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3823, N3824, N3825, N3826, N3827, N3828, N3829, N3830, N3831, N3832, N3833, N3834, N3835, N3836, N3837, N3838, N3839, N3840, N3841, N3842, N3843, N3844, N3845, N3846, N3847, N3848, N3849, N3850, N3851, N3852, N3853, N3854, N3855, N3856, N3857, N3858, N3859, N3860, N3861, N3862, N3863, N3864, N3865, N3866, N3867, N3868, N3869, N3870, N3871, N3872, N3873, N3874, N3875, N3876, N3877, N3878, N3879, N3880, N3881, N3882, N3883, N3884, N3885, N3886, N3887, N3888, N3889, N3890, N3891, N3892, N3893, N3894, N3895, N3896, N3897, N3898, N3899, N3900, N3901, N3902, N3903, N3904, N3905, N3906, N3907, N3908, N3909, N3910, N3911, N3912, N3913, N3914, N3915, N3916, N3917, N3918, N3919, N3920, N3921, N3922, N3923, N3924, N3925, N3926, N3927, N3928, N3929, N3930, N3931, N3932, N3933, N3934, N3935, N3936, N3937, N3938, N3939, N3940, N3941, N3942, N3943, N3944, N3945, N3946, N3947, N3948, N3949, N3950, N3951, N3952, N3953, N3954, N3955, N3956, N3957, N3958, N3959, N3960, N3961, N3962, N3963, N3964, N3965, N3966, N3967, N3968, N3969, N3970, N3971, N3972, N3973, N3974, N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3985, N3986, N3987, N3988, N3989, N3990, N3991, N3992, N3993, N3994, N3995, N3996, N3997, N3998, N3999, N4000, N4001, N4002, N4003, N4004, N4005, N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014, N4015, N4016, N4017, N4018, N4019, N4020, N4021, N4022, N4023, N4024, N4025, N4026, N4027, N4028, N4029, N4030, N4031, N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040, N4041, N4042, N4043, N4044, N4045, N4046, N4047, N4048, N4049, N4050, N4051, N4052, N4053, N4054, N4055, N4056, N4057, N4058, N4059, N4060, N4061, N4062, N4063, N4064, N4065, N4066, N4067, N4068, N4069, N4070, N4071, N4072, N4073, N4074, N4075, N4076, N4077, N4078, N4079, N4080, N4081, N4082, N4083, N4084, N4085, N4086, N4087, N4088, N4089, N4090, N4091, N4092, N4093, N4094, N4095, N4096, N4097, N4098, N4099, N4100, N4101, N4102, N4103, N4104, N4105, N4106, N4107, N4108, N4109, N4110, N4111, N4112, N4113, N4114, N4115, N4116, N4117, N4118, N4119, N4120, N4121, N4122, N4123, N4124, N4125, N4126, N4127, N4128, N4129, N4130, N4131, N4132, N4133, N4134, N4135, N4136, N4137, N4138, N4139, N4140, N4141, N4142, N4143, N4144, N4145, N4146, N4147, N4148, N4149, N4150, N4151, N4152, N4153, N4154, N4155, N4156, N4157, N4158, N4159, N4160, N4161, N4162, N4163, N4164, N4165, N4166, N4167, N4168, N4169, N4170, N4171, N4172, N4173, N4174, N4175, N4176, N4177, N4178, N4179, N4180, N4181, N4182, N4183, N4184, N4185, N4186, N4187, N4188, N4189, N4190, N4191, N4192, N4193, N4194, N4195, N4196, N4197, N4198, N4199, N4200, N4201, N4202, N4203, N4204, N4205, N4206, N4207, N4208, N4209, N4210, N4211, N4212, N4213, N4214, N4215, N4216, N4217, N4218, N4219, N4220, N4221, N4222, N4223, N4224, N4225, N4226, N4227, N4228, N4229, N4230, N4231, N4232, N4233, N4234, N4235, N4236, N4237, N4238, N4239, N4240, N4241, N4242, N4243, N4244, N4245, N4246, N4247, N4248, N4249, N4250, N4251, N4252, N4253, N4254, N4255, N4256, N4257, N4258, N4259, N4260, N4261, N4262, N4263, N4264, N4265, N4266, N4267, N4268, N4269, N4270, N4271, N4272, N4273, N4274, N4275, N4276, N4277, N4278, N4279, N4280, N4281, N4282, N4283, N4284, N4285, N4286, N4287, N4288, N4289, N4290, N4291, N4292, N4293, N4294, N4295, N4296, N4297, N4298, N4299, N4300, N4301, N4302, N4303, N4304, N4305, N4306, N4307, N4308, N4309, N4310, N4311, N4312, N4313, N4314, N4315, N4316, N4317, N4318, N4319, N4320, N4321, N4322, N4323, N4324, N4325, N4326, N4327, N4328, N4329, N4330, N4331, N4332, N4333, N4334, N4335, N4336, N4337, N4338, N4339, N4340, N4341, N4342, N4343, N4344, N4345, N4346, N4347, N4348, N4349, N4350, N4351, N4352, N4353, N4354, N4355, N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363, N4364, N4365, N4366, N4367, N4368, N4369, N4370, N4371, N4372, N4373, N4374, N4375, N4376, N4377, N4378, N4379, N4380, N4381, N4382, N4383, N4384, N4385, N4386, N4387, N4388, N4389, N4390, N4391, N4392, N4393, N4394, N4395, N4396, N4397, N4398, N4399, N4400, N4401, N4402, N4403, N4404, N4405, N4406, N4407, N4408, N4409, N4410, N4411, N4412, N4413, N4414, N4415, N4416, N4417, N4418, N4419, N4420, N4421, N4422, N4423, N4424, N4425, N4426, N4427, N4428, N4429, N4430, N4431, N4432, N4433, N4434, N4435, N4436, N4437, N4438, N4439, N4440, N4441, N4442, N4443, N4444, N4445, N4446, N4447, N4448, N4449, N4450, N4451, N4452, N4453, N4454, N4455, N4456, N4457, N4458, N4459, N4460, N4461, N4462, N4463, N4464, N4465, N4466, N4467, N4468, N4469, N4470, N4471, N4472, N4473, N4474, N4475, N4476, N4477, N4478, N4479, N4480, N4481, N4482, N4483, N4484, N4485, N4486, N4487, N4488, N4489, N4490, N4491, N4492, N4493, N4494, N4495, N4496, N4497, N4498, N4499, N4500, N4501, N4502, N4503, N4504, N4505, N4506, N4507, N4508, N4509, N4510, N4511, N4512, N4513, N4514, N4515, N4516, N4517, N4518, N4519, N4520, N4521, N4522, N4523, N4524, N4525, N4526, N4527, N4528, N4529, N4530, N4531, N4532, N4533, N4534, N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543, N4544, N4545, N4546, N4547, N4548, N4549, N4550, N4551, N4552, N4553, N4554, N4555, N4556, N4557, N4558, N4559, N4560, N4561, N4562, N4563, N4564, N4565, N4566, N4567, N4568, N4569, N4570, N4571, N4572, N4573, N4574, N4575, N4576, N4577, N4578, N4579, N4580, N4581, N4582, N4583, N4584, N4585, N4586, N4587, N4588, N4589, N4590, N4591, N4592, N4593, N4594, N4595, N4596, N4597, N4598, N4599, N4600, N4601, N4602, N4603, N4604, N4605, N4606, N4607, N4608, N4609, N4610, N4611, N4612, N4613, N4614, N4615, N4616, N4617, N4618, N4619, N4620, N4621, N4622, N4623, N4624, N4625, N4626, N4627, N4628, N4629, N4630, N4631, N4632, N4633, N4634, N4635, N4636, N4637, N4638, N4639, N4640, N4641, N4642, N4643, N4644, N4645, N4646, N4647, N4648, N4649, N4650, N4651, N4652, N4653, N4654, N4655, N4656, N4657, N4658, N4659, N4660, N4661, N4662, N4663, N4664, N4665, N4666, N4667, N4668, N4669, N4670, N4671, N4672, N4673, N4674, N4675, N4676, N4677, N4678, N4679, N4680, N4681, N4682, N4683, N4684, N4685, N4686, N4687, N4688, N4689, N4690, N4691, N4692, N4693, N4694, N4695, N4696, N4697, N4698, N4699, N4700, N4701, N4702, N4703, N4704, N4705, N4706, N4707, N4708, N4709, N4710, N4711, N4712, N4713, N4714, N4715, N4716, N4717, N4718, N4719, N4720, N4721, N4722, N4723, N4724, N4725, N4726, N4727, N4728, N4729, N4730, N4731, N4732, N4733, N4734, N4735, N4736, N4737, N4738, N4739, N4740, N4741, N4742, N4743, N4744, N4745, N4746, N4747, N4748, N4749, N4750, N4751, N4752, N4753, N4754, N4755, N4756, N4757, N4758, N4759, N4760, N4761, N4762, N4763, N4764, N4765, N4766, N4767, N4768, N4769, N4770, N4771, N4772, N4773, N4774, N4775, N4776, N4777, N4778, N4779, N4780, N4781, N4782, N4783, N4784, N4785, N4786, N4787, N4788, N4789, N4790, N4791, N4792, N4793, N4794, N4795, N4796, N4797, N4798, N4799, N4800, N4801, N4802, N4803, N4804, N4805, N4806, N4807, N4808, N4809, N4810, N4811, N4812, N4813, N4814, N4815, N4816, N4817, N4818, N4819, N4820, N4821, N4822, N4823, N4824, N4825, N4826, N4827, N4828, N4829, N4830, N4831, N4832, N4833, N4834, N4835, N4836, N4837, N4838, N4839, N4840, N4841, N4842, N4843, N4844, N4845, N4846, N4847, N4848, N4849, N4850, N4851, N4852, N4853, N4854, N4855, N4856, N4857, N4858, N4859, N4860, N4861, N4862, N4863, N4864, N4865, N4866, N4867, N4868, N4869, N4870, N4871, N4872, N4873, N4874, N4875, N4876, N4877, N4878, N4879, N4880, N4881, N4882, N4883, N4884, N4885, N4886, N4887, N4888, N4889, N4890, N4891, N4892, N4893, N4894, N4895, N4896, N4897, N4898, N4899, N4900, N4901, N4902, N4903, N4904, N4905, N4906, N4907, N4908, N4909, N4910, N4911, N4912, N4913, N4914, N4915, N4916, N4917, N4918, N4919, N4920, N4921, N4922, N4923, N4924, N4925, N4926, N4927, N4928, N4929, N4930, N4931, N4932, N4933, N4934, N4935, N4936, N4937, N4938, N4939, N4940, N4941, N4942, N4943, N4944, N4945, N4946, N4947, N4948, N4949, N4950, N4951, N4952, N4953, N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4962, N4963, N4964, N4965, N4966, N4967, N4968, N4969, N4970, N4971, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N4988, N4989, N4990, N4991, N4992, N4993, N4994, N4995, N4996, N4997, N4998, N4999, N5000, N5001, N5002, N5003, N5004, N5005, N5006, N5007, N5008, N5009, N5010, N5011, N5012, N5013, N5014, N5015, N5016, N5017, N5018, N5019, N5020, N5021, N5022, N5023, N5024, N5025, N5026, N5027, N5028, N5029, N5030, N5031, N5032, N5033, N5034, N5035, N5036, N5037, N5038, N5039, N5040, N5041, N5042, N5043, N5044, N5045, N5046, N5047, N5048, N5049, N5050, N5051, N5052, N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062, N5063, N5064, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5074, N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083, N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093, N5094, N5095, N5096, N5097, N5098, N5099, N5100, N5101, N5102, N5103, N5104, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113, N5114, N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123, N5124, N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, N5134, N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144, N5145, N5146, N5147, N5148, N5149, N5150, N5151, N5152, N5153, N5154, N5155, N5156, N5157, N5158, N5159, N5160, N5161, N5162, N5163, N5164, N5165, N5166, N5167, N5168, N5169, N5170, N5171, N5172, N5173, N5174, N5175, N5176, N5177, N5178, N5179, N5180, N5181, N5182, N5183, N5184, N5185, N5186, N5187, N5188, N5189, N5190, N5191, N5192, N5193, N5194, N5195, N5196, N5197, N5198, N5199, N5200, N5201, N5202, N5203, N5204, N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212, N5213, N5214, N5215, N5216, N5217, N5218, N5219, N5220, N5221, N5222, N5223, N5224, N5225, N5226, N5227, N5228, N5229, N5230, N5231, N5232, N5233, N5234, N5235, N5236, N5237, N5238, N5239, N5240, N5241, N5242, N5243, N5244, N5245, N5246, N5247, N5248, N5249, N5250, N5251, N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262, N5263, N5264, N5265, N5266, N5267, N5268, N5269, N5270, N5271, N5272, N5273, N5274, N5275, N5276, N5277, N5278, N5279, N5280, N5281, N5282, N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290, N5291, N5292, N5293, N5294, N5295, N5296, N5297, N5298, N5299, N5300, N5301, N5302, N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310, N5311, N5312, N5313, N5314, N5315, N5316, N5317, N5318, N5319, N5320, N5321, N5322, N5323, N5324, N5325, N5326, N5327, N5328, N5329, N5330, N5331, N5332, N5333, N5334, N5335, N5336, N5337, N5338, N5339, N5340, N5341, N5342, N5343, N5344, N5345, N5346, N5347, N5348, N5349, N5350, N5351, N5352, N5353, N5354, N5355, N5356, N5357, N5358, N5359, N5360, N5361, N5362, N5363, N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5372, N5373, N5374, N5375, N5376, N5377, N5378, N5379, N5380, N5381, N5382, N5383, N5384, N5385, N5386, N5387, N5388, N5389, N5390, N5391, N5392, N5393, N5394, N5395, N5396, N5397, N5398, N5399, N5400, N5401, N5402, N5403, N5404, N5405, N5406, N5407, N5408, N5409, N5410, N5411, N5412, N5413, N5414, N5415, N5416, N5417, N5418, N5419, N5420, N5421, N5422, N5423, N5424, N5425, N5426, N5427, N5428, N5429, N5430, N5431, N5432, N5433, N5434, N5435, N5436, N5437, N5438, N5439, N5440, N5441, N5442, N5443, N5444, N5445, N5446, N5447, N5448, N5449, N5450, N5451, N5452, N5453, N5454, N5455, N5456, N5457, N5458, N5459, N5460, N5461, N5462, N5463, N5464, N5465, N5466, N5467, N5468, N5469, N5470, N5471, N5472, N5473, N5474, N5475, N5476, N5477, N5478, N5479, N5480, N5481, N5482, N5483, N5484, N5485, N5486, N5487, N5488, N5489, N5490, N5491, N5492, N5493, N5494, N5495, N5496, N5497, N5498, N5499, N5500, N5501, N5502, N5503, N5504, N5505, N5506, N5507, N5508, N5509, N5510, N5511, N5512, N5513, N5514, N5515, N5516, N5517, N5518, N5519, N5520, N5521, N5522, N5523, N5524, N5525, N5526, N5527, N5528, N5529, N5530, N5531, N5532, N5533, N5534, N5535, N5536, N5537, N5538, N5539, N5540, N5541, N5542, N5543, N5544, N5545, N5546, N5547, N5548, N5549, N5550, N5551, N5552, N5553, N5554, N5555, N5556, N5557, N5558, N5559, N5560, N5561, N5562, N5563, N5564, N5565, N5566, N5567, N5568, N5569, N5570, N5571, N5572, N5573, N5574, N5575, N5576, N5577, N5578, N5579, N5580, N5581, N5582, N5583, N5584, N5585, N5586, N5587, N5588, N5589, N5590, N5591, N5592, N5593, N5594, N5595, N5596, N5597, N5598, N5599, N5600, N5601, N5602, N5603, N5604, N5605, N5606, N5607, N5608, N5609, N5610, N5611, N5612, N5613, N5614, N5615, N5616, N5617, N5618, N5619, N5620, N5621, N5622, N5623, N5624, N5625, N5626, N5627, N5628, N5629, N5630, N5631, N5632, N5633, N5634, N5635, N5636, N5637, N5638, N5639, N5640, N5641, N5642, N5643, N5644, N5645, N5646, N5647, N5648, N5649, N5650, N5651, N5652, N5653, N5654, N5655, N5656, N5657, N5658, N5659, N5660, N5661, N5662, N5663, N5664, N5665, N5666, N5667, N5668, N5669, N5670, N5671, N5672, N5673, N5674, N5675, N5676, N5677, N5678, N5679, N5680, N5681, N5682, N5683, N5684, N5685, N5686, N5687, N5688, N5689, N5690, N5691, N5692, N5693, N5694, N5695, N5696, N5697, N5698, N5699, N5700, N5701, N5702, N5703, N5704, N5705, N5706, N5707, N5708, N5709, N5710, N5711, N5712, N5713, N5714, N5715, N5716, N5717, N5718, N5719, N5720, N5721, N5722, N5723, N5724, N5725, N5726, N5727, N5728, N5729, N5730, N5731, N5732, N5733, N5734, N5735, N5736, N5737, N5738, N5739, N5740, N5741, N5742, N5743, N5744, N5745, N5746, N5747, N5748, N5749, N5750, N5751, N5752, N5753, N5754, N5755, N5756, N5757, N5758, N5759, N5760, N5761, N5762, N5763, N5764, N5765, N5766, N5767, N5768, N5769, N5770, N5771, N5772, N5773, N5774, N5775, N5776, N5777, N5778, N5779, N5780, N5781, N5782, N5783, N5784, N5785, N5786, N5787, N5788, N5789, N5790, N5791, N5792, N5793, N5794, N5795, N5796, N5797, N5798, N5799, N5800, N5801, N5802, N5803, N5804, N5805, N5806, N5807, N5808, N5809, N5810, N5811, N5812, N5813, N5814, N5815, N5816, N5817, N5818, N5819, N5820, N5821, N5822, N5823, N5824, N5825, N5826, N5827, N5828, N5829, N5830, N5831, N5832, N5833, N5834, N5835, N5836, N5837, N5838, N5839, N5840, N5841, N5842, N5843, N5844, N5845, N5846, N5847, N5848, N5849, N5850, N5851, N5852, N5853, N5854, N5855, N5856, N5857, N5858, N5859, N5860, N5861, N5862, N5863, N5864, N5865, N5866, N5867, N5868, N5869, N5870, N5871, N5872, N5873, N5874, N5875, N5876, N5877, N5878, N5879, N5880, N5881, N5882, N5883, N5884, N5885, N5886, N5887, N5888, N5889, N5890, N5891, N5892, N5893, N5894, N5895, N5896, N5897, N5898, N5899, N5900, N5901, N5902, N5903, N5904, N5905, N5906, N5907, N5908, N5909, N5910, N5911, N5912, N5913, N5914, N5915, N5916, N5917, N5918, N5919, N5920, N5921, N5922, N5923, N5924, N5925, N5926, N5927, N5928, N5929, N5930, N5931, N5932, N5933, N5934, N5935, N5936, N5937, N5938, N5939, N5940, N5941, N5942, N5943, N5944, N5945, N5946, N5947, N5948, N5949, N5950, N5951, N5952, N5953, N5954, N5955, N5956, N5957, N5958, N5959, N5960, N5961, N5962, N5963, N5964, N5965, N5966, N5967, N5968, N5969, N5970, N5971, N5972, N5973, N5974, N5975, N5976, N5977, N5978, N5979, N5980, N5981, N5982, N5983, N5984, N5985, N5986, N5987, N5988, N5989, N5990, N5991, N5992, N5993, N5994, N5995, N5996, N5997, N5998, N5999, N6000, N6001, N6002, N6003, N6004, N6005, N6006, N6007, N6008, N6009, N6010, N6011, N6012, N6013, N6014, N6015, N6016, N6017, N6018, N6019, N6020, N6021, N6022, N6023, N6024, N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032, N6033, N6034, N6035, N6036, N6037, N6038, N6039, N6040, N6041, N6042, N6043, N6044, N6045, N6046, N6047, N6048, N6049, N6050, N6051, N6052, N6053, N6054, N6055, N6056, N6057, N6058, N6059, N6060, N6061, N6062, N6063, N6064, N6065, N6066, N6067, N6068, N6069, N6070, N6071, N6072, N6073, N6074, N6075, N6076, N6077, N6078, N6079, N6080, N6081, N6082, N6083, N6084, N6085, N6086, N6087, N6088, N6089, N6090, N6091, N6092, N6093, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6109, N6110, N6111, N6112, N6113, N6114, N6115, N6116, N6117, N6118, N6119, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134, N6135, N6136, N6137, N6138, N6139, N6140, N6141, N6142, N6143, N6144, N6145, N6146, N6147, N6148, N6149, N6150, N6151, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6165, N6166, N6167, N6168, N6169, N6170, N6171, N6172, N6173, N6174, N6175, N6176, N6177, N6178, N6179, N6180, N6181, N6182, N6183, N6184, N6185, N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6195, N6196, N6197, N6198, N6199, N6200, N6201, N6202, N6203, N6204, N6205, N6206, N6207, N6208, N6209, N6210, N6211, N6212, N6213, N6214, N6215, N6216, N6217, N6218, N6219, N6220, N6221, N6222, N6223, N6224, N6225, N6226, N6227, N6228, N6229, N6230, N6231, N6232, N6233, N6234, N6235, N6236, N6237, N6238, N6239, N6240, N6241, N6242, N6243, N6244, N6245, N6246, N6247, N6248, N6249, N6250, N6251, N6252, N6253, N6254, N6255, N6256, N6257, N6258, N6259, N6260, N6261, N6262, N6263, N6264, N6265, N6266, N6267, N6268, N6269, N6270, N6271, N6272, N6273, N6274, N6275, N6276, N6277, N6278, N6279, N6280, N6281, N6282, N6283, N6284, N6285, N6286, N6287, N6288, N6289, N6290, N6291, N6292, N6293, N6294, N6295, N6296, N6297, N6298, N6299, N6300, N6301, N6302, N6303, N6304, N6305, N6306, N6307, N6308, N6309, N6310, N6311, N6312, N6313, N6314, N6315, N6316, N6317, N6318, N6319, N6320, N6321, N6322, N6323, N6324, N6325, N6326, N6327, N6328, N6329, N6330, N6331, N6332, N6333, N6334, N6335, N6336, N6337, N6338, N6339, N6340, N6341, N6342, N6343, N6344, N6345, N6346, N6347, N6348, N6349, N6350, N6351, N6352, N6353, N6354, N6355, N6356, N6357, N6358, N6359, N6360, N6361, N6362, N6363, N6364, N6365, N6366, N6367, N6368, N6369, N6370, N6371, N6372, N6373, N6374, N6375, N6376, N6377, N6378, N6379, N6380, N6381, N6382, N6383, N6384, N6385, N6386, N6387, N6388, N6389, N6390, N6391, N6392, N6393, N6394, N6395, N6396, N6397, N6398, N6399, N6400, N6401, N6402, N6403, N6404, N6405, N6406, N6407, N6408, N6409, N6410, N6411, N6412, N6413, N6414, N6415, N6416, N6417, N6418, N6419, N6420, N6421, N6422, N6423, N6424, N6425, N6426, N6427, N6428, N6429, N6430, N6431, N6432, N6433, N6434, N6435, N6436, N6437, N6438, N6439, N6440, N6441, N6442, N6443, N6444, N6445, N6446, N6447, N6448, N6449, N6450, N6451, N6452, N6453, N6454, N6455, N6456, N6457, N6458, N6459, N6460, N6461, N6462, N6463, N6464, N6465, N6466, N6467, N6468, N6469, N6470, N6471, N6472, N6473, N6474, N6475, N6476, N6477, N6478, N6479, N6480, N6481, N6482, N6483, N6484, N6485, N6486, N6487, N6488, N6489, N6490, N6491, N6492, N6493, N6494, N6495, N6496, N6497, N6498, N6499, N6500, N6501, N6502, N6503, N6504, N6505, N6506, N6507, N6508, N6509, N6510, N6511, N6512, N6513, N6514, N6515, N6516, N6517, N6518, N6519, N6520, N6521, N6522, N6523, N6524, N6525, N6526, N6527, N6528, N6529, N6530, N6531, N6532, N6533, N6534, N6535, N6536, N6537, N6538, N6539, N6540, N6541, N6542, N6543, N6544, N6545, N6546, N6547, N6548, N6549, N6550, N6551, N6552, N6553, N6554, N6555, N6556, N6557, N6558, N6559, N6560, N6561, N6562, N6563, N6564, N6565, N6566, N6567, N6568, N6569, N6570, N6571, N6572, N6573, N6574, N6575, N6576, N6577, N6578, N6579, N6580, N6581, N6582, N6583, N6584, N6585, N6586, N6587, N6588, N6589, N6590, N6591, N6592, N6593, N6594, N6595, N6596, N6597, N6598, N6599, N6600, N6601, N6602, N6603, N6604, N6605, N6606, N6607, N6608, N6609, N6610, N6611, N6612, N6613, N6614, N6615, N6616, N6617, N6618, N6619, N6620, N6621, N6622, N6623, N6624, N6625, N6626, N6627, N6628, N6629, N6630, N6631, N6632, N6633, N6634, N6635, N6636, N6637, N6638, N6639, N6640, N6641, N6642, N6643, N6644, N6645, N6646, N6647, N6648, N6649, N6650, N6651, N6652, N6653, N6654, N6655, N6656, N6657, N6658, N6659, N6660, N6661, N6662, N6663, N6664, N6665, N6666, N6667, N6668, N6669, N6670, N6671, N6672, N6673, N6674, N6675, N6676, N6677, N6678, N6679, N6680, N6681, N6682, N6683, N6684, N6685, N6686, N6687, N6688, N6689, N6690, N6691, N6692, N6693, N6694, N6695, N6696, N6697, N6698, N6699, N6700, N6701, N6702, N6703, N6704, N6705, N6706, N6707, N6708, N6709, N6710, N6711, N6712, N6713, N6714, N6715, N6716, N6717, N6718, N6719, N6720, N6721, N6722, N6723, N6724, N6725, N6726, N6727, N6728, N6729, N6730, N6731, N6732, N6733, N6734, N6735, N6736, N6737, N6738, N6739, N6740, N6741, N6742, N6743, N6744, N6745, N6746, N6747, N6748, N6749, N6750, N6751, N6752, N6753, N6754, N6755, N6756, N6757, N6758, N6759, N6760, N6761, N6762, N6763, N6764, N6765, N6766, N6767, N6768, N6769, N6770, N6771, N6772, N6773, N6774, N6775, N6776, N6777, N6778, N6779, N6780, N6781, N6782, N6783, N6784, N6785, N6786, N6787, N6788, N6789, N6790, N6791, N6792, N6793, N6794, N6795, N6796, N6797, N6798, N6799, N6800, N6801, N6802, N6803, N6804, N6805, N6806, N6807, N6808, N6809, N6810, N6811, N6812, N6813, N6814, N6815, N6816, N6817, N6818, N6819, N6820, N6821, N6822, N6823, N6824, N6825, N6826, N6827, N6828, N6829, N6830, N6831, N6832, N6833, N6834, N6835, N6836, N6837, N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6845, N6846, N6847, N6848, N6849, N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857, N6858, N6859, N6860, N6861, N6862, N6863, N6864, N6865, N6866, N6867, N6868, N6869, N6870, N6871, N6872, N6873, N6874, N6875, N6876, N6877, N6878, N6879, N6880, N6881, N6882, N6883, N6884, N6885, N6886, N6887, N6888, N6889, N6890, N6891, N6892, N6893, N6894, N6895, N6896, N6897, N6898, N6899, N6900, N6901, N6902, N6903, N6904, N6905, N6906, N6907, N6908, N6909, N6910, N6911, N6912, N6913, N6914, N6915, N6916, N6917, N6918, N6919, N6920, N6921, N6922, N6923, N6924, N6925, N6926, N6927, N6928, N6929, N6930, N6931, N6932, N6933, N6934, N6935, N6936, N6937, N6938, N6939, N6940, N6941, N6942, N6943, N6944, N6945, N6946, N6947, N6948, N6949, N6950, N6951, N6952, N6953, N6954, N6955, N6956, N6957, N6958, N6959, N6960, N6961, N6962, N6963, N6964, N6965, N6966, N6967, N6968, N6969, N6970, N6971, N6972, N6973, N6974, N6975, N6976, N6977, N6978, N6979, N6980, N6981, N6982, N6983, N6984, N6985, N6986, N6987, N6988, N6989, N6990, N6991, N6992, N6993, N6994, N6995, N6996, N6997, N6998, N6999, N7000, N7001, N7002, N7003, N7004, N7005, N7006, N7007, N7008, N7009, N7010, N7011, N7012, N7013, N7014, N7015, N7016, N7017, N7018, N7019, N7020, N7021, N7022, N7023, N7024, N7025, N7026, N7027, N7028, N7029, N7030, N7031, N7032, N7033, N7034, N7035, N7036, N7037, N7038, N7039, N7040, N7041, N7042, N7043, N7044, N7045, N7046, N7047, N7048, N7049, N7050, N7051, N7052, N7053, N7054, N7055, N7056, N7057, N7058, N7059, N7060, N7061, N7062, N7063, N7064, N7065, N7066, N7067, N7068, N7069, N7070, N7071, N7072, N7073, N7074, N7075, N7076, N7077, N7078, N7079, N7080, N7081, N7082, N7083, N7084, N7085, N7086, N7087, N7088, N7089, N7090, N7091, N7092, N7093, N7094, N7095, N7096, N7097, N7098, N7099, N7100, N7101, N7102, N7103, N7104, N7105, N7106, N7107, N7108, N7109, N7110, N7111, N7112, N7113, N7114, N7115, N7116, N7117, N7118, N7119, N7120, N7121, N7122, N7123, N7124, N7125, N7126, N7127, N7128, N7129, N7130, N7131, N7132, N7133, N7134, N7135, N7136, N7137, N7138, N7139, N7140, N7141, N7142, N7143, N7144, N7145, N7146, N7147, N7148, N7149, N7150, N7151, N7152, N7153, N7154, N7155, N7156, N7157, N7158, N7159, N7160, N7161, N7162, N7163, N7164, N7165, N7166, N7167, N7168, N7169, N7170, N7171, N7172, N7173, N7174, N7175, N7176, N7177, N7178, N7179, N7180, N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188, N7189, N7190, N7191, N7192, N7193, N7194, N7195, N7196, N7197, N7198, N7199, N7200, N7201, N7202, N7203, N7204, N7205, N7206, N7207, N7208, N7209, N7210, N7211, N7212, N7213, N7214, N7215, N7216, N7217, N7218, N7219, N7220, N7221, N7222, N7223, N7224, N7225, N7226, N7227, N7228, N7229, N7230, N7231, N7232, N7233, N7234, N7235, N7236, N7237, N7238, N7239, N7240, N7241, N7242, N7243, N7244, N7245, N7246, N7247, N7248, N7249, N7250, N7251, N7252, N7253, N7254, N7255, N7256, N7257, N7258, N7259, N7260, N7261, N7262, N7263, N7264, N7265, N7266, N7267, N7268, N7269, N7270, N7271, N7272, N7273, N7274, N7275, N7276, N7277, N7278, N7279, N7280, N7281, N7282, N7283, N7284, N7285, N7286, N7287, N7288, N7289, N7290, N7291, N7292, N7293, N7294, N7295, N7296, N7297, N7298, N7299, N7300, N7301, N7302, N7303, N7304, N7305, N7306, N7307, N7308, N7309, N7310, N7311, N7312, N7313, N7314, N7315, N7316, N7317, N7318, N7319, N7320, N7321, N7322, N7323, N7324, N7325, N7326, N7327, N7328, N7329, N7330, N7331, N7332, N7333, N7334, N7335, N7336, N7337, N7338, N7339, N7340, N7341, N7342, N7343, N7344, N7345, N7346, N7347, N7348, N7349, N7350, N7351, N7352, N7353, N7354, N7355, N7356, N7357, N7358, N7359, N7360, N7361, N7362, N7363, N7364, N7365, N7366, N7367, N7368, N7369, N7370, N7371, N7372, N7373, N7374, N7375, N7376, N7377, N7378, N7379, N7380, N7381, N7382, N7383, N7384, N7385, N7386, N7387, N7388, N7389, N7390, N7391, N7392, N7393, N7394, N7395, N7396, N7397, N7398, N7399, N7400, N7401, N7402, N7403, N7404, N7405, N7406, N7407, N7408, N7409, N7410, N7411, N7412, N7413, N7414, N7415, N7416, N7417, N7418, N7419, N7420, N7421, N7422, N7423, N7424, N7425, N7426, N7427, N7428, N7429, N7430, N7431, N7432, N7433, N7434, N7435, N7436, N7437, N7438, N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447, N7448, N7449, N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7457, N7458, N7459, N7460, N7461, N7462, N7463, N7464, N7465, N7466, N7467, N7468, N7469, N7470, N7471, N7472, N7473, N7474, N7475, N7476, N7477, N7478, N7479, N7480, N7481, N7482, N7483, N7484, N7485, N7486, N7487, N7488, N7489, N7490, N7491, N7492, N7493, N7494, N7495, N7496, N7497, N7498, N7499, N7500, N7501, N7502, N7503, N7504, N7505, N7506, N7507, N7508, N7509, N7510, N7511, N7512, N7513, N7514, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7523, N7524, N7525, N7526, N7527, N7528, N7529, N7530, N7531, N7532, N7533, N7534, N7535, N7536, N7537, N7538, N7539, N7540, N7541, N7542, N7543, N7544, N7545, N7546, N7547, N7548, N7549, N7550, N7551, N7552, N7553, N7554, N7555, N7556, N7557, N7558, N7559, N7560, N7561, N7562, N7563, N7564, N7565, N7566, N7567, N7568, N7569, N7570, N7571, N7572, N7573, N7574, N7575, N7576, N7577, N7578, N7579, N7580, N7581, N7582, N7583, N7584, N7585, N7586, N7587, N7588, N7589, N7590, N7591, N7592, N7593, N7594, N7595, N7596, N7597, N7598, N7599, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7608, N7609, N7610, N7611, N7612, N7613, N7614, N7615, N7616, N7617, N7618, N7619, N7620, N7621, N7622, N7623, N7624, N7625, N7626, N7627, N7628, N7629, N7630, N7631, N7632, N7633, N7634, N7635, N7636, N7637, N7638, N7639, N7640, N7641, N7642, N7643, N7644, N7645, N7646, N7647, N7648, N7649, N7650, N7651, N7652, N7653, N7654, N7655, N7656, N7657, N7658, N7659, N7660, N7661, N7662, N7663, N7664, N7665, N7666, N7667, N7668, N7669, N7670, N7671, N7672, N7673, N7674, N7675, N7676, N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684, N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692, N7693, N7694, N7695, N7696, N7697, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7708, N7709, N7710, N7711, N7712, N7713, N7714, N7715, N7716, N7717, N7718, N7719, N7720, N7721, N7722, N7723, N7724, N7725, N7726, N7727, N7728, N7729, N7730, N7731, N7732, N7733, N7734, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7743, N7744, N7745, N7746, N7747, N7748, N7749, N7750, N7751, N7752, N7753, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N7762, N7763, N7764, N7765, N7766, N7767, N7768, N7769, N7770, N7771, N7772, N7773, N7774, N7775, N7776, N7777, N7778, N7779, N7780, N7781, N7782, N7783, N7784, N7785, N7786, N7787, N7788, N7789, N7790, N7791, N7792, N7793, N7794, N7795, N7796, N7797, N7798, N7799, N7800, N7801, N7802, N7803, N7804, N7805, N7806, N7807, N7808, N7809, N7810, N7811, N7812, N7813, N7814, N7815, N7816, N7817, N7818, N7819, N7820, N7821, N7822, N7823, N7824, N7825, N7826, N7827, N7828, N7829, N7830, N7831, N7832, N7833, N7834, N7835, N7836, N7837, N7838, N7839, N7840, N7841, N7842, N7843, N7844, N7845, N7846, N7847, N7848, N7849, N7850, N7851, N7852, N7853, N7854, N7855, N7856, N7857, N7858, N7859, N7860, N7861, N7862, N7863, N7864, N7865, N7866, N7867, N7868, N7869, N7870, N7871, N7872, N7873, N7874, N7875, N7876, N7877, N7878, N7879, N7880, N7881, N7882, N7883, N7884, N7885, N7886, N7887, N7888, N7889, N7890, N7891, N7892, N7893, N7894, N7895, N7896, N7897, N7898, N7899, N7900, N7901, N7902, N7903, N7904, N7905, N7906, N7907, N7908, N7909, N7910, N7911, N7912, N7913, N7914, N7915, N7916, N7917, N7918, N7919, N7920, N7921, N7922, N7923, N7924, N7925, N7926, N7927, N7928, N7929, N7930, N7931, N7932, N7933, N7934, N7935, N7936, N7937, N7938, N7939, N7940, N7941, N7942, N7943, N7944, N7945, N7946, N7947, N7948, N7949, N7950, N7951, N7952, N7953, N7954, N7955, N7956, N7957, N7958, N7959, N7960, N7961, N7962, N7963, N7964, N7965, N7966, N7967, N7968, N7969, N7970, N7971, N7972, N7973, N7974, N7975, N7976, N7977, N7978, N7979, N7980, N7981, N7982, N7983, N7984, N7985, N7986, N7987, N7988, N7989, N7990, N7991, N7992, N7993, N7994, N7995, N7996, N7997, N7998, N7999, N8000, N8001, N8002, N8003, N8004, N8005, N8006, N8007, N8008, N8009, N8010, N8011, N8012, N8013, N8014, N8015, N8016, N8017, N8018, N8019, N8020, N8021, N8022, N8023, N8024, N8025, N8026, N8027, N8028, N8029, N8030, N8031, N8032, N8033, N8034, N8035, N8036, N8037, N8038, N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8046, N8047, N8048, N8049, N8050, N8051, N8052, N8053, N8054, N8055, N8056, N8057, N8058, N8059, N8060, N8061, N8062, N8063, N8064, N8065, N8066, N8067, N8068, N8069, N8070, N8071, N8072, N8073, N8074, N8075, N8076, N8077, N8078, N8079, N8080, N8081, N8082, N8083, N8084, N8085, N8086, N8087, N8088, N8089, N8090, N8091, N8092, N8093, N8094, N8095, N8096, N8097, N8098, N8099, N8100, N8101, N8102, N8103, N8104, N8105, N8106, N8107, N8108, N8109, N8110, N8111, N8112, N8113, N8114, N8115, N8116, N8117, N8118, N8119, N8120, N8121, N8122, N8123, N8124, N8125, N8126, N8127, N8128, N8129, N8130, N8131, N8132, N8133, N8134, N8135, N8136, N8137, N8138, N8139, N8140, N8141, N8142, N8143, N8144, N8145, N8146, N8147, N8148, N8149, N8150, N8151, N8152, N8153, N8154, N8155, N8156, N8157, N8158, N8159, N8160, N8161, N8162, N8163, N8164, N8165, N8166, N8167, N8168, N8169, N8170, N8171, N8172, N8173, N8174, N8175, N8176, N8177, N8178, N8179, N8180, N8181, N8182, N8183, N8184, N8185, N8186, N8187, N8188, N8189, N8190, N8191, N8192, N8193, N8194, N8195, N8196, N8197, N8198, N8199, N8200, N8201, N8202, N8203, N8204, N8205, N8206, N8207, N8208, N8209, N8210, N8211, N8212, N8213, N8214, N8215, N8216, N8217, N8218, N8219, N8220, N8221, N8222, N8223, N8224, N8225, N8226, N8227, N8228, N8229, N8230, N8231, N8232, N8233, N8234, N8235, N8236, N8237, N8238, N8239, N8240, N8241, N8242, N8243, N8244, N8245, N8246, N8247, N8248, N8249, N8250, N8251, N8252, N8253, N8254, N8255, N8256, N8257, N8258, N8259, N8260, N8261, N8262, N8263, N8264, N8265, N8266, N8267, N8268, N8269, N8270, N8271, N8272, N8273, N8274, N8275, N8276, N8277, N8278, N8279, N8280, N8281, N8282, N8283, N8284, N8285, N8286, N8287, N8288, N8289, N8290, N8291, N8292, N8293, N8294, N8295, N8296, N8297, N8298, N8299, N8300, N8301, N8302, N8303, N8304, N8305, N8306, N8307, N8308, N8309, N8310, N8311, N8312, N8313, N8314, N8315, N8316, N8317, N8318, N8319, N8320, N8321, N8322, N8323, N8324, N8325, N8326, N8327, N8328, N8329, N8330, N8331, N8332, N8333, N8334, N8335, N8336, N8337, N8338, N8339, N8340, N8341, N8342, N8343, N8344, N8345, N8346, N8347, N8348, N8349, N8350, N8351, N8352, N8353, N8354, N8355, N8356, N8357, N8358, N8359, N8360, N8361, N8362, N8363, N8364, N8365, N8366, N8367, N8368, N8369, N8370, N8371, N8372, N8373, N8374, N8375, N8376, N8377, N8378, N8379, N8380, N8381, N8382, N8383, N8384, N8385, N8386, N8387, N8388, N8389, N8390, N8391, N8392, N8393, N8394, N8395, N8396, N8397, N8398, N8399, N8400, N8401, N8402, N8403, N8404, N8405, N8406, N8407, N8408, N8409, N8410, N8411, N8412, N8413, N8414, N8415, N8416, N8417, N8418, N8419, N8420, N8421, N8422, N8423, N8424, N8425, N8426, N8427, N8428, N8429, N8430, N8431, N8432, N8433, N8434, N8435, N8436, N8437, N8438, N8439, N8440, N8441, N8442, N8443, N8444, N8445, N8446, N8447, N8448, N8449, N8450, N8451, N8452, N8453, N8454, N8455, N8456, N8457, N8458, N8459, N8460, N8461, N8462, N8463, N8464, N8465, N8466, N8467, N8468, N8469, N8470, N8471, N8472, N8473, N8474, N8475, N8476, N8477, N8478, N8479, N8480, N8481, N8482, N8483, N8484, N8485, N8486, N8487, N8488, N8489, N8490, N8491, N8492, N8493, N8494, N8495, N8496, N8497, N8498, N8499, N8500, N8501, N8502, N8503, N8504, N8505, N8506, N8507, N8508, N8509, N8510, N8511, N8512, N8513, N8514, N8515, N8516, N8517, N8518, N8519, N8520, N8521, N8522, N8523, N8524, N8525, N8526, N8527, N8528, N8529, N8530, N8531, N8532, N8533, N8534, N8535, N8536, N8537, N8538, N8539, N8540, N8541, N8542, N8543, N8544, N8545, N8546, N8547, N8548, N8549, N8550, N8551, N8552, N8553, N8554, N8555, N8556, N8557, N8558, N8559, N8560, N8561, N8562, N8563, N8564, N8565, N8566, N8567, N8568, N8569, N8570, N8571, N8572, N8573, N8574, N8575, N8576, N8577, N8578, N8579, N8580, N8581, N8582, N8583, N8584, N8585, N8586, N8587, N8588, N8589, N8590, N8591, N8592, N8593, N8594, N8595, N8596, N8597, N8598, N8599, N8600, N8601, N8602, N8603, N8604, N8605, N8606, N8607, N8608, N8609, N8610, N8611, N8612, N8613, N8614, N8615, N8616, N8617, N8618, N8619, N8620, N8621, N8622, N8623, N8624, N8625, N8626, N8627, N8628, N8629, N8630, N8631, N8632, N8633, N8634, N8635, N8636, N8637, N8638, N8639, N8640, N8641, N8642, N8643, N8644, N8645, N8646, N8647, N8648, N8649, N8650, N8651, N8652, N8653, N8654, N8655, N8656, N8657, N8658, N8659, N8660, N8661, N8662, N8663, N8664, N8665, N8666, N8667, N8668, N8669, N8670, N8671, N8672, N8673, N8674, N8675, N8676, N8677, N8678, N8679, N8680, N8681, N8682, N8683, N8684, N8685, N8686, N8687, N8688, N8689, N8690, N8691, N8692, N8693, N8694, N8695, N8696, N8697, N8698, N8699, N8700, N8701, N8702, N8703, N8704, N8705, N8706, N8707, N8708, N8709, N8710, N8711, N8712, N8713, N8714, N8715, N8716, N8717, N8718, N8719, N8720, N8721, N8722, N8723, N8724, N8725, N8726, N8727, N8728, N8729, N8730, N8731, N8732, N8733, N8734, N8735, N8736, N8737, N8738, N8739, N8740, N8741, N8742, N8743, N8744, N8745, N8746, N8747, N8748, N8749, N8750, N8751, N8752, N8753, N8754, N8755, N8756, N8757, N8758, N8759, N8760, N8761, N8762, N8763, N8764, N8765, N8766, N8767, N8768, N8769, N8770, N8771, N8772, N8773, N8774, N8775, N8776, N8777, N8778, N8779, N8780, N8781, N8782, N8783, N8784, N8785, N8786, N8787, N8788, N8789, N8790, N8791, N8792, N8793, N8794, N8795, N8796, N8797, N8798, N8799, N8800, N8801, N8802, N8803, N8804, N8805, N8806, N8807, N8808, N8809, N8810, N8811, N8812, N8813, N8814, N8815, N8816, N8817, N8818, N8819, N8820, N8821, N8822, N8823, N8824, N8825, N8826, N8827, N8828, N8829, N8830, N8831, N8832, N8833, N8834, N8835, N8836, N8837, N8838, N8839, N8840, N8841, N8842, N8843, N8844, N8845, N8846, N8847, N8848, N8849, N8850, N8851, N8852, N8853, N8854, N8855, N8856, N8857, N8858, N8859, N8860, N8861, N8862, N8863, N8864, N8865, N8866, N8867, N8868, N8869, N8870, N8871, N8872, N8873, N8874, N8875, N8876, N8877, N8878, N8879, N8880, N8881, N8882, N8883, N8884, N8885, N8886, N8887, N8888, N8889, N8890, N8891, N8892, N8893, N8894, N8895, N8896, N8897, N8898, N8899, N8900, N8901, N8902, N8903, N8904, N8905, N8906, N8907, N8908, N8909, N8910, N8911, N8912, N8913, N8914, N8915, N8916, N8917, N8918, N8919, N8920, N8921, N8922, N8923, N8924, N8925, N8926, N8927, N8928, N8929, N8930, N8931, N8932, N8933, N8934, N8935, N8936, N8937, N8938, N8939, N8940, N8941, N8942, N8943, N8944, N8945, N8946, N8947, N8948, N8949, N8950, N8951, N8952, N8953, N8954, N8955, N8956, N8957, N8958, N8959, N8960, N8961, N8962, N8963, N8964, N8965, N8966, N8967, N8968, N8969, N8970, N8971, N8972, N8973, N8974, N8975, N8976, N8977, N8978, N8979, N8980, N8981, N8982, N8983, N8984, N8985, N8986, N8987, N8988, N8989, N8990, N8991, N8992, N8993, N8994, N8995, N8996, N8997, N8998, N8999, N9000, N9001, N9002, N9003, N9004, N9005, N9006, N9007, N9008, N9009, N9010, N9011, N9012, N9013, N9014, N9015, N9016, N9017, N9018, N9019, N9020, N9021, N9022, N9023, N9024, N9025, N9026, N9027, N9028, N9029, N9030, N9031, N9032, N9033, N9034, N9035, N9036, N9037, N9038, N9039, N9040, N9041, N9042, N9043, N9044, N9045, N9046, N9047, N9048, N9049, N9050, N9051, N9052, N9053, N9054, N9055, N9056, N9057, N9058, N9059, N9060, N9061, N9062, N9063, N9064, N9065, N9066, N9067, N9068, N9069, N9070, N9071, N9072, N9073, N9074, N9075, N9076, N9077, N9078, N9079, N9080, N9081, N9082, N9083, N9084, N9085, N9086, N9087, N9088, N9089, N9090, N9091, N9092, N9093, N9094, N9095, N9096, N9097, N9098, N9099, N9100, N9101, N9102, N9103, N9104, N9105, N9106, N9107, N9108, N9109, N9110, N9111, N9112, N9113, N9114, N9115, N9116, N9117, N9118, N9119, N9120, N9121, N9122, N9123, N9124, N9125, N9126, N9127, N9128, N9129, N9130, N9131, N9132, N9133, N9134, N9135, N9136, N9137, N9138, N9139, N9140, N9141, N9142, N9143, N9144, N9145, N9146, N9147, N9148, N9149, N9150, N9151, N9152, N9153, N9154, N9155, N9156, N9157, N9158, N9159, N9160, N9161, N9162, N9163, N9164, N9165, N9166, N9167, N9168, N9169, N9170, N9171, N9172, N9173, N9174, N9175, N9176, N9177, N9178, N9179, N9180, N9181, N9182, N9183, N9184, N9185, N9186, N9187, N9188, N9189, N9190, N9191, N9192, N9193, N9194, N9195, N9196, N9197, N9198, N9199, N9200, N9201, N9202, N9203, N9204, N9205, N9206, N9207, N9208, N9209, N9210, N9211, N9212, N9213, N9214, N9215, N9216, N9217, N9218, N9219, N9220, N9221, N9222, N9223, N9224, N9225, N9226, N9227, N9228, N9229, N9230, N9231, N9232, N9233, N9234, N9235, N9236, N9237, N9238, N9239, N9240, N9241, N9242, N9243, N9244, N9245, N9246, N9247, N9248, N9249, N9250, N9251, N9252, N9253, N9254, N9255, N9256, N9257, N9258, N9259, N9260, N9261, N9262, N9263, N9264, N9265, N9266, N9267, N9268, N9269, N9270, N9271, N9272, N9273, N9274, N9275, N9276, N9277, N9278, N9279, N9280, N9281, N9282, N9283, N9284, N9285, N9286, N9287, N9288, N9289, N9290, N9291, N9292, N9293, N9294, N9295, N9296, N9297, N9298, N9299, N9300, N9301, N9302, N9303, N9304, N9305, N9306, N9307, N9308, N9309, N9310, N9311, N9312, N9313, N9314, N9315, N9316, N9317, N9318, N9319, N9320, N9321, N9322, N9323, N9324, N9325, N9326, N9327, N9328, N9329, N9330, N9331, N9332, N9333, N9334, N9335, N9336, N9337, N9338, N9339, N9340, N9341, N9342, N9343, N9344, N9345, N9346, N9347, N9348, N9349, N9350, N9351, N9352, N9353, N9354, N9355, N9356, N9357, N9358, N9359, N9360, N9361, N9362, N9363, N9364, N9365, N9366, N9367, N9368, N9369, N9370, N9371, N9372, N9373, N9374, N9375, N9376, N9377, N9378, N9379, N9380, N9381, N9382, N9383, N9384, N9385, N9386, N9387, N9388, N9389, N9390, N9391, N9392, N9393, N9394, N9395, N9396, N9397, N9398, N9399, N9400, N9401, N9402, N9403, N9404, N9405, N9406, N9407, N9408, N9409, N9410, N9411, N9412, N9413, N9414, N9415, N9416, N9417, N9418, N9419, N9420, N9421, N9422, N9423, N9424, N9425, N9426, N9427, N9428, N9429, N9430, N9431, N9432, N9433, N9434, N9435, N9436, N9437, N9438, N9439, N9440, N9441, N9442, N9443, N9444, N9445, N9446, N9447, N9448, N9449, N9450, N9451, N9452, N9453, N9454, N9455, N9456, N9457, N9458, N9459, N9460, N9461, N9462, N9463, N9464, N9465, N9466, N9467, N9468, N9469, N9470, N9471, N9472, N9473, N9474, N9475, N9476, N9477, N9478, N9479, N9480, N9481, N9482, N9483, N9484, N9485, N9486, N9487, N9488, N9489, N9490, N9491, N9492, N9493, N9494, N9495, N9496, N9497, N9498, N9499, N9500, N9501, N9502, N9503, N9504, N9505, N9506, N9507, N9508, N9509, N9510, N9511, N9512, N9513, N9514, N9515, N9516, N9517, N9518, N9519, N9520, N9521, N9522, N9523, N9524, N9525, N9526, N9527, N9528, N9529, N9530, N9531, N9532, N9533, N9534, N9535, N9536, N9537, N9538, N9539, N9540, N9541, N9542, N9543, N9544, N9545, N9546, N9547, N9548, N9549, N9550, N9551, N9552, N9553, N9554, N9555, N9556, N9557, N9558, N9559, N9560, N9561, N9562, N9563, N9564, N9565, N9566, N9567, N9568, N9569, N9570, N9571, N9572, N9573, N9574, N9575, N9576, N9577, N9578, N9579, N9580, N9581, N9582, N9583, N9584, N9585, N9586, N9587, N9588, N9589, N9590, N9591, N9592, N9593, N9594, N9595, N9596, N9597, N9598, N9599, N9600, N9601, N9602, N9603, N9604, N9605, N9606, N9607, N9608, N9609, N9610, N9611, N9612, N9613, N9614, N9615, N9616, N9617, N9618, N9619, N9620, N9621, N9622, N9623, N9624, N9625, N9626, N9627, N9628, N9629, N9630, N9631, N9632, N9633, N9634, N9635, N9636, N9637, N9638, N9639, N9640, N9641, N9642, N9643, N9644, N9645, N9646, N9647, N9648, N9649, N9650, N9651, N9652, N9653, N9654, N9655, N9656, N9657, N9658, N9659, N9660, N9661, N9662, N9663, N9664, N9665, N9666, N9667, N9668, N9669, N9670, N9671, N9672, N9673, N9674, N9675, N9676, N9677, N9678, N9679, N9680, N9681, N9682, N9683, N9684, N9685, N9686, N9687, N9688, N9689, N9690, N9691, N9692, N9693, N9694, N9695, N9696, N9697, N9698, N9699, N9700, N9701, N9702, N9703, N9704, N9705, N9706, N9707, N9708, N9709, N9710, N9711, N9712, N9713, N9714, N9715, N9716, N9717, N9718, N9719, N9720, N9721, N9722, N9723, N9724, N9725, N9726, N9727, N9728, N9729, N9730, N9731, N9732, N9733, N9734, N9735, N9736, N9737, N9738, N9739, N9740, N9741, N9742, N9743, N9744, N9745, N9746, N9747, N9748, N9749, N9750, N9751, N9752, N9753, N9754, N9755, N9756, N9757, N9758, N9759, N9760, N9761, N9762, N9763, N9764, N9765, N9766, N9767, N9768, N9769, N9770, N9771, N9772, N9773, N9774, N9775, N9776, N9777, N9778, N9779, N9780, N9781, N9782, N9783, N9784, N9785, N9786, N9787, N9788, N9789, N9790, N9791, N9792, N9793, N9794, N9795, N9796, N9797, N9798, N9799, N9800, N9801, N9802, N9803, N9804, N9805, N9806, N9807, N9808, N9809, N9810, N9811, N9812, N9813, N9814, N9815, N9816, N9817, N9818, N9819, N9820, N9821, N9822, N9823, N9824, N9825, N9826, N9827, N9828, N9829, N9830, N9831, N9832, N9833, N9834, N9835, N9836, N9837, N9838, N9839, N9840, N9841, N9842, N9843, N9844, N9845, N9846, N9847, N9848, N9849, N9850, N9851, N9852, N9853, N9854, N9855, N9856, N9857, N9858, N9859, N9860, N9861, N9862, N9863, N9864, N9865, N9866, N9867, N9868, N9869, N9870, N9871, N9872, N9873, N9874, N9875, N9876, N9877, N9878, N9879, N9880, N9881, N9882, N9883, N9884, N9885, N9886, N9887, N9888, N9889, N9890, N9891, N9892, N9893, N9894, N9895, N9896, N9897, N9898, N9899, N9900, N9901, N9902, N9903, N9904, N9905, N9906, N9907, N9908, N9909, N9910, N9911, N9912, N9913, N9914, N9915, N9916, N9917, N9918, N9919, N9920, N9921, N9922, N9923, N9924, N9925, N9926, N9927, N9928, N9929, N9930, N9931, N9932, N9933, N9934, N9935, N9936, N9937, N9938, N9939, N9940, N9941, N9942, N9943, N9944, N9945, N9946, N9947, N9948, N9949, N9950, N9951, N9952, N9953, N9954, N9955, N9956, N9957, N9958, N9959, N9960, N9961, N9962, N9963, N9964, N9965, N9966, N9967, N9968, N9969, N9970, N9971, N9972, N9973, N9974, N9975, N9976, N9977, N9978, N9979, N9980, N9981, N9982, N9983, N9984, N9985, N9986, N9987, N9988, N9989, N9990, N9991, N9992, N9993, N9994, N9995, N9996, N9997, N9998, N9999, N10000, N10001, N10002, N10003, N10004, N10005, N10006, N10007, N10008, N10009, N10010, N10011, N10012, N10013, N10014, N10015, N10016, N10017, N10018, N10019, N10020, N10021, N10022, N10023, N10024, N10025, N10026, N10027, N10028, N10029, N10030, N10031, N10032, N10033, N10034, N10035, N10036, N10037, N10038, N10039, N10040, N10041, N10042, N10043, N10044, N10045, N10046, N10047, N10048, N10049, N10050, N10051, N10052, N10053, N10054, N10055, N10056, N10057, N10058, N10059, N10060, N10061, N10062, N10063, N10064, N10065, N10066, N10067, N10068, N10069, N10070, N10071, N10072, N10073, N10074, N10075, N10076, N10077, N10078, N10079, N10080, N10081, N10082, N10083, N10084, N10085, N10086, N10087, N10088, N10089, N10090, N10091, N10092, N10093, N10094, N10095, N10096, N10097, N10098, N10099, N10100, N10101, N10102, N10103, N10104, N10105, N10106, N10107, N10108, N10109, N10110, N10111, N10112, N10113, N10114, N10115, N10116, N10117, N10118, N10119, N10120, N10121, N10122, N10123, N10124, N10125, N10126, N10127, N10128, N10129, N10130, N10131, N10132, N10133, N10134, N10135, N10136, N10137, N10138, N10139, N10140, N10141, N10142, N10143, N10144, N10145, N10146, N10147, N10148, N10149, N10150, N10151, N10152, N10153, N10154, N10155, N10156, N10157, N10158, N10159, N10160, N10161, N10162, N10163, N10164, N10165, N10166, N10167, N10168, N10169, N10170, N10171, N10172, N10173, N10174, N10175, N10176, N10177, N10178, N10179, N10180, N10181, N10182, N10183, N10184, N10185, N10186, N10187, N10188, N10189, N10190, N10191, N10192, N10193, N10194, N10195, N10196, N10197, N10198, N10199, N10200, N10201, N10202, N10203, N10204, N10205, N10206, N10207, N10208, N10209, N10210, N10211, N10212, N10213, N10214, N10215, N10216, N10217, N10218, N10219, N10220, N10221, N10222, N10223, N10224, N10225, N10226, N10227, N10228, N10229, N10230, N10231, N10232, N10233, N10234, N10235, N10236, N10237, N10238, N10239, N10240, N10241, N10242, N10243, N10244, N10245, N10246, N10247, N10248, N10249, N10250, N10251, N10252, N10253, N10254, N10255, N10256, N10257, N10258, N10259, N10260, N10261, N10262, N10263, N10264, N10265, N10266, N10267, N10268, N10269, N10270, N10271, N10272, N10273, N10274, N10275, N10276, N10277, N10278, N10279, N10280, N10281, N10282, N10283, N10284, N10285, N10286, N10287, N10288, N10289, N10290, N10291, N10292, N10293, N10294, N10295, N10296, N10297, N10298, N10299, N10300, N10301, N10302, N10303, N10304, N10305, N10306, N10307, N10308, N10309, N10310, N10311, N10312, N10313, N10314, N10315, N10316, N10317, N10318, N10319, N10320, N10321, N10322, N10323, N10324, N10325, N10326, N10327, N10328, N10329, N10330, N10331, N10332, N10333, N10334, N10335, N10336, N10337, N10338, N10339, N10340, N10341, N10342, N10343, N10344, N10345, N10346, N10347, N10348, N10349, N10350, N10351, N10352, N10353, N10354, N10355, N10356, N10357, N10358, N10359, N10360, N10361, N10362, N10363, N10364, N10365, N10366, N10367, N10368, N10369, N10370, N10371, N10372, N10373, N10374, N10375, N10376, N10377, N10378, N10379, N10380, N10381, N10382, N10383, N10384, N10385, N10386, N10387, N10388, N10389, N10390, N10391, N10392, N10393, N10394, N10395, N10396, N10397, N10398, N10399, N10400, N10401, N10402, N10403, N10404, N10405, N10406, N10407, N10408, N10409, N10410, N10411, N10412, N10413, N10414, N10415, N10416, N10417, N10418, N10419, N10420, N10421, N10422, N10423, N10424, N10425, N10426, N10427, N10428, N10429, N10430, N10431, N10432, N10433, N10434, N10435, N10436, N10437, N10438, N10439, N10440, N10441, N10442, N10443, N10444, N10445, N10446, N10447, N10448, N10449, N10450, N10451, N10452, N10453, N10454, N10455, N10456, N10457, N10458, N10459, N10460, N10461, N10462, N10463, N10464, N10465, N10466, N10467, N10468, N10469, N10470, N10471, N10472, N10473, N10474, N10475, N10476, N10477, N10478, N10479, N10480, N10481, N10482, N10483, N10484, N10485, N10486, N10487, N10488, N10489, N10490, N10491, N10492, N10493, N10494, N10495, N10496, N10497, N10498, N10499, N10500, N10501, N10502, N10503, N10504, N10505, N10506, N10507, N10508, N10509, N10510, N10511, N10512, N10513, N10514, N10515, N10516, N10517, N10518, N10519, N10520, N10521, N10522, N10523, N10524, N10525, N10526, N10527, N10528, N10529, N10530, N10531, N10532, N10533, N10534, N10535, N10536, N10537, N10538, N10539, N10540, N10541, N10542, N10543, N10544, N10545, N10546, N10547, N10548, N10549, N10550, N10551, N10552, N10553, N10554, N10555, N10556, N10557, N10558, N10559, N10560, N10561, N10562, N10563, N10564, N10565, N10566, N10567, N10568, N10569, N10570, N10571, N10572, N10573, N10574, N10575, N10576, N10577, N10578, N10579, N10580, N10581, N10582, N10583, N10584, N10585, N10586, N10587, N10588, N10589, N10590, N10591, N10592, N10593, N10594, N10595, N10596, N10597, N10598, N10599, N10600, N10601, N10602, N10603, N10604, N10605, N10606, N10607, N10608, N10609, N10610, N10611, N10612, N10613, N10614, N10615, N10616, N10617, N10618, N10619, N10620, N10621, N10622, N10623, N10624, N10625, N10626, N10627, N10628, N10629, N10630, N10631, N10632, N10633, N10634, N10635, N10636, N10637, N10638, N10639, N10640, N10641, N10642, N10643, N10644, N10645, N10646, N10647, N10648, N10649, N10650, N10651, N10652, N10653, N10654, N10655, N10656, N10657, N10658, N10659, N10660, N10661, N10662, N10663, N10664, N10665, N10666, N10667, N10668, N10669, N10670, N10671, N10672, N10673, N10674, N10675, N10676, N10677, N10678, N10679, N10680, N10681, N10682, N10683, N10684, N10685, N10686, N10687, N10688, N10689, N10690, N10691, N10692, N10693, N10694, N10695, N10696, N10697, N10698, N10699, N10700, N10701, N10702, N10703, N10704, N10705, N10706, N10707, N10708, N10709, N10710, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10719, N10720, N10721, N10722, N10723, N10724, N10725, N10726, N10727, N10728, N10729, N10730, N10731, N10732, N10733, N10734, N10735, N10736, N10737, N10738, N10739, N10740, N10741, N10742, N10743, N10744, N10745, N10746, N10747, N10748, N10749, N10750, N10751, N10752, N10753, N10754, N10755, N10756, N10757, N10758, N10759, N10760, N10761, N10762, N10763, N10764, N10765, N10766, N10767, N10768, N10769, N10770, N10771, N10772, N10773, N10774, N10775, N10776, N10777, N10778, N10779, N10780, N10781, N10782, N10783, N10784, N10785, N10786, N10787, N10788, N10789, N10790, N10791, N10792, N10793, N10794, N10795, N10796, N10797, N10798, N10799, N10800, N10801, N10802, N10803, N10804, N10805, N10806, N10807, N10808, N10809, N10810, N10811, N10812, N10813, N10814, N10815, N10816, N10817, N10818, N10819, N10820, N10821, N10822, N10823, N10824, N10825, N10826, N10827, N10828, N10829, N10830, N10831, N10832, N10833, N10834, N10835, N10836, N10837, N10838, N10839, N10840, N10841, N10842, N10843, N10844, N10845, N10846, N10847, N10848, N10849, N10850, N10851, N10852, N10853, N10854, N10855, N10856, N10857, N10858, N10859, N10860, N10861, N10862, N10863, N10864, N10865, N10866, N10867, N10868, N10869, N10870, N10871, N10872, N10873, N10874, N10875, N10876, N10877, N10878, N10879, N10880, N10881, N10882, N10883, N10884, N10885, N10886, N10887, N10888, N10889, N10890, N10891, N10892, N10893, N10894, N10895, N10896, N10897, N10898, N10899, N10900, N10901, N10902, N10903, N10904, N10905, N10906, N10907, N10908, N10909, N10910, N10911, N10912, N10913, N10914, N10915, N10916, N10917, N10918, N10919, N10920, N10921, N10922, N10923, N10924, N10925, N10926, N10927, N10928, N10929, N10930, N10931, N10932, N10933, N10934, N10935, N10936, N10937, N10938, N10939, N10940, N10941, N10942, N10943, N10944, N10945, N10946, N10947, N10948, N10949, N10950, N10951, N10952, N10953, N10954, N10955, N10956, N10957, N10958, N10959, N10960, N10961, N10962, N10963, N10964, N10965, N10966, N10967, N10968, N10969, N10970, N10971, N10972, N10973, N10974, N10975, N10976, N10977, N10978, N10979, N10980, N10981, N10982, N10983, N10984, N10985, N10986, N10987, N10988, N10989, N10990, N10991, N10992, N10993, N10994, N10995, N10996, N10997, N10998, N10999, N11000, N11001, N11002, N11003, N11004, N11005, N11006, N11007, N11008, N11009, N11010, N11011, N11012, N11013, N11014, N11015, N11016, N11017, N11018, N11019, N11020, N11021, N11022, N11023, N11024, N11025, N11026, N11027, N11028, N11029, N11030, N11031, N11032, N11033, N11034, N11035, N11036, N11037, N11038, N11039, N11040, N11041, N11042, N11043, N11044, N11045, N11046, N11047, N11048, N11049, N11050, N11051, N11052, N11053, N11054, N11055, N11056, N11057, N11058, N11059, N11060, N11061, N11062, N11063, N11064, N11065, N11066, N11067, N11068, N11069, N11070, N11071, N11072, N11073, N11074, N11075, N11076, N11077, N11078, N11079, N11080, N11081, N11082, N11083, N11084, N11085, N11086, N11087, N11088, N11089, N11090, N11091, N11092, N11093, N11094, N11095, N11096, N11097, N11098, N11099, N11100, N11101, N11102, N11103, N11104, N11105, N11106, N11107, N11108, N11109, N11110, N11111, N11112, N11113, N11114, N11115, N11116, N11117, N11118, N11119, N11120, N11121, N11122, N11123, N11124, N11125, N11126, N11127, N11128, N11129, N11130, N11131, N11132, N11133, N11134, N11135, N11136, N11137, N11138, N11139, N11140, N11141, N11142, N11143, N11144, N11145, N11146, N11147, N11148, N11149, N11150, N11151, N11152, N11153, N11154, N11155, N11156, N11157, N11158, N11159, N11160, N11161, N11162, N11163, N11164, N11165, N11166, N11167, N11168, N11169, N11170, N11171, N11172, N11173, N11174, N11175, N11176, N11177, N11178, N11179, N11180, N11181, N11182, N11183, N11184, N11185, N11186, N11187, N11188, N11189, N11190, N11191, N11192, N11193, N11194, N11195, N11196, N11197, N11198, N11199, N11200, N11201, N11202, N11203, N11204, N11205, N11206, N11207, N11208, N11209, N11210, N11211, N11212, N11213, N11214, N11215, N11216, N11217, N11218, N11219, N11220, N11221, N11222, N11223, N11224, N11225, N11226, N11227, N11228, N11229, N11230, N11231, N11232, N11233, N11234, N11235, N11236, N11237, N11238, N11239, N11240, N11241, N11242, N11243, N11244, N11245, N11246, N11247, N11248, N11249, N11250, N11251, N11252, N11253, N11254, N11255, N11256, N11257, N11258, N11259, N11260, N11261, N11262, N11263, N11264, N11265, N11266, N11267, N11268, N11269, N11270, N11271, N11272, N11273, N11274, N11275, N11276, N11277, N11278, N11279, N11280, N11281, N11282, N11283, N11284, N11285, N11286, N11287, N11288, N11289, N11290, N11291, N11292, N11293, N11294, N11295, N11296, N11297, N11298, N11299, N11300, N11301, N11302, N11303, N11304, N11305, N11306, N11307, N11308, N11309, N11310, N11311, N11312, N11313, N11314, N11315, N11316, N11317, N11318, N11319, N11320, N11321, N11322, N11323, N11324, N11325, N11326, N11327, N11328, N11329, N11330, N11331, N11332, N11333, N11334, N11335, N11336, N11337, N11338, N11339, N11340, N11341, N11342, N11343, N11344, N11345, N11346, N11347, N11348, N11349, N11350, N11351, N11352, N11353, N11354, N11355, N11356, N11357, N11358, N11359, N11360, N11361, N11362, N11363, N11364, N11365, N11366, N11367, N11368, N11369, N11370, N11371, N11372, N11373, N11374, N11375, N11376, N11377, N11378, N11379, N11380, N11381, N11382, N11383, N11384, N11385, N11386, N11387, N11388, N11389, N11390, N11391, N11392, N11393, N11394, N11395, N11396, N11397, N11398, N11399, N11400, N11401, N11402, N11403, N11404, N11405, N11406, N11407, N11408, N11409, N11410, N11411, N11412, N11413, N11414, N11415, N11416, N11417, N11418, N11419, N11420, N11421, N11422, N11423, N11424, N11425, N11426, N11427, N11428, N11429, N11430, N11431, N11432, N11433, N11434, N11435, N11436, N11437, N11438, N11439, N11440, N11441, N11442, N11443, N11444, N11445, N11446, N11447, N11448, N11449, N11450, N11451, N11452, N11453, N11454, N11455, N11456, N11457, N11458, N11459, N11460, N11461, N11462, N11463, N11464, N11465, N11466, N11467, N11468, N11469, N11470, N11471, N11472, N11473, N11474, N11475, N11476, N11477, N11478, N11479, N11480, N11481, N11482, N11483, N11484, N11485, N11486, N11487, N11488, N11489, N11490, N11491, N11492, N11493, N11494, N11495, N11496, N11497, N11498, N11499, N11500, N11501, N11502, N11503, N11504, N11505, N11506, N11507, N11508, N11509, N11510, N11511, N11512, N11513, N11514, N11515, N11516, N11517, N11518, N11519, N11520, N11521, N11522, N11523, N11524, N11525, N11526, N11527, N11528, N11529, N11530, N11531, N11532, N11533, N11534, N11535, N11536, N11537, N11538, N11539, N11540, N11541, N11542, N11543, N11544, N11545, N11546, N11547, N11548, N11549, N11550, N11551, N11552, N11553, N11554, N11555, N11556, N11557, N11558, N11559, N11560, N11561, N11562, N11563, N11564, N11565, N11566, N11567, N11568, N11569, N11570, N11571, N11572, N11573, N11574, N11575, N11576, N11577, N11578, N11579, N11580, N11581, N11582, N11583, N11584, N11585, N11586, N11587, N11588, N11589, N11590, N11591, N11592, N11593, N11594, N11595, N11596, N11597, N11598, N11599, N11600, N11601, N11602, N11603, N11604, N11605, N11606, N11607, N11608, N11609, N11610, N11611, N11612, N11613, N11614, N11615, N11616, N11617, N11618, N11619, N11620, N11621, N11622, N11623, N11624, N11625, N11626, N11627, N11628, N11629, N11630, N11631, N11632, N11633, N11634, N11635, N11636, N11637, N11638, N11639, N11640, N11641, N11642, N11643, N11644, N11645, N11646, N11647, N11648, N11649, N11650, N11651, N11652, N11653, N11654, N11655, N11656, N11657, N11658, N11659, N11660, N11661, N11662, N11663, N11664, N11665, N11666, N11667, N11668, N11669, N11670, N11671, N11672, N11673, N11674, N11675, N11676, N11677, N11678, N11679, N11680, N11681, N11682, N11683, N11684, N11685, N11686, N11687, N11688, N11689, N11690, N11691, N11692, N11693, N11694, N11695, N11696, N11697, N11698, N11699, N11700, N11701, N11702, N11703, N11704, N11705, N11706, N11707, N11708, N11709, N11710, N11711, N11712, N11713, N11714, N11715, N11716, N11717, N11718, N11719, N11720, N11721, N11722, N11723, N11724, N11725, N11726, N11727, N11728, N11729, N11730, N11731, N11732, N11733, N11734, N11735, N11736, N11737, N11738, N11739, N11740, N11741, N11742, N11743, N11744, N11745, N11746, N11747, N11748, N11749, N11750, N11751, N11752, N11753, N11754, N11755, N11756, N11757, N11758, N11759, N11760, N11761, N11762, N11763, N11764, N11765, N11766, N11767, N11768, N11769, N11770, N11771, N11772, N11773, N11774, N11775, N11776, N11777, N11778, N11779, N11780, N11781, N11782, N11783, N11784, N11785, N11786, N11787, N11788, N11789, N11790, N11791, N11792, N11793, N11794, N11795, N11796, N11797, N11798, N11799, N11800, N11801, N11802, N11803, N11804, N11805, N11806, N11807, N11808, N11809, N11810, N11811, N11812, N11813, N11814, N11815, N11816, N11817, N11818, N11819, N11820, N11821, N11822, N11823, N11824, N11825, N11826, N11827, N11828, N11829, N11830, N11831, N11832, N11833, N11834, N11835, N11836, N11837, N11838, N11839, N11840, N11841, N11842, N11843, N11844, N11845, N11846, N11847, N11848, N11849, N11850, N11851, N11852, N11853, N11854, N11855, N11856, N11857, N11858, N11859, N11860, N11861, N11862, N11863, N11864, N11865, N11866, N11867, N11868, N11869, N11870, N11871, N11872, N11873, N11874, N11875, N11876, N11877, N11878, N11879, N11880, N11881, N11882, N11883, N11884, N11885, N11886, N11887, N11888, N11889, N11890, N11891, N11892, N11893, N11894, N11895, N11896, N11897, N11898, N11899, N11900, N11901, N11902, N11903, N11904, N11905, N11906, N11907, N11908, N11909, N11910, N11911, N11912, N11913, N11914, N11915, N11916, N11917, N11918, N11919, N11920, N11921, N11922, N11923, N11924, N11925, N11926, N11927, N11928, N11929, N11930, N11931, N11932, N11933, N11934, N11935, N11936, N11937, N11938, N11939, N11940, N11941, N11942, N11943, N11944, N11945, N11946, N11947, N11948, N11949, N11950, N11951, N11952, N11953, N11954, N11955, N11956, N11957, N11958, N11959, N11960, N11961, N11962, N11963, N11964, N11965, N11966, N11967, N11968, N11969, N11970, N11971, N11972, N11973, N11974, N11975, N11976, N11977, N11978, N11979, N11980, N11981, N11982, N11983, N11984, N11985, N11986, N11987, N11988, N11989, N11990, N11991, N11992, N11993, N11994, N11995, N11996, N11997, N11998, N11999, N12000, N12001, N12002, N12003, N12004, N12005, N12006, N12007, N12008, N12009, N12010, N12011, N12012, N12013, N12014, N12015, N12016, N12017, N12018, N12019, N12020, N12021, N12022, N12023, N12024, N12025, N12026, N12027, N12028, N12029, N12030, N12031, N12032, N12033, N12034, N12035, N12036, N12037, N12038, N12039, N12040, N12041, N12042, N12043, N12044, N12045, N12046, N12047, N12048, N12049, N12050, N12051, N12052, N12053, N12054, N12055, N12056, N12057, N12058, N12059, N12060, N12061, N12062, N12063, N12064, N12065, N12066, N12067, N12068, N12069, N12070, N12071, N12072, N12073, N12074, N12075, N12076, N12077, N12078, N12079, N12080, N12081, N12082, N12083, N12084, N12085, N12086, N12087, N12088, N12089, N12090, N12091, N12092, N12093, N12094, N12095, N12096, N12097, N12098, N12099, N12100, N12101, N12102, N12103, N12104, N12105, N12106, N12107, N12108, N12109, N12110, N12111, N12112, N12113, N12114, N12115, N12116, N12117, N12118, N12119, N12120, N12121, N12122, N12123, N12124, N12125, N12126, N12127, N12128, N12129, N12130, N12131, N12132, N12133, N12134, N12135, N12136, N12137, N12138, N12139, N12140, N12141, N12142, N12143, N12144, N12145, N12146, N12147, N12148, N12149, N12150, N12151, N12152, N12153, N12154, N12155, N12156, N12157, N12158, N12159, N12160, N12161, N12162, N12163, N12164, N12165, N12166, N12167, N12168, N12169, N12170, N12171, N12172, N12173, N12174, N12175, N12176, N12177, N12178, N12179, N12180, N12181, N12182, N12183, N12184, N12185, N12186, N12187, N12188, N12189, N12190, N12191, N12192, N12193, N12194, N12195, N12196, N12197, N12198, N12199, N12200, N12201, N12202, N12203, N12204, N12205, N12206, N12207, N12208, N12209, N12210, N12211, N12212, N12213, N12214, N12215, N12216, N12217, N12218, N12219, N12220, N12221, N12222, N12223, N12224, N12225, N12226, N12227, N12228, N12229, N12230, N12231, N12232, N12233, N12234, N12235, N12236, N12237, N12238, N12239, N12240, N12241, N12242, N12243, N12244, N12245, N12246, N12247, N12248, N12249, N12250, N12251, N12252, N12253, N12254, N12255, N12256, N12257, N12258, N12259, N12260, N12261, N12262, N12263, N12264, N12265, N12266, N12267, N12268, N12269, N12270, N12271, N12272, N12273, N12274, N12275, N12276, N12277, N12278, N12279, N12280, N12281, N12282, N12283, N12284, N12285, N12286, N12287, N12288, N12289, N12290, N12291, N12292, N12293, N12294, N12295, N12296, N12297, N12298, N12299, N12300, N12301, N12302, N12303, N12304, N12305, N12306, N12307, N12308, N12309, N12310, N12311, N12312, N12313, N12314, N12315, N12316, N12317, N12318, N12319, N12320, N12321, N12322, N12323, N12324, N12325, N12326, N12327, N12328, N12329, N12330, N12331, N12332, N12333, N12334, N12335, N12336, N12337, N12338, N12339, N12340, N12341, N12342, N12343, N12344, N12345, N12346, N12347, N12348, N12349, N12350, N12351, N12352, N12353, N12354, N12355, N12356, N12357, N12358, N12359, N12360, N12361, N12362, N12363, N12364, N12365, N12366, N12367, N12368, N12369, N12370, N12371, N12372, N12373, N12374, N12375, N12376, N12377, N12378, N12379, N12380, N12381, N12382, N12383, N12384, N12385, N12386, N12387, N12388, N12389, N12390, N12391, N12392, N12393, N12394, N12395, N12396, N12397, N12398, N12399, N12400, N12401, N12402, N12403, N12404, N12405, N12406, N12407, N12408, N12409, N12410, N12411, N12412, N12413, N12414, N12415, N12416, N12417, N12418, N12419, N12420, N12421, N12422, N12423, N12424, N12425, N12426, N12427, N12428, N12429, N12430, N12431, N12432, N12433, N12434, N12435, N12436, N12437, N12438, N12439, N12440, N12441, N12442, N12443, N12444, N12445, N12446, N12447, N12448, N12449, N12450, N12451, N12452, N12453, N12454, N12455, N12456, N12457, N12458, N12459, N12460, N12461, N12462, N12463, N12464, N12465, N12466, N12467, N12468, N12469, N12470, N12471, N12472, N12473, N12474, N12475, N12476, N12477, N12478, N12479, N12480, N12481, N12482, N12483, N12484, N12485, N12486, N12487, N12488, N12489, N12490, N12491, N12492, N12493, N12494, N12495, N12496, N12497, N12498, N12499, N12500, N12501, N12502, N12503, N12504, N12505, N12506, N12507, N12508, N12509, N12510, N12511, N12512, N12513, N12514, N12515, N12516, N12517, N12518, N12519, N12520, N12521, N12522, N12523, N12524, N12525, N12526, N12527, N12528, N12529, N12530, N12531, N12532, N12533, N12534, N12535, N12536, N12537, N12538, N12539, N12540, N12541, N12542, N12543, N12544, N12545, N12546, N12547, N12548, N12549, N12550, N12551, N12552, N12553, N12554, N12555, N12556, N12557, N12558, N12559, N12560, N12561, N12562, N12563, N12564, N12565, N12566, N12567, N12568, N12569, N12570, N12571, N12572, N12573, N12574, N12575, N12576, N12577, N12578, N12579, N12580, N12581, N12582, N12583, N12584, N12585, N12586, N12587, N12588, N12589, N12590, N12591, N12592, N12593, N12594, N12595, N12596, N12597, N12598, N12599, N12600, N12601, N12602, N12603, N12604, N12605, N12606, N12607, N12608, N12609, N12610, N12611, N12612, N12613, N12614, N12615, N12616, N12617, N12618, N12619, N12620, N12621, N12622, N12623, N12624, N12625, N12626, N12627, N12628, N12629, N12630, N12631, N12632, N12633, N12634, N12635, N12636, N12637, N12638, N12639, N12640, N12641, N12642, N12643, N12644, N12645, N12646, N12647, N12648, N12649, N12650, N12651, N12652, N12653, N12654, N12655, N12656, N12657, N12658, N12659, N12660, N12661, N12662, N12663, N12664, N12665, N12666, N12667, N12668, N12669, N12670, N12671, N12672, N12673, N12674, N12675, N12676, N12677, N12678, N12679, N12680, N12681, N12682, N12683, N12684, N12685, N12686, N12687, N12688, N12689, N12690, N12691, N12692, N12693, N12694, N12695, N12696, N12697, N12698, N12699, N12700, N12701, N12702, N12703, N12704, N12705, N12706, N12707, N12708, N12709, N12710, N12711, N12712, N12713, N12714, N12715, N12716, N12717, N12718, N12719, N12720, N12721, N12722, N12723, N12724, N12725, N12726, N12727, N12728, N12729, N12730, N12731, N12732, N12733, N12734, N12735, N12736, N12737, N12738, N12739, N12740, N12741, N12742, N12743, N12744, N12745, N12746, N12747, N12748, N12749, N12750, N12751, N12752, N12753, N12754, N12755, N12756, N12757, N12758, N12759, N12760, N12761, N12762, N12763, N12764, N12765, N12766, N12767, N12768, N12769, N12770, N12771, N12772, N12773, N12774, N12775, N12776, N12777, N12778, N12779, N12780, N12781, N12782, N12783, N12784, N12785, N12786, N12787, N12788, N12789, N12790, N12791, N12792, N12793, N12794, N12795, N12796, N12797, N12798, N12799, N12800, N12801, N12802, N12803, N12804, N12805, N12806, N12807, N12808, N12809, N12810, N12811, N12812, N12813, N12814, N12815, N12816, N12817, N12818, N12819, N12820, N12821, N12822, N12823, N12824, N12825, N12826, N12827, N12828, N12829, N12830, N12831, N12832, N12833, N12834, N12835, N12836, N12837, N12838, N12839, N12840, N12841, N12842, N12843, N12844, N12845, N12846, N12847, N12848, N12849, N12850, N12851, N12852, N12853, N12854, N12855, N12856, N12857, N12858, N12859, N12860, N12861, N12862, N12863, N12864, N12865, N12866, N12867, N12868, N12869, N12870, N12871, N12872;
    output N12874, N12877, N12881, N12891, N12892, N12897, N12899, N12905, N12908, N12911, N12916, N12918, N12920, N12924, N12925, N12931, N12933, N12943, N12949, N12952, N12958, N12965, N12969, N12973, N12980, N12981, N12991, N12995, N12996, N13008, N13015, N13021, N13023, N13024, N13028, N13033, N13035, N13040, N13043, N13065, N13071, N13084, N13096, N13110, N13118, N13120, N13123, N13124, N13132, N13144, N13154, N13157, N13165, N13168, N13170, N13182, N13189, N13200, N13206, N13211, N13217, N13225, N13228, N13233, N13241, N13242, N13250, N13257, N13276, N13277, N13283, N13307, N13309, N13310, N13326, N13327, N13330, N13339, N13342, N13348, N13353, N13360, N13361, N13362, N13369, N13373, N13376, N13377, N13381, N13396, N13408, N13410, N13415, N13420, N13421, N13431, N13434, N13442, N13443, N13444, N13446, N13448, N13456, N13457, N13458, N13465, N13466, N13482, N13483, N13490, N13492, N13505, N13512, N13514, N13517, N13524, N13527, N13533, N13536, N13547, N13548, N13551, N13556, N13563, N13566, N13577, N13589, N13594, N13595, N13608, N13610, N13611, N13612, N13615, N13616, N13628, N13633, N13647, N13650, N13651, N13663, N13666, N13673, N13674, N13679, N13681, N13684, N13686, N13691, N13699, N13700, N13707, N13711, N13718, N13719, N13734, N13737, N13741, N13742, N13761, N13767, N13770, N13775, N13776, N13781, N13785, N13789, N13803, N13806, N13809, N13811, N13819, N13820, N13828, N13838, N13842, N13844, N13847, N13852, N13858, N13867, N13869, N13870, N13873, N13880, N13885, N13893, N13896, N13901, N13905, N13906, N13910, N13915, N13920, N13921, N13929, N13932, N13934, N13941, N13956, N13959, N13965, N13969, N13972, N13991, N14000, N14005, N14018, N14019, N14033, N14034, N14037, N14040, N14045, N14052, N14056, N14060, N14079, N14084, N14087, N14100, N14101, N14104, N14107, N14113, N14119, N14124, N14125, N14126, N14147, N14151, N14158, N14159, N14161, N14165, N14171, N14174, N14180, N14185, N14186, N14187, N14203, N14205, N14207, N14208, N14212, N14214, N14215, N14216, N14217, N14219, N14222, N14234, N14243, N14269, N14274, N14275, N14280, N14288, N14289, N14291, N14296, N14298, N14311, N14318, N14321, N14337, N14347, N14352, N14354, N14355, N14359, N14361, N14368, N14382, N14385, N14416, N14417, N14424, N14428, N14429, N14433, N14436, N14441, N14443, N14444, N14453, N14455, N14462, N14469, N14471, N14480, N14481, N14490, N14499, N14502, N14507, N14515, N14518, N14519, N14528, N14546, N14553, N14563, N14568, N14570, N14577, N14578, N14594, N14600, N14603, N14604, N14606, N14608, N14613, N14623, N14637, N14638, N14653, N14663, N14666, N14671, N14679, N14680, N14685, N14691, N14694, N14698, N14709, N14715, N14725, N14733, N14736, N14744, N14752, N14755, N14756, N14767, N14775, N14783, N14785, N14791, N14812, N14824, N14826, N14831, N14837, N14839, N14840, N14848, N14849, N14850, N14863, N14867, N14876, N14881, N14890, N14898, N14899, N14920, N14922, N14931, N14936, N14939, N14947, N14953, N14958, N14961, N14968, N14969, N14971, N14978, N14991, N14992, N15002, N15005, N15006, N15013, N15015, N15018, N15032, N15035, N15038, N15071, N15075, N15078, N15085, N15090, N15100, N15101, N15104, N15105, N15107, N15110, N15111, N15114, N15126, N15134, N15144, N15148, N15152, N15156, N15158, N15169, N15170, N15171, N15173, N15174, N15183, N15185, N15199, N15201, N15209, N15214, N15217, N15224, N15228, N15233, N15249, N15254, N15255, N15257, N15259, N15260, N15274, N15278, N15291, N15294, N15296, N15303, N15304, N15307, N15308, N15310, N15313, N15317, N15319, N15323, N15331, N15346, N15353, N15354, N15362, N15366, N15379, N15390, N15402, N15403, N15410, N15422, N15434, N15442, N15444, N15453, N15455, N15469, N15473, N15485, N15489, N15494, N15496, N15497, N15500, N15501, N15504, N15513, N15516, N15519, N15520, N15522, N15529, N15532, N15534, N15537, N15540, N15541, N15543, N15545, N15550, N15556, N15561, N15564, N15572, N15575, N15591, N15592, N15600, N15622, N15638, N15643, N15646, N15653, N15660, N15664, N15670, N15673, N15677, N15678, N15680, N15691, N15693, N15705, N15708, N15709, N15711, N15715, N15719, N15722, N15724, N15738, N15740, N15741, N15748, N15756, N15761, N15766, N15774, N15788, N15793, N15795, N15798, N15799, N15818, N15819, N15823, N15828, N15831, N15835, N15836, N15837, N15844, N15847, N15852, N15854, N15878, N15889, N15890, N15893, N15908, N15910, N15916, N15929, N15934, N15948, N15951, N15963, N15969, N15970, N15975, N15984, N15991, N16008, N16009, N16010, N16012, N16014, N16020, N16022, N16026, N16029, N16035, N16036, N16042, N16046, N16050, N16057, N16058, N16060, N16068, N16079, N16081, N16095, N16110, N16111, N16112, N16113, N16116, N16118, N16121, N16123, N16133, N16138, N16142, N16154, N16160, N16170, N16177, N16183, N16191, N16193, N16197, N16198, N16201, N16202, N16210, N16215, N16231, N16233, N16255, N16256, N16266, N16274, N16278, N16282, N16283, N16289, N16290, N16301, N16303, N16323, N16326, N16328, N16330, N16332, N16334, N16341, N16353, N16364, N16367, N16379, N16385, N16394, N16398, N16400, N16402, N16403, N16409, N16416, N16417, N16421, N16428, N16442, N16450, N16453, N16457, N16458, N16462, N16466, N16474, N16480, N16487, N16494, N16499, N16516, N16519, N16527, N16529, N16533, N16537, N16551, N16556, N16560, N16565, N16571, N16576, N16578, N16582, N16586, N16591, N16592, N16598, N16601, N16602, N16616, N16629, N16631, N16632, N16634, N16642, N16645, N16649, N16666, N16667, N16674, N16677, N16682, N16684, N16687, N16695, N16709, N16717, N16725, N16730, N16738, N16742, N16747, N16760, N16765, N16782, N16796, N16797, N16801, N16803, N16806, N16809, N16814, N16818, N16828, N16830, N16839, N16841, N16846, N16847, N16848, N16854, N16867, N16871, N16879, N16883, N16891, N16906, N16911, N16920, N16925, N16939, N16940, N16942, N16949, N16954, N16956, N16971, N16981, N16984, N16990, N16996, N16999, N17002, N17004, N17017, N17018, N17019, N17024, N17041, N17043, N17052, N17053, N17063, N17066, N17076, N17082, N17083, N17091, N17095, N17098, N17102, N17106, N17107, N17110, N17115, N17124, N17127, N17141, N17148, N17156, N17169, N17181, N17182, N17183, N17188, N17191, N17193, N17203, N17209, N17210, N17214, N17216, N17219, N17221, N17223, N17236, N17243, N17250, N17251, N17252, N17255, N17260, N17264, N17274, N17278, N17285, N17291, N17301, N17304, N17310, N17318, N17323, N17335, N17337, N17342, N17360, N17362, N17367, N17369, N17375, N17384, N17393, N17397, N17399, N17400, N17413, N17425, N17428, N17431, N17444, N17445, N17446, N17451, N17459, N17460, N17464, N17480, N17482, N17494, N17495, N17512, N17521, N17523, N17526, N17529, N17536, N17537, N17542, N17544, N17548, N17550, N17555, N17571, N17578, N17579, N17582, N17586, N17590, N17591, N17593, N17601, N17604, N17609, N17612, N17614, N17619, N17633, N17642, N17649, N17650, N17662, N17665, N17673, N17674, N17675, N17685, N17686, N17701, N17707, N17709, N17711, N17719, N17723, N17727, N17728, N17735, N17745, N17749, N17753, N17766, N17770, N17794, N17800, N17804, N17806, N17832, N17838, N17843, N17847, N17852, N17858, N17885, N17888, N17894, N17895, N17897, N17903, N17905, N17908, N17911, N17912, N17917, N17918, N17922, N17925, N17927, N17931, N17934, N17935, N17943, N17944, N17945, N17948, N17966, N17971, N17972, N17983, N17993, N17997, N17999, N18005, N18007, N18010, N18016, N18022, N18027, N18029, N18042, N18054, N18058, N18060, N18081, N18097, N18101, N18109, N18110, N18112, N18120, N18126, N18138, N18144, N18149, N18153, N18157, N18159, N18166, N18172, N18173, N18174, N18189, N18201, N18203, N18219, N18234, N18240, N18245, N18249, N18261, N18264, N18267, N18271, N18279, N18281, N18285, N18303, N18310, N18322, N18338, N18339, N18350, N18351, N18354, N18362, N18364, N18372, N18375, N18379, N18400, N18416, N18420, N18430, N18436, N18445, N18461, N18464, N18467, N18484, N18488, N18493, N18495, N18502, N18506, N18510, N18519, N18524, N18526, N18528, N18544, N18549, N18561, N18563, N18566, N18576, N18578, N18583, N18587, N18619, N18622, N18627, N18641, N18649, N18665, N18668, N18671, N18685, N18688, N18693, N18723, N18724, N18730, N18737, N18739, N18741, N18743, N18751, N18754, N18776, N18781, N18783, N18799, N18805, N18820, N18822, N18825, N18834, N18838, N18848, N18850, N18855, N18866, N18867, N18881, N18883, N18884, N18887, N18899, N18907, N18912, N18919, N18921, N18924, N18929, N18937, N18939, N18944, N18949, N18955, N18971, N18980, N18981, N18983, N18984, N18988, N18991, N18999, N19007, N19008, N19011, N19017, N19033, N19038, N19048, N19051, N19056, N19057, N19058, N19063, N19066, N19068, N19070, N19076, N19087, N19088, N19095, N19097, N19100, N19104, N19105, N19108, N19109, N19112, N19113, N19116, N19129, N19130, N19139, N19160, N19174, N19175, N19178, N19182, N19187, N19190, N19194, N19207, N19209, N19212, N19213, N19215, N19220, N19224, N19241, N19242, N19246, N19247, N19248, N19251, N19265, N19274, N19277, N19279, N19296, N19303, N19306, N19314, N19324, N19326, N19329, N19334, N19340, N19341, N19346, N19347, N19350, N19375, N19380, N19386, N19388, N19399, N19402, N19409, N19430, N19445, N19447, N19457, N19459, N19474, N19481, N19482, N19484, N19493, N19499, N19524, N19527, N19531, N19532, N19534, N19536, N19537, N19543, N19549, N19561, N19564, N19567, N19568, N19570, N19577, N19583, N19585, N19593, N19596, N19617, N19622, N19623, N19630, N19633, N19657, N19658, N19668, N19670, N19673, N19676, N19678, N19686, N19693, N19696, N19714, N19729, N19743, N19744, N19746, N19747, N19748, N19751, N19763, N19780, N19785, N19816, N19819, N19822, N19823, N19824, N19829, N19832, N19839, N19844, N19851, N19852, N19859, N19864, N19870, N19871, N19872, N19881, N19892, N19893, N19897, N19905, N19909, N19918, N19920, N19921, N19927, N19937, N19938, N19939, N19942, N19948, N19951, N19953, N19960, N19968, N19969, N19978, N19986, N19988, N19995, N19998, N20002, N20003, N20007, N20010, N20018, N20019, N20036, N20042, N20047, N20048, N20055, N20057, N20059, N20060, N20066, N20068, N20069, N20072, N20074, N20077, N20082, N20087, N20089, N20099, N20105, N20108, N20119, N20123, N20125, N20135, N20138, N20146, N20154, N20158, N20164, N20186, N20189, N20190, N20191, N20192, N20197, N20199, N20203, N20208, N20217, N20218, N20227, N20249, N20270, N20277, N20278, N20279, N20281, N20284, N20286, N20287, N20291, N20292, N20295, N20299, N20300, N20309, N20314, N20333, N20345, N20354, N20359, N20360, N20367, N20369, N20376, N20394, N20396, N20403, N20404, N20407, N20408, N20409, N20411, N20413, N20422, N20425, N20429, N20445, N20455, N20458, N20479, N20484, N20493, N20495, N20507, N20508, N20515, N20522, N20523, N20533, N20534, N20536, N20541, N20545, N20547, N20567, N20576, N20577, N20586, N20588, N20594, N20598, N20601, N20602, N20604, N20606, N20607, N20610, N20613, N20618, N20619, N20629, N20637, N20638, N20640, N20650, N20652, N20653, N20661, N20663, N20668, N20680, N20685, N20692, N20703, N20710, N20727, N20744, N20747, N20748, N20771, N20773, N20776, N20783, N20787, N20791, N20799, N20803, N20806, N20807, N20808, N20816, N20818, N20823, N20824, N20843, N20851, N20863, N20864, N20870, N20873, N20874, N20888, N20893, N20900, N20902, N20906, N20911, N20916, N20921, N20924, N20933, N20935, N20938, N20941, N20952, N20958, N20963, N20970, N20971, N21001, N21019, N21022, N21023, N21024, N21036, N21037, N21038, N21041, N21050, N21051, N21064, N21065, N21074, N21085, N21086, N21094, N21095, N21096, N21106, N21115, N21116, N21119, N21122, N21134, N21140, N21145, N21150, N21157, N21161, N21170, N21191, N21192, N21203, N21206, N21211, N21213, N21214, N21217, N21219, N21226, N21227, N21228, N21231, N21235, N21238, N21241, N21248, N21251, N21252, N21254, N21257, N21261, N21264, N21270, N21274, N21276, N21284, N21285, N21287, N21291, N21292, N21296, N21302, N21304, N21306, N21307, N21316, N21323, N21325, N21327, N21330, N21331, N21332, N21333, N21334, N21336, N21349, N21350, N21352, N21354, N21356, N21357, N21362, N21368, N21371, N21372, N21377, N21382, N21386, N21388, N21395, N21397, N21399, N21402, N21404, N21406, N21416, N21421, N21426, N21432, N21433, N21438, N21445, N21450, N21452, N21457, N21459, N21465, N21466, N21467, N21468, N21469, N21470, N21481, N21483, N21485, N21491, N21498, N21503, N21509, N21516, N21518, N21521, N21523, N21527, N21530, N21537, N21538, N21540, N21546, N21547, N21555, N21561, N21562, N21566, N21567, N21569, N21571, N21582, N21584, N21585, N21586, N21590, N21591, N21597, N21598, N21607, N21609, N21610, N21611, N21613, N21617, N21622, N21624, N21629, N21631, N21636, N21637, N21641, N21654, N21669, N21672, N21675, N21684, N21685, N21686, N21687, N21688, N21692, N21694, N21698, N21705, N21712, N21715, N21717, N21719, N21721, N21727, N21739, N21741, N21742, N21745, N21746, N21753, N21758, N21769, N21770, N21772, N21773, N21781, N21786, N21788, N21795, N21796, N21797, N21798, N21813, N21833, N21835, N21842, N21852, N21857, N21860, N21862, N21864, N21868, N21869, N21871, N21876, N21882, N21885, N21889, N21891, N21898, N21902, N21908, N21909, N21914, N21916, N21918, N21930, N21935, N21943, N21954, N21957, N21958, N21959, N21964, N21966, N21971, N21978, N21982, N21983, N21987, N21989, N21991, N21994, N21995, N21996, N21998, N21999, N22003, N22008, N22014, N22018, N22019, N22023, N22024, N22026, N22029, N22032, N22037, N22040, N22043, N22049, N22052, N22053, N22058, N22059, N22060, N22064, N22066, N22067, N22068, N22069, N22070, N22071, N22073, N22076, N22077, N22080, N22081, N22084, N22100, N22102, N22104, N22105, N22116, N22117, N22121, N22123, N22126, N22132, N22140, N22142, N22145, N22147, N22150, N22157, N22161, N22167, N22173, N22177, N22183, N22185, N22186, N22188, N22191, N22197, N22199, N22204, N22206, N22213, N22215, N22217, N22218, N22221, N22222, N22223, N22225, N22234, N22235, N22237, N22240, N22241, N22243, N22244, N22248, N22249, N22251, N22257, N22262, N22263, N22266, N22272, N22284, N22287, N22302, N22303, N22307, N22311, N22312, N22315, N22317, N22324, N22327, N22329, N22330, N22332, N22334, N22340, N22341, N22342, N22343, N22344, N22350, N22354, N22363, N22365, N22368, N22372, N22377, N22380, N22382, N22391, N22397, N22398, N22400, N22401, N22420, N22424, N22430, N22432, N22435, N22439, N22440, N22446, N22454, N22460, N22467, N22470, N22472, N22473, N22488, N22489, N22490, N22495, N22498, N22503, N22510, N22511, N22512, N22516, N22517, N22520, N22521, N22523, N22528, N22537, N22541, N22547, N22549, N22551, N22552, N22560, N22561, N22563, N22568, N22578, N22589, N22595, N22597, N22606, N22618, N22621, N22622, N22629, N22631, N22634, N22638, N22648, N22650, N22656, N22659, N22664, N22676, N22677, N22682, N22683, N22684, N22693, N22694, N22699, N22704, N22705, N22706, N22709, N22714, N22715, N22724, N22727, N22730, N22737, N22749, N22761, N22764, N22769, N22779, N22780, N22782, N22783, N22790, N22792, N22794, N22797, N22804, N22806, N22809, N22810, N22818, N22819, N22821, N22822, N22823, N22824, N22827, N22829, N22831, N22834, N22840, N22842, N22846, N22850, N22860, N22861, N22873, N22876, N22880, N22884, N22888, N22893, N22895, N22900, N22901, N22902, N22911, N22914, N22916, N22918, N22920, N22922, N22934, N22941, N22942, N22947, N22951, N22955, N22959, N22968, N22978, N22980, N22984, N22991, N22994, N22997, N22998, N23000, N23001, N23007, N23008, N23009, N23018, N23019, N23026, N23028, N23029, N23032, N23038, N23054, N23056, N23057, N23058, N23059, N23064, N23068, N23072, N23076, N23081, N23086, N23087, N23090, N23092, N23093, N23101, N23102, N23110, N23111, N23112, N23114, N23116, N23117, N23121, N23126, N23129, N23133, N23135, N23137, N23141, N23142, N23147, N23148, N23157, N23159, N23165, N23170, N23178, N23186, N23188, N23194, N23196, N23197, N23198, N23199, N23201, N23214, N23217, N23218, N23221, N23222, N23223, N23224, N23225, N23228, N23231, N23232, N23241, N23244, N23245, N23246, N23247, N23251, N23259, N23261, N23262, N23269, N23277, N23280, N23283, N23287, N23289, N23297, N23300, N23312, N23315, N23316, N23320, N23324, N23331, N23336, N23349, N23351, N23359, N23365, N23366, N23367, N23369, N23370, N23374, N23376, N23378, N23390, N23391, N23392, N23395, N23397, N23406, N23413, N23415, N23420, N23433, N23439, N23447, N23455, N23456, N23457, N23458, N23459, N23468, N23475, N23478, N23481, N23482, N23486, N23489, N23492, N23493, N23494, N23506, N23508, N23515, N23517, N23521, N23522, N23528, N23535, N23537, N23540, N23547, N23554, N23558, N23559, N23560, N23563, N23567, N23575, N23579, N23587, N23588, N23590, N23592, N23594, N23597, N23600, N23602, N23607, N23610, N23611, N23613, N23622, N23630, N23634, N23636, N23641, N23646, N23655, N23656, N23660, N23661, N23667, N23671, N23675, N23680, N23685, N23693, N23699, N23700, N23701, N23702, N23705, N23708, N23712, N23732, N23738, N23739, N23746, N23749, N23755, N23758, N23759, N23760, N23769, N23770, N23771, N23772, N23774, N23778, N23783, N23791, N23795, N23800, N23803, N23805, N23815, N23817, N23819, N23824, N23830, N23831, N23832, N23843, N23844, N23845, N23846, N23847, N23848, N23852, N23853, N23858, N23861, N23869, N23870, N23872, N23874, N23878, N23889, N23891, N23894, N23896, N23897, N23905, N23908, N23922, N23925, N23926, N23942, N23944, N23947, N23951, N23954, N23963, N23967, N23975, N23978, N23981, N23983, N23988, N23991, N23994, N24010, N24023, N24024, N24027, N24028, N24033, N24041, N24043, N24047, N24052, N24053, N24061, N24062, N24065, N24066, N24068, N24069, N24079, N24080, N24081, N24084, N24092, N24097, N24098, N24104, N24115, N24117, N24130, N24131, N24133, N24134, N24137, N24138, N24139, N24140, N24143, N24144, N24151, N24153, N24161, N24162, N24164, N24168, N24172, N24173, N24178, N24188, N24192, N24196, N24214, N24221, N24222, N24230, N24234, N24238, N24241, N24244, N24246, N24249, N24254, N24259, N24266, N24273, N24274, N24277, N24279, N24283, N24286, N24290, N24295, N24297, N24298, N24299, N24302, N24305, N24309, N24312, N24314, N24315, N24325, N24327, N24342, N24347, N24352, N24360, N24362, N24372, N24374, N24380, N24381, N24393, N24399, N24403, N24404, N24407, N24420, N24426, N24436, N24440, N24443, N24445, N24446, N24454, N24457, N24466, N24468, N24472, N24483, N24486, N24489, N24493, N24506, N24512, N24515, N24516, N24519, N24527, N24530, N24531, N24534, N24535, N24539, N24544, N24552, N24555, N24557, N24574, N24578, N24582, N24584, N24590, N24592, N24593, N24598, N24599, N24603, N24607, N24609, N24613, N24615, N24619, N24621, N24622, N24624, N24628, N24633, N24638, N24642, N24644, N24646, N24647, N24650, N24651, N24657, N24663, N24675, N24696, N24706, N24711, N24715, N24717, N24724, N24732, N24736, N24739, N24742, N24747, N24749, N24752, N24757, N24761, N24775, N24776, N24777, N24782, N24783, N24784, N24785, N24807, N24813, N24814, N24815, N24823, N24824, N24826, N24829, N24830, N24832, N24840, N24844, N24847, N24848, N24855, N24856, N24858, N24859, N24864, N24869, N24870, N24871, N24872, N24877, N24884, N24885, N24887, N24890, N24894, N24895, N24896, N24903, N24917, N24922, N24927, N24929, N24933, N24937, N24938, N24939, N24941, N24943, N24945, N24946, N24950, N24954, N24956, N24964, N24968, N24969, N24973, N24975, N24978, N24979, N24983, N24990, N24992, N25003, N25006, N25012, N25016, N25017, N25021, N25033, N25042, N25045, N25054, N25057, N25062, N25064, N25066, N25067, N25069, N25079, N25080, N25088, N25091, N25092, N25113, N25114, N25115, N25118, N25120, N25121, N25122, N25123, N25132, N25135, N25136, N25143, N25144, N25157, N25158, N25165, N25170, N25171, N25172, N25179, N25181, N25186, N25190, N25192, N25193, N25199, N25200, N25207, N25210, N25229, N25233, N25235, N25237, N25238, N25239, N25240, N25247, N25256, N25257, N25260, N25265, N25266, N25267, N25268, N25272, N25278, N25281, N25282, N25285, N25288, N25295, N25296, N25309, N25310, N25313, N25316, N25318, N25319, N25324, N25330, N25337, N25339, N25340, N25345, N25347, N25350, N25356, N25358, N25359, N25368, N25373, N25375, N25376, N25380, N25381, N25390, N25396, N25397, N25399, N25400, N25401, N25407, N25412, N25420, N25425, N25426, N25429, N25430, N25431, N25434, N25437, N25439, N25443, N25448, N25451, N25452, N25456, N25458, N25461, N25464, N25468, N25470, N25472, N25473, N25480, N25483, N25489, N25491, N25500, N25501, N25505, N25506, N25512, N25514, N25520, N25521, N25523, N25527, N25530, N25535, N25538, N25540, N25541, N25542, N25543, N25545, N25549, N25552, N25554, N25556, N25558, N25559, N25560, N25575, N25576, N25577, N25578, N25585, N25587, N25589, N25595, N25596, N25599, N25606, N25609, N25610, N25611, N25612, N25616, N25617, N25618, N25620, N25622, N25623, N25628, N25629, N25634, N25637, N25643, N25645, N25646, N25647, N25648, N25652, N25655, N25659, N25666, N25667, N25670, N25673, N25674, N25675, N25678, N25682, N25684, N25686, N25687, N25688, N25690, N25695, N25705, N25709, N25711, N25713, N25714, N25715, N25722, N25724, N25726, N25727, N25729, N25733, N25735, N25736, N25737, N25739, N25740, N25742, N25744, N25746, N25749, N25752, N25755, N25757, N25761, N25762, N25763, N25767, N25769, N25770, N25772, N25779, N25780, N25781, N25791, N25793, N25797, N25798, N25807, N25809, N25811, N25812, N25818, N25828, N25835, N25838, N25840, N25843, N25848, N25851, N25853, N25854, N25855, N25859, N25861, N25867, N25870, N25888, N25892, N25896, N25907, N25908, N25910, N25913, N25914, N25918, N25923, N25928, N25935, N25936, N25944, N25946, N25948, N25958, N25959, N25960, N25968, N25970, N25971, N25972, N25976, N25978, N25988, N26000, N26002, N26005, N26006, N26009, N26010, N26020, N26023, N26024, N26028, N26029, N26032, N26034, N26039, N26042, N26048, N26050, N26052, N26053, N26055, N26056, N26058, N26062, N26065, N26072, N26073, N26076, N26077, N26078, N26079, N26080, N26091, N26094, N26096, N26097, N26100, N26103, N26104, N26106, N26112, N26113, N26116, N26118, N26120, N26123, N26124, N26131, N26132, N26134, N26137, N26138, N26139, N26141, N26146, N26152, N26153, N26154, N26161, N26162, N26163, N26166, N26170, N26171, N26181, N26183, N26188, N26189, N26191, N26192, N26197, N26199, N26200, N26201, N26204, N26206, N26208, N26214, N26215, N26219, N26221, N26223, N26227, N26228, N26230, N26231, N26234, N26235, N26236, N26237, N26238, N26244, N26246, N26247, N26249, N26251, N26254, N26259, N26261, N26264, N26273, N26274, N26276, N26277, N26279, N26284, N26285, N26286, N26288, N26289, N26298, N26304, N26317, N26322, N26326, N26329, N26337, N26339, N26346, N26347, N26349, N26351, N26353, N26354, N26358, N26359, N26361, N26363, N26365, N26367, N26369, N26372, N26374, N26375, N26378, N26384, N26385, N26386, N26387, N26397, N26399, N26400, N26402, N26403, N26406, N26408, N26409, N26410, N26413, N26429, N26432, N26434, N26435, N26436, N26440, N26442, N26446, N26452, N26453, N26454, N26461, N26467, N26470, N26475, N26477, N26478, N26480, N26483, N26490, N26492, N26494, N26496, N26499, N26500, N26503, N26505, N26514, N26515, N26518, N26521, N26522, N26523, N26524, N26528, N26529, N26531, N26534, N26535, N26537, N26540, N26541, N26551, N26553, N26558, N26562, N26563, N26570, N26571, N26573, N26574, N26575, N26577, N26592, N26593, N26594, N26603, N26609, N26611, N26620, N26625, N26629, N26630, N26631, N26637, N26640, N26644, N26649, N26656, N26659, N26660, N26662, N26668, N26672, N26681, N26692, N26698, N26699, N26701, N26702, N26705, N26706, N26710, N26712, N26714, N26717, N26718, N26721, N26726, N26728, N26736, N26739, N26741, N26743, N26745, N26747, N26757, N26760, N26765, N26766, N26771, N26776, N26777, N26781, N26784, N26785, N26787, N26789, N26790, N26794, N26798, N26799, N26800, N26803, N26809, N26816, N26820, N26821, N26822, N26823, N26825, N26828, N26830, N26832, N26837, N26844, N26845, N26851, N26854, N26855, N26857, N26864, N26865, N26880, N26885, N26886, N26895, N26896, N26899, N26903, N26904, N26905, N26907, N26909, N26912, N26913, N26921, N26923, N26924, N26930, N26931, N26939, N26940, N26942, N26945, N26950, N26954, N26955, N26957, N26961, N26964, N26971, N26973, N26984, N26986, N26987, N26988, N26989, N26991, N26992, N26993, N26997, N26999, N27001, N27002, N27004, N27010, N27013, N27014, N27016, N27021, N27023, N27024, N27025, N27027, N27034, N27035, N27036, N27038, N27040, N27041, N27042, N27045, N27046, N27047, N27048, N27058, N27061, N27063, N27065, N27071, N27073, N27074, N27075, N27078, N27079, N27088, N27090, N27091, N27094, N27106, N27114, N27118, N27120, N27128, N27129, N27130, N27133, N27134, N27135, N27136, N27142, N27148, N27150, N27158, N27159, N27166, N27169, N27172, N27180, N27187, N27188, N27189, N27192, N27193, N27194, N27195, N27198, N27200, N27202, N27203, N27204, N27208, N27212, N27216, N27222, N27224, N27227, N27228, N27230, N27233, N27238, N27242, N27243, N27244, N27246, N27248, N27251, N27253, N27254, N27258, N27263, N27273, N27277, N27284, N27292, N27295, N27299, N27302, N27306, N27307, N27311, N27312, N27313, N27315, N27322, N27323, N27326, N27330, N27333, N27335, N27338, N27341, N27343, N27344, N27345, N27348, N27350, N27351, N27352, N27356, N27359, N27363, N27364, N27367, N27371, N27372, N27375, N27381, N27383, N27385, N27386, N27388, N27390, N27395, N27398, N27400, N27409, N27410, N27414, N27415, N27418, N27424, N27430, N27432, N27435, N27437, N27441, N27443, N27446, N27447, N27450, N27451, N27457, N27458, N27460, N27461, N27466, N27468, N27469, N27470, N27471, N27475, N27476, N27481, N27485, N27487, N27490, N27491, N27493, N27494, N27495, N27497, N27502, N27504, N27505, N27529, N27530, N27531, N27539, N27542, N27548, N27550, N27551, N27555, N27559, N27563, N27568, N27569, N27570, N27576, N27579, N27580, N27586, N27587, N27590, N27591, N27603, N27611, N27612, N27613, N27614, N27618, N27622, N27626, N27627, N27628, N27629, N27630, N27632, N27633, N27635, N27636, N27646, N27647, N27648, N27649, N27650, N27653, N27654, N27655, N27660, N27662, N27664, N27665, N27671, N27672, N27675, N27676, N27681, N27682, N27685, N27686, N27689, N27693, N27699, N27701, N27704, N27708, N27711, N27713, N27716, N27719, N27720, N27721, N27722, N27728, N27729, N27731, N27733, N27735, N27738, N27744, N27748, N27751, N27752, N27756, N27757, N27762, N27764, N27769, N27770, N27775, N27778, N27780, N27783, N27786, N27787, N27788, N27789, N27790, N27792, N27794, N27798, N27804, N27805, N27807, N27809, N27811, N27813, N27818, N27828, N27829, N27830, N27833, N27835, N27837, N27841, N27842, N27844, N27848, N27849, N27850, N27854, N27856, N27861, N27868, N27873, N27879, N27883, N27886, N27887, N27890, N27894, N27896, N27900, N27903, N27906, N27907, N27915, N27918, N27922, N27931, N27932, N27935, N27941, N27942, N27944, N27947, N27949, N27954, N27955, N27958, N27959, N27965, N27967, N27974, N27976, N27977, N27984, N27986, N27988, N27990, N27994, N28000, N28001, N28003, N28005, N28007, N28012, N28026, N28030, N28032, N28033, N28035, N28038, N28039, N28040, N28048, N28051, N28054, N28059, N28062, N28065, N28067, N28068, N28071, N28073, N28074, N28075, N28080, N28084, N28085, N28099, N28100, N28108, N28117, N28119, N28120, N28123, N28128, N28129, N28130, N28131, N28134, N28140, N28145, N28149, N28152, N28153, N28155, N28157, N28166, N28167, N28168, N28173, N28175, N28180, N28181, N28184, N28187, N28188, N28189, N28196, N28200, N28207, N28209, N28210, N28212, N28213, N28216, N28221, N28223, N28224, N28225, N28228, N28230, N28231, N28236, N28239, N28240, N28243, N28247, N28249, N28251, N28255, N28259, N28261, N28262, N28263, N28266, N28268, N28274, N28275, N28278, N28280, N28281, N28283, N28285, N28286, N28288, N28291, N28292, N28293, N28296, N28300, N28306, N28315, N28316, N28319, N28322, N28323, N28327, N28330, N28331, N28332, N28333, N28337, N28338, N28340, N28341, N28343, N28351, N28355, N28357, N28360, N28362, N28366, N28367, N28369, N28370, N28373, N28376, N28377, N28378, N28383, N28388, N28391, N28394, N28395, N28398, N28400, N28402, N28407, N28413, N28414, N28415, N28416, N28420, N28424, N28425, N28428, N28433, N28438, N28442, N28447, N28449, N28453, N28454, N28462, N28464, N28468, N28470, N28473, N28474, N28480, N28482, N28484, N28489, N28492, N28502, N28504, N28505, N28509, N28517, N28518, N28519, N28524, N28525, N28527, N28530, N28533, N28534, N28535, N28536, N28539, N28541, N28542, N28543, N28549, N28550, N28552, N28558, N28562, N28563, N28573, N28576, N28579, N28580, N28583, N28584, N28591, N28592, N28593, N28595, N28597, N28598, N28604, N28605, N28607, N28608, N28609, N28612, N28613, N28621, N28623, N28624, N28626, N28632, N28638, N28641, N28647, N28648, N28658, N28661, N28666, N28670, N28671, N28672, N28676, N28683, N28694, N28696, N28700, N28707, N28713, N28715, N28722, N28723, N28725, N28728, N28733, N28734, N28735, N28736, N28745, N28748, N28751, N28752, N28755, N28759, N28765, N28775, N28778, N28780, N28784, N28790, N28791, N28792, N28799, N28800, N28802, N28806, N28811, N28812, N28814, N28816, N28818, N28824, N28826, N28827, N28829, N28830, N28834, N28835, N28849, N28851, N28852, N28853, N28858, N28862, N28863, N28866, N28869, N28872, N28875, N28879, N28881, N28883, N28887, N28890, N28898, N28899, N28900, N28902, N28903, N28917, N28918, N28924, N28926, N28928, N28929, N28931, N28932, N28934, N28935, N28936, N28940, N28941, N28947, N28955, N28961, N28967, N28971, N28972, N28976, N28985, N28992, N28994, N29001, N29002, N29003, N29017, N29020, N29023, N29029, N29034, N29042, N29045, N29053, N29054, N29056, N29057, N29059, N29060, N29062, N29067, N29068, N29070, N29073, N29074, N29076, N29077, N29080, N29081, N29086, N29092, N29095, N29096, N29103, N29111, N29112, N29115, N29121, N29123, N29124, N29126, N29127, N29128, N29137, N29138, N29140, N29141, N29142, N29143, N29145, N29152, N29155, N29161, N29166, N29171, N29177, N29178, N29184, N29187, N29189, N29192, N29194, N29199, N29200, N29202, N29203, N29204, N29206, N29209, N29213, N29215, N29218, N29220, N29224, N29229, N29234, N29237, N29252, N29256, N29258, N29261, N29267, N29268, N29269, N29273, N29277, N29283, N29288, N29290, N29291, N29297, N29301, N29302, N29303, N29306, N29307, N29312, N29328, N29334, N29336, N29338, N29341, N29342, N29345, N29348, N29349, N29350, N29356, N29357, N29360, N29361, N29362, N29368, N29369, N29370, N29373, N29378, N29379, N29380, N29381, N29387, N29390, N29395, N29396, N29404, N29411, N29414, N29415, N29417, N29421, N29426, N29427, N29429, N29439, N29447, N29448, N29452, N29461, N29462, N29466, N29469, N29471, N29473, N29476, N29478, N29482, N29488, N29493, N29497, N29498, N29499, N29501, N29507, N29520, N29527, N29529, N29530, N29533, N29534, N29537, N29538, N29539, N29543, N29549, N29550, N29552, N29554, N29558, N29562, N29563, N29568, N29570, N29571, N29572, N29573, N29576, N29579, N29581, N29584, N29585, N29588, N29590, N29594, N29601, N29605, N29606, N29610, N29614, N29620, N29624, N29627, N29628, N29631, N29632, N29633, N29640, N29641, N29643, N29645, N29646, N29648, N29649, N29651, N29652, N29654, N29655, N29657, N29658, N29659, N29662, N29663, N29666, N29668, N29669, N29670, N29676, N29679, N29682, N29686, N29690, N29691, N29693, N29699, N29700, N29703, N29711, N29712, N29713, N29724, N29726, N29727, N29729, N29731, N29734, N29742, N29746, N29747, N29748, N29750, N29751, N29760, N29764, N29765, N29767, N29768, N29779, N29785, N29786, N29787, N29789, N29794, N29795, N29796, N29798, N29802, N29804, N29808, N29811, N29812, N29813, N29816, N29817, N29820, N29822, N29825, N29829, N29833, N29836, N29837, N29840, N29843, N29845, N29846, N29849, N29850, N29852, N29853, N29855, N29857, N29863, N29866, N29873, N29874, N29875, N29876, N29878, N29879, N29885, N29886, N29894, N29899, N29901, N29907, N29913, N29918, N29923, N29925, N29926, N29927, N29928, N29931, N29934, N29935, N29942, N29944, N29946, N29947, N29948, N29952, N29953, N29955, N29956, N29957, N29959, N29960, N29965, N29966, N29969, N29972, N29975, N29976, N29980, N29981, N29984, N29987, N29988, N30007, N30008, N30009, N30012, N30015, N30027, N30031, N30034, N30035, N30036, N30042, N30044, N30045, N30046, N30050, N30057, N30059, N30060, N30064, N30066, N30070, N30077, N30079, N30080, N30084, N30085, N30091, N30093, N30096, N30097, N30098, N30102, N30104, N30105, N30108, N30109, N30110, N30111, N30116, N30118, N30119, N30123, N30124, N30127, N30135, N30137, N30138, N30139, N30140, N30141, N30142, N30143, N30144, N30146, N30148, N30149, N30150, N30155, N30157, N30158, N30161, N30162, N30163, N30164, N30165, N30169, N30170, N30171, N30174, N30176, N30177, N30178, N30179, N30180, N30181, N30183, N30184, N30186, N30187, N30188, N30189, N30190, N30191, N30192, N30193, N30194, N30195, N30196, N30197, N30198, N30199, N30201, N30203, N30205, N30206, N30208, N30210, N30212, N30213, N30214, N30215, N30216, N30217, N30218, N30219, N30221, N30222, N30223, N30224, N30225, N30226, N30227, N30228, N30230, N30233, N30236, N30237, N30239, N30241, N30242, N30243, N30245, N30247, N30248, N30249, N30252, N30253, N30255, N30256, N30258, N30259, N30260, N30262, N30263, N30264, N30265, N30266, N30267, N30268, N30270, N30272, N30273, N30275, N30278, N30279, N30280, N30281, N30283, N30284, N30286, N30288, N30292, N30293, N30295, N30296, N30297, N30298, N30301, N30303, N30305, N30307, N30309, N30313, N30314, N30316, N30317, N30319, N30321, N30322, N30323, N30325, N30326, N30330, N30331, N30333, N30334, N30336, N30337, N30338, N30339, N30341, N30343, N30344, N30345, N30347, N30348, N30350, N30352, N30354, N30357, N30358, N30359, N30361, N30363, N30364, N30365, N30366, N30367, N30369, N30370, N30372, N30373, N30374, N30375, N30376, N30377, N30378, N30381, N30382, N30383, N30386, N30389, N30391, N30393, N30395, N30396, N30398, N30401, N30404, N30405, N30406, N30407, N30411, N30412, N30413, N30414, N30415, N30416, N30418, N30419, N30420, N30421, N30424, N30426, N30427, N30428, N30432, N30434, N30435, N30437, N30438, N30440, N30442, N30443, N30444, N30446, N30447, N30448, N30449, N30452, N30453, N30454, N30455, N30456, N30457, N30458, N30459, N30460, N30461, N30462, N30463, N30466, N30467, N30468, N30469, N30470, N30471, N30474, N30476, N30477, N30479, N30480, N30481, N30484, N30485, N30487, N30488, N30491, N30493, N30495, N30496, N30497, N30498, N30499, N30500, N30502, N30503, N30504, N30505, N30506, N30507, N30508, N30509, N30510, N30514, N30515, N30517, N30519, N30520, N30521, N30522, N30523, N30524, N30527, N30528, N30529, N30530, N30531, N30532, N30533, N30534, N30536, N30537, N30539, N30540, N30544, N30545, N30546, N30551, N30553, N30554, N30557, N30559, N30560, N30561, N30564, N30572, N30575, N30577, N30578, N30579, N30580, N30582, N30584, N30585, N30586, N30588, N30589, N30590, N30591, N30592, N30593, N30595, N30596, N30597, N30598, N30601, N30602, N30603, N30605, N30608, N30609, N30611, N30612, N30613, N30615, N30616, N30617, N30618, N30620, N30621, N30622, N30623, N30625, N30627, N30628, N30631, N30633, N30634, N30635, N30636, N30638, N30639, N30641, N30642, N30643, N30644, N30649, N30650, N30651, N30652, N30654, N30655, N30656, N30658, N30659, N30660, N30662, N30663, N30664, N30665, N30666, N30667, N30668, N30669, N30670, N30671, N30672, N30673, N30674, N30675, N30676, N30677, N30678, N30679, N30681, N30682, N30683, N30685, N30687, N30688, N30689, N30691, N30692, N30693, N30694, N30696, N30699, N30703, N30704, N30705, N30706, N30710, N30712, N30713, N30714, N30716, N30717, N30718, N30719, N30721, N30724, N30725, N30726, N30727, N30730, N30731, N30732, N30735, N30737, N30739, N30741, N30742, N30743, N30744, N30747, N30749, N30750, N30751, N30753, N30755, N30756, N30758, N30759, N30761, N30763, N30766, N30767, N30768, N30769, N30772, N30773, N30774, N30777, N30779, N30780, N30781, N30782, N30784, N30785, N30786, N30787, N30789, N30790, N30791, N30792, N30793, N30794, N30795, N30796, N30801, N30803, N30804, N30806, N30808, N30809, N30810, N30813, N30815, N30816, N30817, N30818, N30819, N30822, N30823, N30824, N30826, N30827, N30828, N30829, N30832, N30833, N30834, N30836, N30837, N30838, N30839, N30840, N30842, N30843, N30845, N30846, N30847, N30849, N30850, N30851, N30852, N30853, N30855, N30856, N30858, N30861, N30862, N30863, N30864, N30865, N30866, N30869, N30871, N30872, N30873, N30875, N30876, N30877, N30879, N30880, N30881, N30882, N30883, N30885, N30886, N30887, N30888, N30890, N30893, N30895, N30896, N30898, N30900, N30901, N30902, N30903, N30904, N30905, N30907, N30908, N30912, N30913, N30914, N30915, N30916, N30917, N30918, N30919, N30921, N30922, N30923, N30925, N30926, N30930, N30933, N30934, N30935, N30936, N30937, N30939, N30942, N30944, N30945, N30946, N30947, N30948, N30949, N30950, N30952, N30953, N30957, N30959, N30960, N30962, N30963, N30964, N30965, N30966, N30968, N30970, N30971, N30972, N30974, N30975, N30976, N30977, N30979, N30981, N30982, N30983, N30986, N30987, N30988, N30991, N30992, N30993, N30994, N30998, N30999, N31000, N31003, N31004, N31005, N31006, N31007, N31009, N31010, N31016, N31017, N31018, N31019, N31020, N31021, N31022, N31023, N31028, N31029, N31032, N31033, N31035, N31036, N31037, N31038, N31039, N31041, N31043, N31045, N31047, N31048, N31050, N31051, N31052, N31053, N31054, N31056, N31057, N31058, N31059, N31061, N31062, N31064, N31065, N31068, N31069, N31071, N31072, N31077, N31078, N31080, N31081, N31082, N31083, N31085, N31088, N31089, N31093, N31094, N31096, N31097, N31098, N31101, N31103, N31105, N31107, N31108, N31110, N31111, N31112, N31113, N31115, N31116, N31117, N31118, N31123, N31125, N31127, N31128, N31129, N31131, N31133, N31134, N31137, N31138, N31141, N31145, N31148, N31149, N31152, N31153, N31155, N31157, N31158, N31159, N31160, N31163, N31164, N31165, N31166, N31167, N31169, N31171, N31172, N31174, N31176, N31178, N31180, N31182, N31184, N31185, N31186, N31188, N31189, N31192, N31193, N31194, N31196, N31197, N31199, N31200, N31202, N31203, N31204, N31205, N31206, N31207, N31210, N31211, N31212, N31213, N31218, N31219, N31220, N31221, N31223, N31224, N31225, N31227, N31229, N31230, N31231, N31232, N31233, N31235, N31236, N31240, N31241, N31243, N31246, N31248, N31251, N31252, N31253, N31255, N31258, N31259, N31260, N31262, N31263, N31266, N31269, N31270, N31271, N31272, N31273, N31274, N31275, N31277, N31280, N31282, N31283, N31284, N31285, N31286, N31287, N31290, N31291, N31293, N31294, N31295, N31297, N31299, N31301, N31308, N31309, N31310, N31312, N31313, N31315, N31317, N31319, N31320, N31321, N31324, N31325, N31326, N31328, N31329, N31332, N31333, N31335, N31336, N31337, N31338, N31339, N31340, N31341, N31342, N31343, N31346, N31350, N31352, N31355, N31356, N31357, N31361, N31362, N31364, N31365, N31367, N31368, N31370, N31371, N31372, N31374, N31375, N31376, N31377, N31378, N31379, N31382, N31383, N31385, N31386, N31387, N31388, N31389, N31390, N31391, N31392, N31393, N31395, N31396, N31397, N31398, N31401, N31402, N31403, N31404, N31405, N31406, N31407, N31408, N31409, N31412, N31414, N31415, N31416, N31417, N31418, N31420, N31421, N31422, N31424, N31425, N31428, N31430, N31431, N31432, N31433, N31434, N31438, N31439, N31441, N31443, N31447, N31448, N31450, N31451, N31452, N31453, N31459, N31463, N31464, N31465, N31466, N31467, N31469, N31471, N31472, N31473, N31474, N31475, N31477, N31478, N31479, N31481, N31482, N31483, N31484, N31485, N31488, N31489, N31490, N31491, N31492, N31495, N31496, N31497, N31498, N31499, N31501, N31502, N31505, N31506, N31507, N31508, N31511, N31512, N31513, N31514, N31516, N31517, N31518, N31519, N31520, N31521, N31522, N31524, N31525, N31527, N31528, N31529, N31532, N31533, N31535, N31536, N31537, N31538, N31540, N31541, N31542, N31543, N31544, N31546, N31548, N31550, N31551, N31553, N31554, N31556, N31557, N31560, N31561, N31562, N31563, N31565, N31566, N31567, N31568, N31570, N31571, N31573, N31574, N31575, N31576, N31579, N31580, N31581, N31582, N31583, N31584, N31586, N31587, N31588, N31589, N31591, N31593, N31594, N31595, N31596, N31597, N31598, N31600, N31603, N31605, N31606, N31608, N31610, N31614, N31615, N31617, N31618, N31619, N31620, N31621, N31622, N31624, N31627, N31628, N31629, N31630, N31632, N31637, N31638, N31642, N31643, N31645, N31647, N31648, N31649, N31651, N31652, N31653, N31654, N31655, N31656, N31657, N31658, N31659, N31660, N31664, N31665, N31666, N31667, N31668, N31670, N31672, N31673, N31674, N31677, N31679, N31681, N31682, N31684, N31685, N31686, N31687, N31688, N31689, N31691, N31692, N31693, N31694, N31695, N31696, N31697, N31698, N31699, N31700, N31701, N31703, N31704, N31705, N31706, N31707, N31708, N31710, N31711, N31712, N31714, N31715, N31717, N31718, N31719, N31720, N31724, N31725, N31728, N31731, N31734, N31736, N31737, N31738, N31740, N31742, N31744, N31745, N31746, N31749, N31752, N31753, N31754, N31757, N31759, N31760, N31761, N31762, N31763, N31764, N31765, N31766, N31767, N31768, N31771, N31772, N31773, N31775, N31776, N31777, N31778, N31781, N31783, N31785, N31787, N31788, N31789, N31790, N31791, N31793, N31794, N31797, N31801, N31802, N31803, N31805, N31806, N31807, N31808, N31810, N31811, N31812, N31813, N31814, N31815, N31817, N31818, N31819, N31820, N31821, N31822, N31823, N31824, N31825, N31826, N31827, N31828, N31829, N31830, N31831, N31833, N31834, N31836, N31837, N31840, N31841, N31842, N31843, N31845, N31846, N31848, N31849, N31850, N31851, N31852, N31854, N31855, N31857, N31858, N31859, N31860, N31865, N31867, N31868, N31870, N31871, N31872, N31873, N31875, N31876, N31880, N31881, N31882, N31883, N31884, N31885, N31887, N31888, N31890, N31891, N31892, N31895, N31896, N31899, N31900, N31903, N31904, N31906, N31907, N31908, N31910, N31911, N31912, N31913, N31915, N31916, N31918, N31920, N31922, N31924, N31925, N31928, N31929, N31930, N31932, N31933, N31937, N31939, N31940, N31941, N31942, N31944, N31945, N31946, N31947, N31948, N31949, N31950, N31953, N31954, N31956, N31957, N31959, N31960, N31962, N31963, N31964, N31965, N31966, N31967, N31969, N31971, N31973, N31974, N31976, N31977, N31979, N31981, N31982, N31983, N31984, N31985, N31988, N31989, N31990, N31991, N31992, N31994, N31996, N31998, N31999, N32000, N32001, N32002, N32004, N32007, N32010, N32012, N32013, N32014, N32015, N32017, N32018, N32019, N32020, N32021, N32026, N32027, N32028, N32030, N32032, N32034, N32036, N32037, N32038, N32040, N32041, N32042, N32045, N32047, N32048, N32050, N32051, N32053, N32054, N32055, N32056, N32057, N32058, N32059, N32062, N32064, N32065, N32066, N32068, N32069, N32070, N32073, N32075, N32076, N32077, N32078, N32079, N32080, N32081, N32082, N32083, N32084, N32087, N32088, N32089, N32090, N32092, N32093, N32097, N32098, N32099, N32101, N32104, N32105, N32106, N32108, N32109, N32110, N32111, N32114, N32117, N32118, N32119, N32121, N32124, N32127, N32129, N32130, N32134, N32135, N32136, N32137, N32138, N32141, N32143, N32144, N32145, N32146, N32147, N32148, N32150, N32151, N32152, N32153, N32154, N32155, N32160, N32161, N32162, N32164, N32165, N32167, N32171, N32173, N32174, N32175, N32176, N32177, N32179, N32182, N32183, N32184, N32186, N32187, N32189, N32190, N32192, N32193, N32195, N32199, N32200, N32201, N32203, N32209, N32210, N32212, N32214, N32216, N32218, N32219, N32222, N32223, N32224, N32225, N32226, N32228, N32229, N32230, N32232, N32233, N32234, N32235, N32236, N32237, N32238, N32240, N32243, N32244, N32246, N32247, N32249, N32250, N32251, N32252, N32253, N32255, N32257, N32259, N32260, N32262, N32263, N32264, N32265, N32266, N32267, N32269, N32272, N32273, N32274, N32275, N32276, N32277, N32278, N32279, N32280, N32282, N32283, N32287, N32288, N32290, N32291, N32292, N32293, N32294, N32295, N32296, N32298, N32301, N32302, N32303, N32304, N32305, N32308, N32309, N32310, N32311, N32312, N32313, N32314, N32315, N32316, N32317, N32318, N32319, N32320, N32321, N32325, N32327, N32328, N32329, N32330, N32333, N32336, N32337, N32339, N32340, N32341, N32342, N32343, N32345, N32346, N32347, N32348, N32349, N32350, N32351, N32352, N32353, N32354, N32355, N32356, N32357, N32359, N32361, N32362, N32363, N32365, N32367, N32369, N32370, N32372, N32373, N32374, N32377, N32378, N32379, N32380, N32382, N32383, N32384, N32385, N32386, N32387, N32388, N32389, N32392, N32393, N32394, N32396, N32397, N32399, N32400, N32401, N32404, N32405, N32406, N32407, N32408, N32409, N32410, N32411, N32412, N32416, N32418, N32419, N32420, N32421, N32422, N32424, N32425, N32426, N32427, N32428, N32429, N32430, N32431, N32432, N32433, N32434, N32435, N32437, N32438, N32439, N32440, N32441, N32442, N32444, N32445, N32446, N32447, N32448, N32449, N32451, N32454, N32455, N32456, N32459, N32460, N32461, N32464, N32465, N32466, N32469, N32471, N32472, N32473, N32474, N32475, N32476, N32480, N32481, N32482, N32483, N32489, N32490, N32491, N32492, N32494, N32496, N32498, N32500, N32501, N32502, N32505, N32506, N32507, N32508, N32511, N32513, N32514, N32517, N32519, N32521, N32522, N32525, N32526, N32527, N32528, N32531, N32532, N32535, N32539, N32540, N32542, N32543, N32544, N32547, N32548, N32550, N32552, N32553, N32554, N32557, N32558, N32559, N32560, N32562, N32563, N32564, N32565, N32567, N32568, N32570, N32573, N32575, N32576, N32577, N32579, N32581, N32582, N32583, N32584, N32585, N32586, N32587, N32589, N32590, N32592, N32593, N32595, N32597, N32598, N32599, N32600, N32602, N32603, N32604, N32606, N32607, N32608, N32610, N32613, N32615, N32616, N32617, N32618, N32619, N32621, N32622, N32623, N32624, N32625, N32626, N32628, N32629, N32631, N32633, N32634, N32635, N32637, N32638, N32639, N32640, N32641, N32642, N32643, N32644, N32645, N32650, N32652, N32653, N32654, N32655, N32656, N32657, N32658, N32661, N32662, N32663, N32665, N32666, N32667, N32668, N32669, N32670, N32671, N32673, N32674, N32676, N32677, N32678, N32679, N32682, N32685, N32686, N32689, N32690, N32691, N32693, N32694, N32695, N32696, N32698, N32700, N32702, N32703, N32704, N32705, N32706, N32707, N32709, N32710, N32712, N32713, N32714, N32716, N32718, N32719, N32720, N32722, N32723, N32725, N32726, N32728, N32730, N32731, N32732, N32733, N32735, N32736, N32737, N32738, N32740, N32741, N32742, N32743, N32744, N32745, N32747, N32748, N32749, N32750, N32752, N32754, N32755, N32756, N32758, N32759, N32760, N32762, N32763, N32764, N32765, N32769, N32770, N32771, N32772, N32773, N32774, N32777, N32778, N32779, N32781, N32782, N32784, N32785, N32786, N32787, N32788, N32789, N32790, N32792, N32793, N32794, N32795, N32796, N32797, N32798, N32799, N32800, N32801, N32802, N32804, N32807, N32809, N32810, N32811, N32812, N32813, N32814, N32817, N32818, N32819, N32820, N32821, N32822, N32823, N32824, N32825, N32828, N32829, N32830, N32832, N32833, N32834, N32837, N32838, N32841, N32842, N32846, N32848, N32849, N32850, N32851, N32852, N32853, N32854, N32858, N32859, N32860, N32862, N32863, N32866, N32867, N32868, N32869, N32871, N32872, N32873, N32874, N32875, N32876, N32877, N32878, N32879, N32880, N32881, N32882, N32883, N32884, N32885, N32886, N32887, N32888, N32890, N32892, N32893, N32896, N32899, N32900, N32901, N32905, N32906, N32907, N32908, N32909, N32911, N32912, N32916, N32917, N32918, N32920, N32923, N32924, N32926, N32930, N32931, N32935, N32936, N32937, N32939, N32940, N32942, N32943, N32944, N32946, N32947, N32948, N32949, N32950, N32952, N32953, N32956, N32957, N32958, N32960, N32965, N32966, N32968, N32969, N32970, N32971, N32972, N32973, N32977, N32978, N32979, N32980, N32982, N32983, N32985, N32986, N32987, N32988, N32990, N32991, N32993, N32994, N32995, N32998, N32999, N33000, N33001, N33002, N33005, N33006, N33007, N33009, N33010, N33012, N33013, N33016, N33018, N33020, N33021, N33022, N33024, N33025, N33026, N33027, N33028, N33029, N33031, N33032, N33034, N33035, N33036, N33037, N33038, N33040, N33044, N33045, N33046, N33047, N33049, N33054, N33055, N33056, N33057, N33058, N33061, N33063, N33064, N33068, N33072, N33073, N33075, N33077, N33078, N33079, N33082, N33083, N33084, N33085, N33087, N33088, N33091, N33092, N33093, N33096, N33098, N33099, N33101, N33105, N33107, N33108, N33109, N33110, N33111, N33112, N33113, N33114, N33115, N33116, N33117, N33119, N33120, N33122, N33124, N33125, N33126, N33127, N33129, N33131, N33132, N33133, N33136, N33138, N33141, N33142, N33143, N33144, N33145, N33146, N33149, N33150, N33151, N33152, N33156, N33157, N33158, N33159, N33160, N33162, N33163, N33164, N33165, N33167, N33168, N33170, N33171, N33173, N33174, N33175, N33177, N33178, N33179, N33180, N33181, N33182, N33183, N33185, N33186, N33188, N33189, N33190, N33191, N33192, N33193, N33194, N33195, N33196, N33197, N33198, N33202, N33203, N33206, N33208, N33209, N33211, N33215, N33216, N33217, N33220, N33221, N33223, N33224, N33226, N33227, N33229, N33231, N33232, N33233, N33234, N33236, N33238, N33240, N33241, N33242, N33244, N33245, N33247, N33248, N33249, N33250, N33253, N33254, N33256, N33257, N33259, N33262, N33263, N33264, N33265, N33266, N33267, N33269, N33274, N33277, N33279, N33282, N33284, N33285, N33287, N33288, N33289, N33291, N33292, N33293, N33294, N33295, N33297, N33299, N33300, N33301, N33302, N33304, N33305, N33306, N33307, N33309, N33310, N33311, N33313, N33315, N33316, N33317, N33318, N33319, N33320, N33321, N33324, N33325, N33327, N33329, N33330, N33331, N33332, N33335, N33336, N33337, N33338, N33339, N33340, N33341, N33342, N33343, N33344, N33345, N33346, N33347, N33348, N33349, N33351, N33352, N33353, N33354, N33355, N33356, N33358, N33359, N33360, N33361, N33362, N33363, N33364, N33365, N33366, N33367, N33368, N33369, N33372, N33373, N33374, N33377, N33378, N33379, N33380, N33384, N33385, N33386, N33387, N33388, N33392, N33396, N33398, N33400, N33401, N33404, N33405, N33406, N33407, N33408, N33410, N33411, N33413, N33414, N33415, N33416, N33418, N33419, N33422, N33423, N33424, N33427, N33431, N33432, N33433, N33434, N33436, N33437, N33441, N33442, N33443, N33446, N33447, N33448, N33450, N33451, N33452, N33453, N33455, N33457, N33458, N33462, N33463, N33464, N33466, N33467, N33468, N33469, N33474, N33476, N33477, N33479, N33481, N33485, N33486, N33487, N33489, N33490, N33491, N33492, N33493, N33496, N33497, N33500, N33501, N33502, N33503, N33504, N33506, N33508, N33509, N33510, N33511, N33513, N33514, N33515, N33516, N33517, N33518, N33519, N33521, N33522, N33524, N33526, N33527, N33528, N33529, N33530, N33531, N33532, N33534, N33536, N33537, N33538, N33539, N33540, N33543, N33546, N33547, N33548, N33550, N33551, N33552, N33553, N33554, N33555, N33556, N33557, N33559, N33560, N33561, N33562, N33563, N33564, N33565, N33568, N33570, N33573, N33574, N33576, N33577, N33578, N33579, N33583, N33584, N33586, N33587, N33588, N33590, N33593, N33594, N33599, N33606, N33609, N33610, N33611, N33613, N33614, N33616, N33618, N33619, N33620, N33621, N33622, N33623, N33625, N33626, N33627, N33628, N33629, N33630, N33631, N33635, N33637, N33639, N33640, N33641, N33642, N33643, N33646, N33647, N33650, N33651, N33652, N33653, N33654, N33655, N33656, N33657, N33658, N33659, N33660, N33661, N33663, N33670, N33672, N33673, N33674, N33675, N33677, N33678, N33679, N33680, N33681, N33683, N33684, N33685, N33687, N33689, N33691, N33692, N33693, N33694, N33695, N33697, N33700, N33701, N33703, N33705, N33706, N33707, N33708, N33709, N33710, N33711, N33712, N33713, N33714, N33718, N33720, N33721, N33722, N33723, N33724, N33725, N33726, N33727, N33729, N33730, N33731, N33733, N33734, N33735, N33738, N33740, N33741, N33742, N33743, N33745, N33746, N33747, N33749, N33750, N33751, N33752, N33753, N33754, N33755, N33757, N33758, N33759, N33761, N33763, N33764, N33765, N33766, N33767, N33769, N33772, N33773, N33774, N33775, N33776, N33777, N33778, N33779, N33780, N33782, N33783, N33784, N33785, N33786, N33787, N33788, N33789, N33792, N33793, N33794, N33795, N33796, N33797, N33798, N33799, N33800, N33801, N33802, N33803, N33804, N33805, N33807, N33809, N33811, N33812, N33813, N33814, N33815, N33818, N33820, N33821, N33822, N33824, N33825, N33826, N33827, N33828, N33829, N33830, N33832, N33833, N33835, N33836, N33837, N33839, N33841, N33842, N33844, N33846, N33848, N33849, N33850, N33851, N33852, N33853, N33854, N33856, N33858, N33859, N33861, N33862, N33863, N33864, N33866, N33867, N33869, N33870, N33871, N33872, N33873, N33875, N33876, N33877, N33878, N33879, N33880, N33881, N33882, N33884, N33888, N33889, N33890, N33891, N33892, N33896, N33897, N33898, N33899, N33900, N33901, N33903, N33904, N33905, N33906, N33907, N33908, N33909, N33911, N33914, N33915, N33916, N33917, N33919, N33921, N33922, N33925, N33927, N33928, N33929, N33930, N33933, N33934, N33935, N33936, N33937, N33940, N33943, N33944, N33945, N33946, N33947, N33948, N33949, N33950, N33951, N33952, N33953, N33955, N33956, N33960, N33961, N33963, N33965, N33966, N33967, N33968, N33969, N33970, N33971, N33972, N33973, N33974, N33975, N33976, N33977, N33978, N33979, N33980, N33983, N33984, N33985, N33986, N33987, N33990, N33992, N33993, N33994, N33995, N33996, N33997, N33998, N34000, N34001, N34002, N34003, N34004, N34005, N34006, N34008, N34009, N34010, N34011, N34016, N34019, N34020, N34021, N34023, N34024, N34025, N34026, N34028, N34031, N34032, N34033, N34035, N34036, N34037, N34039, N34040, N34042, N34043, N34044, N34045, N34046, N34047, N34049, N34050, N34052, N34053, N34054, N34055, N34057, N34058, N34059, N34060, N34061, N34062, N34063, N34065, N34066, N34067, N34068, N34070, N34072, N34073, N34074, N34076, N34077, N34081, N34082, N34084, N34085, N34088, N34090, N34092, N34093, N34095, N34096, N34097, N34098, N34100, N34102, N34103, N34105, N34106, N34107, N34108, N34109, N34110, N34112, N34114, N34115, N34116, N34117, N34118, N34119, N34120, N34121, N34122, N34123, N34124, N34125, N34127, N34128, N34129, N34130, N34131, N34132, N34133, N34135, N34136, N34137, N34141, N34142, N34143, N34145, N34146, N34147, N34148, N34149, N34150, N34151, N34153, N34155, N34156, N34158, N34160, N34161, N34163, N34165, N34166, N34170, N34171, N34174, N34177, N34178, N34179, N34180, N34181, N34183, N34184, N34185, N34186, N34187, N34188, N34189, N34193, N34195, N34196, N34197, N34198, N34199, N34201, N34202, N34205, N34206, N34209, N34210, N34212, N34214, N34217, N34218, N34221, N34223, N34225, N34228, N34229, N34231, N34232, N34233, N34235, N34236, N34237, N34239, N34240, N34242, N34243, N34244, N34245, N34246, N34247, N34248, N34250, N34251, N34252, N34253, N34257, N34259, N34260, N34261, N34263, N34265, N34266, N34267, N34270, N34271, N34274, N34276, N34277, N34278, N34279, N34281, N34282, N34284, N34285, N34287, N34289, N34290, N34292, N34293, N34294, N34295, N34296, N34298, N34299, N34300, N34301, N34302, N34303, N34305, N34306, N34307, N34309, N34310, N34312, N34313, N34314, N34316, N34318, N34319, N34321, N34322, N34323, N34324, N34325, N34330, N34331, N34334, N34336, N34337, N34338, N34341, N34343, N34344, N34345, N34346, N34347, N34350, N34351, N34352, N34355, N34356, N34358, N34359, N34361, N34363, N34364, N34365, N34369, N34371, N34372, N34373, N34374, N34375, N34376, N34378, N34379, N34380, N34384, N34386, N34388, N34389, N34390, N34392, N34393, N34396, N34397, N34399, N34400, N34401, N34403, N34405, N34406, N34409, N34410, N34411, N34412, N34413, N34414, N34416, N34417, N34418, N34419, N34420, N34421, N34422, N34424, N34425, N34426, N34427, N34430, N34432, N34433, N34435, N34436, N34437, N34439, N34440, N34442, N34445, N34446, N34447, N34448, N34449, N34450, N34451, N34454, N34455, N34456, N34457, N34458, N34459, N34460, N34461, N34462, N34463, N34466, N34467, N34468, N34469, N34470, N34471, N34473, N34478, N34480, N34481, N34484, N34487, N34488, N34490, N34493, N34494, N34495, N34496, N34497, N34498, N34499, N34500, N34501, N34502, N34503, N34505, N34508, N34512, N34514, N34517, N34519, N34521, N34522, N34523, N34525, N34526, N34527, N34528, N34531, N34532, N34533, N34534, N34535, N34536, N34537, N34539, N34540, N34541, N34542, N34544, N34545, N34546, N34547, N34548, N34549, N34552, N34554, N34555, N34556, N34557, N34558, N34560, N34561, N34563, N34564, N34565, N34566, N34567, N34568, N34569, N34570, N34571, N34572, N34574, N34576, N34577, N34578, N34579, N34580, N34581, N34583, N34585, N34586, N34587, N34589, N34590, N34591, N34593, N34594, N34595, N34596, N34597, N34598, N34599, N34600, N34602, N34604, N34605, N34606, N34608, N34612, N34613, N34614, N34616, N34618, N34619, N34622, N34623, N34624, N34625, N34626, N34627, N34628, N34629, N34630, N34631, N34633, N34636, N34637, N34638, N34640, N34641, N34642, N34643, N34644, N34646, N34647, N34648, N34649, N34650, N34653, N34655, N34657, N34659, N34660, N34662, N34663, N34665, N34667, N34670, N34671, N34672, N34673, N34674, N34675, N34677, N34678, N34679, N34680, N34681, N34682, N34683, N34685, N34686, N34687, N34688, N34689, N34693, N34697, N34698, N34699, N34701, N34703, N34704, N34705, N34707, N34708, N34711, N34712, N34713, N34719, N34720, N34722, N34724, N34725, N34726, N34727, N34728, N34729, N34730, N34731, N34732, N34735, N34738, N34741, N34742, N34743, N34744, N34745, N34746, N34748, N34749, N34750, N34751, N34752, N34753, N34754, N34756, N34758, N34763, N34764, N34766, N34767, N34769, N34771, N34772, N34773, N34774, N34775, N34777, N34778, N34780, N34781, N34787, N34788, N34789, N34794, N34795, N34796, N34797, N34799, N34800, N34804, N34806, N34807, N34808, N34809, N34810, N34811, N34814, N34815, N34818, N34821, N34822, N34823, N34826, N34827, N34829, N34830, N34831, N34832, N34833, N34836, N34837, N34839, N34840, N34841, N34842, N34844, N34845, N34847, N34848, N34850, N34851, N34853, N34854, N34855, N34856, N34857, N34861, N34863, N34865, N34867, N34868, N34869, N34870, N34871, N34874, N34877, N34878, N34879, N34881, N34882, N34883, N34885, N34886, N34889, N34891, N34893, N34895, N34896, N34897, N34898, N34899, N34900, N34901, N34903, N34904, N34906, N34907, N34908, N34909, N34910, N34911, N34912, N34913, N34914, N34915, N34917, N34918, N34919, N34920, N34921, N34922, N34923, N34925, N34926, N34928, N34929, N34932, N34933, N34934, N34937, N34938, N34939, N34940, N34944, N34945, N34946, N34948, N34951, N34953, N34954, N34956, N34957, N34958, N34959, N34960, N34961, N34962, N34963, N34965, N34967, N34968, N34970, N34977, N34978, N34979, N34982, N34983, N34984, N34985, N34986, N34987, N34988, N34990, N34992, N34993, N34994, N34995, N34996, N34999, N35000, N35001, N35002, N35005, N35006, N35007, N35009, N35013, N35015, N35017, N35018, N35019, N35020, N35021, N35022, N35024, N35025, N35026, N35027, N35028, N35029, N35030, N35032, N35033, N35034, N35035, N35036, N35039, N35042, N35043, N35045, N35046, N35048, N35049, N35050, N35052, N35053, N35054, N35055, N35056, N35057, N35058, N35059, N35060, N35062, N35063, N35064, N35065, N35066, N35067, N35069, N35070, N35071, N35073, N35074, N35077, N35078, N35082, N35083, N35085, N35086, N35087, N35088, N35089, N35091, N35092, N35093, N35095, N35096, N35097, N35098, N35099, N35100, N35101, N35103, N35104, N35107, N35108, N35109, N35110, N35111, N35113, N35115, N35117, N35118, N35119, N35120, N35123, N35125, N35126, N35128, N35129, N35131, N35132, N35133, N35134, N35135, N35136, N35139, N35140, N35143, N35144, N35145, N35146, N35147, N35148, N35149, N35150, N35151, N35152, N35153, N35154, N35155, N35156, N35159, N35160, N35161, N35163, N35166, N35167, N35168, N35169, N35171, N35172, N35173, N35174, N35175, N35176, N35177, N35178, N35179, N35180, N35181, N35185, N35186, N35187, N35188, N35189, N35190, N35191, N35192, N35193, N35196, N35197, N35198, N35199, N35200, N35203, N35204, N35206, N35207, N35208, N35209, N35210, N35211, N35212, N35215, N35217, N35218, N35220, N35221, N35222, N35224, N35225, N35227, N35228, N35230, N35232, N35234, N35236, N35237, N35239, N35240, N35241, N35242, N35244, N35246, N35247, N35248, N35249, N35252, N35253, N35254, N35256, N35257, N35258, N35259, N35260, N35261, N35262, N35263, N35264, N35265, N35266, N35267, N35268, N35269, N35275, N35278, N35279, N35280, N35281, N35282, N35283, N35284, N35286, N35288, N35289, N35290, N35291, N35295, N35296, N35298, N35299, N35300, N35301, N35302, N35304, N35305, N35308, N35309, N35310, N35311, N35313, N35314, N35315, N35318, N35319, N35321, N35322, N35323, N35324, N35326, N35327, N35328, N35330, N35331, N35332, N35333, N35334, N35337, N35338, N35340, N35342, N35343, N35344, N35345, N35346, N35349, N35350, N35351, N35352, N35353, N35354, N35355, N35356, N35357, N35358, N35359, N35362, N35363, N35366, N35368, N35370, N35371, N35373, N35374, N35375, N35376, N35377, N35378, N35379, N35380, N35381, N35383, N35384, N35385, N35386, N35387, N35388, N35389, N35391, N35392, N35394, N35395, N35396, N35398, N35399, N35400, N35401, N35402, N35403, N35406, N35407, N35408, N35409, N35411, N35413, N35414, N35415, N35416, N35417, N35418, N35419, N35422, N35423, N35424, N35425, N35427, N35428, N35429, N35431, N35433, N35435, N35436, N35438, N35439, N35440, N35441, N35442, N35443, N35444, N35445, N35446, N35448, N35449, N35453, N35456, N35457, N35458, N35459, N35460, N35463, N35464, N35467, N35468, N35469, N35470, N35471, N35472, N35474, N35476, N35477, N35479, N35481, N35482, N35485, N35486, N35488, N35490, N35492, N35495, N35496, N35497, N35498, N35499, N35500, N35501, N35502, N35503, N35504, N35507, N35508, N35511, N35512, N35513, N35514, N35516, N35517, N35519, N35521, N35522, N35524, N35525, N35526, N35527, N35529, N35530, N35531, N35532, N35533, N35534, N35536, N35538, N35542, N35544, N35545, N35547, N35548, N35549, N35550, N35551, N35553, N35554, N35555, N35557, N35558, N35560, N35561, N35563, N35564, N35565, N35567, N35569, N35570, N35571, N35573, N35574, N35575, N35576, N35577, N35578, N35579, N35582, N35583, N35584, N35585, N35586, N35587, N35588, N35589, N35591, N35592, N35593, N35594, N35595, N35596, N35598, N35600, N35601, N35603, N35604, N35605, N35606, N35608, N35609, N35611, N35612, N35613, N35615, N35618, N35619, N35620, N35621, N35623, N35624, N35625, N35626, N35627, N35629, N35630, N35631, N35632, N35633, N35635, N35637, N35642, N35643, N35645, N35647, N35649, N35650, N35652, N35653, N35655, N35659, N35661, N35663, N35665, N35666, N35668, N35669, N35670, N35672, N35674, N35675, N35676, N35677, N35678, N35680, N35681, N35682, N35684, N35687, N35690, N35691, N35692, N35694, N35695, N35697, N35698, N35700, N35701, N35702, N35703, N35704, N35705, N35707, N35710, N35711, N35715, N35716, N35718, N35720, N35721, N35722, N35723, N35724, N35725, N35726, N35728, N35731, N35732, N35734, N35735, N35737, N35739, N35740, N35743, N35745, N35747, N35749, N35751, N35752, N35754, N35755, N35756, N35757, N35758, N35759, N35760, N35762, N35764, N35766, N35767, N35768, N35769, N35770, N35771, N35776, N35777, N35779, N35781, N35782, N35785, N35786, N35791, N35793, N35795, N35796, N35797, N35798, N35799, N35800, N35801, N35802, N35803, N35804, N35805, N35806, N35807, N35808, N35811, N35814, N35815, N35816, N35818, N35820, N35821, N35822, N35823, N35828, N35831, N35832, N35833, N35835, N35836, N35837, N35838, N35840, N35841, N35842, N35843, N35844, N35845, N35846, N35847, N35848, N35849, N35851, N35852, N35853, N35855, N35856, N35858, N35860, N35861, N35862, N35863, N35864, N35865, N35868, N35869, N35870, N35872, N35875, N35876, N35878, N35880, N35884, N35885, N35889, N35891, N35892, N35893, N35894, N35895, N35896, N35897, N35898, N35899, N35900, N35901, N35903, N35905, N35906, N35907, N35908, N35910, N35911, N35913, N35914, N35917, N35918, N35919, N35921, N35923, N35924, N35926, N35927, N35929, N35931, N35932, N35933, N35934, N35935, N35936, N35938, N35940, N35941, N35943, N35944, N35947, N35948, N35949, N35950, N35952, N35953, N35954, N35955, N35957, N35958, N35959, N35961, N35962, N35965, N35966, N35971, N35972, N35973, N35974, N35975, N35977, N35979, N35980, N35981, N35982, N35983, N35984, N35986, N35987, N35988, N35989, N35992, N35994, N35995, N35996, N35998, N36000, N36001, N36002, N36003, N36004, N36005, N36006, N36008, N36011, N36013, N36016, N36017, N36019, N36020, N36022, N36024, N36025, N36026, N36027, N36029, N36030, N36031, N36035, N36036, N36037, N36038, N36041, N36042, N36043, N36044, N36047, N36048, N36050, N36051, N36052, N36053, N36055, N36057, N36058, N36059, N36060, N36061, N36063, N36065, N36066, N36068, N36069, N36070, N36072, N36073, N36074, N36076, N36077, N36080, N36081, N36083, N36086, N36087, N36089, N36091, N36092, N36093, N36094, N36097, N36098, N36100, N36102, N36103, N36105, N36106, N36107, N36108, N36109, N36111, N36112, N36113, N36114, N36115, N36116, N36117, N36118, N36121, N36122, N36123, N36124, N36125, N36127, N36130, N36131, N36133, N36134, N36135, N36138, N36139, N36140, N36141, N36143, N36145, N36146, N36148, N36150, N36151, N36153, N36154, N36155, N36158, N36159, N36160, N36161, N36163, N36164, N36169, N36170, N36172, N36174, N36175, N36176, N36177, N36178, N36180, N36181, N36182, N36186, N36187, N36188, N36189, N36191, N36192, N36193, N36194, N36195, N36196, N36197, N36198, N36201, N36202, N36205, N36206, N36209, N36210, N36212, N36214, N36215, N36216, N36219, N36222, N36224, N36225, N36226, N36227, N36228, N36229, N36230, N36231, N36232, N36233, N36234, N36235, N36236, N36238, N36239, N36241, N36242, N36246, N36247, N36249, N36250, N36251, N36252, N36256, N36257, N36259, N36260, N36261, N36262, N36263, N36264, N36265, N36266, N36267, N36271, N36272, N36273, N36274, N36275, N36276, N36277, N36278, N36279, N36281, N36282, N36284, N36285, N36286, N36288, N36289, N36293, N36294, N36295, N36296, N36298, N36300, N36301, N36304, N36307, N36308, N36309, N36313, N36315, N36317, N36318, N36319, N36322, N36325, N36326, N36328, N36329, N36330, N36331, N36333, N36336, N36337, N36338, N36339, N36341, N36342, N36344, N36345, N36346, N36347, N36348, N36351, N36353, N36354, N36355, N36356, N36358, N36362, N36363, N36364, N36365, N36366, N36367, N36368, N36371, N36372, N36373, N36374, N36376, N36378, N36380, N36381, N36383, N36385, N36387, N36388, N36390, N36391, N36393, N36394, N36395, N36396, N36398, N36400, N36401, N36403, N36404, N36406, N36408, N36410, N36412, N36413, N36415, N36416, N36419, N36420, N36421, N36422, N36423, N36424, N36425, N36426, N36427, N36428, N36429, N36430, N36431, N36432, N36433, N36434, N36435, N36436, N36437, N36439, N36442, N36443, N36448, N36451, N36452, N36453, N36455, N36456, N36457, N36458, N36463, N36464, N36465, N36466, N36467, N36468, N36469, N36470, N36471, N36472, N36473, N36474, N36475, N36477, N36478, N36480, N36481, N36482, N36483, N36484, N36488, N36489, N36490, N36491, N36492, N36493, N36497, N36498, N36499, N36500, N36501, N36502, N36503, N36505, N36506, N36507, N36512, N36515, N36516, N36518, N36519, N36521, N36522, N36524, N36525, N36526, N36527, N36528, N36529, N36531, N36532, N36534, N36536, N36537, N36539, N36540, N36542, N36543, N36545, N36546, N36548, N36549, N36552, N36553, N36554, N36556, N36557, N36558, N36560, N36561, N36562, N36563, N36564, N36565, N36566, N36567, N36569, N36570, N36571, N36575, N36576, N36577, N36578, N36580, N36583, N36584, N36585, N36587, N36588, N36592, N36594, N36595, N36596, N36597, N36598, N36599, N36600, N36601, N36602, N36603, N36604, N36605, N36607, N36608, N36609, N36610, N36611, N36613, N36615, N36617, N36618, N36619, N36621, N36622, N36623, N36624, N36625, N36626, N36627, N36629, N36630, N36633, N36634, N36635, N36636, N36638, N36639, N36640, N36642, N36644, N36645, N36646, N36647, N36649, N36650, N36651, N36653, N36654, N36655, N36656, N36657, N36661, N36662, N36663, N36664, N36665, N36666, N36667, N36668, N36669, N36671, N36672, N36673, N36674, N36675, N36677, N36678, N36679, N36680, N36682, N36683, N36684, N36686, N36687, N36688, N36689, N36691, N36695, N36697, N36699, N36701, N36702, N36703, N36705, N36706, N36707, N36709, N36711, N36713, N36715, N36716, N36717, N36718, N36719, N36720, N36721, N36722, N36723, N36724, N36725, N36727, N36729, N36730, N36733, N36734, N36735, N36737, N36738, N36740, N36742, N36743, N36744, N36746, N36747, N36748, N36749, N36752, N36754, N36755, N36756, N36758, N36760, N36764, N36765, N36767, N36768, N36769, N36770, N36771, N36773, N36774, N36777, N36778, N36779, N36780, N36782, N36783, N36784, N36785, N36786, N36787, N36788, N36789, N36791, N36793, N36795, N36797, N36798, N36799, N36803, N36804, N36805, N36806, N36807, N36808, N36809, N36810, N36811, N36812, N36813, N36816, N36817, N36818, N36820, N36821, N36822, N36823, N36824, N36825, N36828, N36829, N36831, N36834, N36835, N36839, N36840, N36842, N36845, N36846, N36848, N36850, N36851, N36852, N36853, N36854, N36855, N36858, N36859, N36861, N36862, N36863, N36864, N36865, N36866, N36867, N36869, N36870, N36871, N36872, N36873, N36874, N36879, N36880, N36881, N36882, N36886, N36887, N36888, N36889, N36890, N36891, N36892, N36893, N36896, N36897, N36898, N36900, N36902, N36906, N36907, N36908, N36909, N36910, N36911, N36912, N36915, N36916, N36917, N36918, N36920, N36921, N36922, N36923, N36925, N36926, N36928, N36929, N36930, N36931, N36932, N36933, N36934, N36936, N36937, N36938, N36939, N36946, N36948, N36949, N36950, N36951, N36952, N36954, N36955, N36956, N36958, N36959, N36960, N36961, N36962, N36964, N36967, N36970, N36972, N36977, N36978, N36980, N36981, N36982, N36985, N36990, N36991, N36992, N36995, N36998, N36999, N37000, N37001, N37002, N37003, N37004, N37006, N37011, N37013, N37014, N37016, N37017, N37018, N37019, N37020, N37021, N37023, N37024, N37025, N37026, N37028, N37029, N37031, N37032, N37035, N37037, N37038, N37039, N37042, N37043, N37044, N37046, N37048, N37052, N37053, N37054, N37055, N37059, N37061, N37063, N37065, N37066, N37067, N37068, N37070, N37071, N37075, N37079, N37083, N37084, N37085, N37087, N37088, N37089, N37090, N37091, N37092, N37093, N37094, N37097, N37099, N37100, N37103, N37108, N37109, N37111, N37113, N37115, N37117, N37120, N37121, N37123, N37124, N37125, N37128, N37131, N37137, N37139, N37140, N37141, N37142, N37144, N37145, N37148, N37149, N37150, N37152, N37153, N37154, N37155, N37156, N37157, N37158, N37159, N37161, N37162, N37163, N37164, N37165, N37166, N37167, N37169, N37170, N37171, N37173, N37176, N37177, N37179, N37180, N37181, N37182, N37185, N37186, N37187, N37192, N37193, N37194, N37195, N37196, N37197, N37198, N37199, N37200, N37201, N37202, N37204, N37205, N37206, N37211, N37212, N37213, N37214, N37215, N37216, N37218, N37220, N37222, N37226, N37228, N37230, N37231, N37232, N37234, N37235, N37237, N37238, N37239, N37242, N37243, N37244, N37245, N37247, N37248, N37249, N37251, N37252, N37253, N37254, N37256, N37260, N37264, N37265, N37266, N37267, N37269, N37271, N37272, N37273, N37274, N37275, N37276, N37277, N37278, N37279, N37280, N37282, N37284, N37285, N37286, N37288, N37289, N37290, N37294, N37297, N37299, N37300, N37302, N37304, N37305, N37306, N37307, N37308, N37309, N37310, N37311, N37312, N37313, N37316, N37319, N37320, N37321, N37322, N37324, N37325, N37326, N37327, N37328, N37331, N37334, N37335, N37336, N37338, N37339, N37341, N37342, N37343, N37345, N37346, N37347, N37348, N37349, N37350, N37351, N37352, N37353, N37354, N37355, N37358, N37359, N37360, N37363, N37365, N37366, N37368, N37371, N37373, N37374, N37375, N37376, N37377, N37378, N37379, N37380, N37381, N37382, N37383, N37386, N37387, N37388, N37389, N37390, N37391, N37392, N37393, N37394, N37399, N37401, N37402, N37403, N37404, N37405, N37407, N37408, N37409, N37410, N37411, N37414, N37415, N37417, N37418, N37419, N37420, N37421, N37424, N37425, N37426, N37427, N37428, N37430, N37432, N37433, N37434, N37435, N37437, N37438, N37439, N37440, N37442, N37443, N37444, N37445, N37446, N37448, N37450, N37453, N37454, N37455, N37457, N37460, N37463, N37464, N37466, N37467, N37469, N37470, N37475, N37477, N37479, N37480, N37481, N37482, N37483, N37485, N37486, N37488, N37490, N37492, N37496, N37497, N37498, N37500, N37501, N37502, N37503, N37504, N37505, N37506, N37508, N37509, N37512, N37513, N37514, N37515, N37517, N37518, N37519, N37520, N37521, N37523, N37524, N37526, N37527, N37528, N37529, N37531, N37532, N37533, N37534, N37535, N37536, N37537, N37538, N37540, N37542, N37543, N37545, N37546, N37547, N37548, N37549, N37550, N37551, N37552, N37553, N37554, N37556, N37557, N37558, N37559, N37563, N37564, N37565, N37566, N37571, N37572, N37573, N37574, N37575, N37576, N37578, N37579, N37580, N37581, N37582, N37583, N37584, N37585, N37586, N37588, N37590, N37591, N37592, N37593, N37595, N37596, N37598, N37600, N37601, N37602, N37603, N37604, N37605, N37607, N37608, N37609, N37610, N37611, N37612, N37613, N37614, N37616, N37617, N37618, N37620, N37621, N37622, N37623, N37624, N37625, N37628, N37629, N37630, N37631, N37632, N37633, N37635, N37636, N37638, N37639, N37643, N37644, N37645, N37646, N37647, N37648, N37649, N37650, N37651, N37654, N37655, N37656, N37658, N37659, N37660, N37661, N37663, N37664, N37666, N37668, N37670, N37671, N37672, N37673, N37674, N37677, N37678, N37680, N37684, N37687, N37688, N37690, N37691, N37692, N37693, N37695, N37696, N37697, N37701, N37705, N37707, N37708, N37709, N37710, N37711, N37712, N37713, N37714, N37715, N37716, N37717, N37720, N37723, N37724, N37726, N37727, N37728, N37729, N37730, N37731, N37734, N37736, N37737, N37738, N37739, N37740, N37742, N37743, N37745, N37746, N37747, N37748, N37749, N37750, N37751, N37752, N37753, N37754, N37756, N37757, N37759, N37761, N37763, N37764, N37766, N37768, N37769, N37770, N37772, N37773, N37774, N37775, N37776, N37777, N37778, N37779, N37780, N37781, N37782, N37783, N37786, N37788, N37789, N37790, N37791, N37792, N37793, N37795, N37796, N37797, N37798, N37803, N37804, N37806, N37807, N37808, N37809, N37811, N37813, N37814, N37816, N37819, N37820, N37826, N37827, N37828, N37830, N37831, N37832, N37833, N37837, N37838, N37840, N37841, N37844, N37846, N37847, N37851, N37852, N37853, N37854, N37855, N37857, N37858, N37859, N37860, N37861, N37862, N37863, N37864, N37865, N37866, N37867, N37868, N37869, N37871, N37872, N37874, N37875, N37876, N37877, N37878, N37879, N37882, N37884, N37885, N37887, N37888, N37889, N37890, N37891, N37892, N37893, N37894, N37895, N37896, N37898, N37900, N37903, N37904, N37905, N37907, N37908, N37909, N37911, N37912, N37913, N37914, N37915, N37917, N37918, N37919, N37920, N37921, N37922, N37923, N37924, N37927, N37928, N37929, N37930, N37932, N37933, N37934, N37935, N37937, N37938, N37939, N37940, N37941, N37943, N37944, N37945, N37946, N37948, N37949, N37950, N37952, N37953, N37957, N37959, N37960, N37961, N37964, N37965, N37966, N37967, N37968, N37969, N37970, N37971, N37972, N37973, N37977, N37979, N37980, N37981, N37982, N37983, N37986, N37987, N37988, N37989, N37990, N37994, N37998, N37999, N38000, N38003, N38005, N38006, N38009, N38010, N38011, N38012, N38015, N38016, N38017, N38019, N38022, N38023, N38024, N38025, N38026, N38027, N38029, N38030, N38031, N38032, N38033, N38034, N38035, N38040, N38041, N38043, N38045, N38046, N38047, N38048, N38049, N38050, N38051, N38052, N38053, N38054, N38055, N38056, N38057, N38059, N38062, N38063, N38064, N38065, N38066, N38067, N38069, N38071, N38074, N38075, N38077, N38078, N38080, N38082, N38083, N38084, N38088, N38090, N38091, N38092, N38093, N38094, N38095, N38096, N38097, N38098, N38099, N38100, N38103, N38104, N38105, N38108, N38109, N38111, N38113, N38114, N38116, N38117, N38118, N38119, N38121, N38122, N38124, N38125, N38126, N38127, N38128, N38129, N38132, N38133, N38134, N38135, N38136, N38137, N38139, N38141, N38142, N38143, N38144, N38145, N38146, N38147, N38148, N38149, N38150, N38151, N38152, N38153, N38154, N38155, N38157, N38159, N38160, N38161, N38163, N38164, N38166, N38168, N38171, N38175, N38177, N38178, N38179, N38182, N38183, N38186, N38187, N38188, N38189, N38190, N38191, N38192, N38193, N38194, N38196, N38197, N38199, N38202, N38204, N38205, N38206, N38207, N38209, N38210, N38212, N38213, N38217, N38218, N38220, N38221, N38222, N38224, N38225, N38226, N38227, N38228, N38230, N38232, N38233, N38234, N38235, N38237, N38238, N38240, N38243, N38245, N38246, N38247, N38248, N38249, N38250, N38255, N38259, N38260, N38261, N38262, N38263, N38264, N38267, N38268, N38270, N38271, N38275, N38276, N38277, N38278, N38279, N38281, N38283, N38284, N38285, N38287, N38288, N38289, N38290, N38293, N38294, N38296, N38297, N38299, N38302, N38304, N38305, N38307, N38308, N38309, N38312, N38313, N38314, N38315, N38316, N38318, N38319, N38321, N38322, N38324, N38325, N38326, N38328, N38329, N38331, N38332, N38335, N38336, N38337, N38338, N38339, N38340, N38341, N38342, N38345, N38346, N38349, N38350, N38351, N38353, N38354, N38359, N38360, N38362, N38365, N38368, N38369, N38371, N38372, N38374, N38375, N38376, N38378, N38379, N38380, N38381, N38384, N38385, N38386, N38387, N38388, N38389, N38391, N38392, N38393, N38394, N38396, N38397, N38398, N38399, N38400, N38402, N38403, N38404, N38405, N38407, N38408, N38409, N38410, N38411, N38412, N38413, N38415, N38416, N38418, N38419, N38421, N38422, N38423, N38424, N38426, N38427, N38428, N38429, N38430, N38431, N38433, N38434, N38435, N38436, N38437, N38438, N38439, N38440, N38443, N38444, N38445, N38446, N38447, N38448, N38449, N38452, N38453, N38454, N38455, N38458, N38459, N38460, N38461, N38462, N38464, N38465, N38467, N38468, N38469, N38470, N38471, N38472, N38473, N38474, N38476, N38478, N38479, N38480, N38482, N38483, N38486, N38487, N38488, N38489, N38493, N38494, N38495, N38496, N38497, N38498, N38501, N38504, N38505, N38506, N38507, N38508, N38509, N38510, N38511, N38512, N38515, N38517, N38518, N38520, N38521, N38522, N38524, N38525, N38527, N38528, N38530, N38531, N38533, N38535, N38536, N38538, N38539, N38540, N38541, N38542, N38544, N38545, N38546, N38547, N38548, N38549, N38550, N38551, N38552, N38553, N38555, N38556, N38557, N38558, N38559, N38561, N38562, N38563, N38567, N38569, N38570, N38571, N38572, N38573, N38574, N38575, N38576, N38577, N38579, N38580, N38582, N38583, N38585, N38586, N38587, N38588, N38589, N38591, N38596, N38597, N38598, N38599, N38602, N38604, N38608, N38609, N38614, N38615, N38616, N38618, N38619, N38620, N38622, N38623, N38627, N38628, N38629, N38630, N38631, N38632, N38633, N38634, N38636, N38637, N38638, N38639, N38643, N38646, N38648, N38650, N38652, N38653, N38654, N38655, N38656, N38657, N38658, N38659, N38660, N38662, N38663, N38664, N38665, N38667, N38668, N38669, N38670, N38671, N38672, N38674, N38675, N38676, N38679, N38680, N38682, N38684, N38686, N38687, N38688, N38689, N38695, N38696, N38697, N38699, N38700, N38704, N38705, N38707, N38708, N38710, N38712, N38713, N38714, N38715, N38717, N38718, N38719, N38720, N38721, N38722, N38723, N38725, N38726, N38728, N38730, N38731, N38733, N38734, N38736, N38737, N38739, N38740, N38741, N38744, N38746, N38747, N38749, N38750, N38751, N38753, N38755, N38756, N38757, N38758, N38759, N38761, N38762, N38764, N38765, N38766, N38767, N38768, N38769, N38770, N38771, N38772, N38775, N38776, N38778, N38779, N38780, N38781, N38782, N38784, N38785, N38786, N38788, N38791, N38792, N38793, N38794, N38795, N38796, N38798, N38801, N38802, N38803, N38805, N38806, N38808, N38812, N38813, N38815, N38817, N38819, N38821, N38823, N38826, N38827, N38829, N38830, N38832, N38834, N38835, N38836, N38838, N38840, N38841, N38842, N38844, N38845, N38849, N38850, N38851, N38853, N38856, N38857, N38858, N38859, N38862, N38865, N38867, N38868, N38869, N38870, N38874, N38876, N38877, N38880, N38882, N38883, N38884, N38885, N38886, N38887, N38888, N38889, N38890, N38891, N38892, N38893, N38895, N38897, N38898, N38901, N38903, N38904, N38905, N38906, N38907, N38910, N38911, N38913, N38914, N38915, N38916, N38917, N38918, N38919, N38920, N38921, N38922, N38923, N38924, N38925, N38926, N38928, N38931, N38932, N38933, N38934, N38937, N38938, N38939, N38940, N38941, N38944, N38946, N38947, N38949, N38950, N38951, N38952, N38953, N38954, N38956, N38957, N38960, N38961, N38962, N38964, N38966, N38967, N38968, N38970, N38971, N38972, N38974, N38976, N38977, N38980, N38984, N38986, N38987, N38990, N38993, N38994, N38999, N39000, N39001, N39002, N39003, N39005, N39007, N39008, N39010, N39011, N39014, N39016, N39017, N39019, N39020, N39021, N39023, N39024, N39025, N39026, N39028, N39029, N39030, N39031, N39033, N39034, N39035, N39036, N39037, N39038, N39041, N39042, N39043, N39044, N39045, N39046, N39047, N39048, N39049, N39050, N39051, N39053, N39054, N39055, N39057, N39059, N39060, N39061, N39062, N39063, N39064, N39065, N39066, N39068, N39069, N39070, N39071, N39073, N39074, N39076, N39077, N39078, N39079, N39081, N39082, N39084, N39086, N39089, N39090, N39091, N39092, N39093, N39097, N39098, N39101, N39102, N39103, N39104, N39105, N39106, N39107, N39108, N39109, N39110, N39111, N39112, N39117, N39119, N39122, N39123, N39124, N39125, N39126, N39128, N39129, N39131, N39132, N39133, N39134, N39135, N39136, N39137, N39139, N39142, N39143, N39144, N39148, N39149, N39151, N39153, N39154, N39155, N39156, N39157, N39160, N39161, N39163, N39164, N39165, N39166, N39168, N39169, N39170, N39171, N39172, N39173, N39175, N39176, N39177, N39178, N39181, N39182, N39184, N39185, N39186, N39187, N39188, N39190, N39194, N39195, N39196, N39197, N39200, N39201, N39203, N39204, N39206, N39208, N39209, N39211, N39213, N39214, N39216, N39217, N39218, N39219, N39220, N39222, N39223, N39224, N39225, N39227, N39228, N39229, N39230, N39233, N39234, N39236, N39238, N39241, N39242, N39243, N39244, N39247, N39248, N39249, N39250, N39251, N39252, N39253, N39255, N39257, N39258, N39260, N39261, N39262, N39267, N39268, N39270, N39271, N39272, N39273, N39274, N39277, N39278, N39281, N39283, N39284, N39285, N39286, N39287, N39289, N39290, N39291, N39293, N39294, N39295, N39297, N39298, N39299, N39301, N39303, N39304, N39305, N39306, N39308, N39310, N39311, N39316, N39318, N39320, N39321, N39322, N39324, N39325, N39327, N39328, N39329, N39330, N39331, N39332, N39334, N39335, N39336, N39337, N39338, N39339, N39340, N39342, N39345, N39347, N39348, N39351, N39352, N39353, N39354, N39357, N39358, N39359, N39360, N39361, N39366, N39368, N39369, N39372, N39373, N39375, N39376, N39378, N39379, N39380, N39383, N39384, N39388, N39389, N39390, N39391, N39393, N39394, N39395, N39396, N39398, N39401, N39403, N39404, N39406, N39407, N39409, N39410, N39411, N39413, N39414, N39417, N39418, N39419, N39420, N39421, N39422, N39423, N39425, N39429, N39431, N39432, N39433, N39436, N39437, N39438, N39439, N39440, N39441, N39442, N39443, N39444, N39445, N39450, N39451, N39452, N39453, N39456, N39459, N39461, N39463, N39465, N39467, N39468, N39472, N39473, N39475, N39477, N39480, N39482, N39484, N39485, N39486, N39487, N39488, N39489, N39490, N39491, N39494, N39496, N39497, N39499, N39500, N39501, N39502, N39503, N39506, N39507, N39508, N39509, N39511, N39512, N39516, N39517, N39519, N39521, N39522, N39524, N39526, N39527, N39528, N39530, N39531, N39533, N39534, N39535, N39536, N39537, N39539, N39540, N39543, N39544, N39545, N39547, N39548, N39551, N39552, N39553, N39554, N39555, N39556, N39557, N39558, N39560, N39561, N39563, N39564, N39565, N39566, N39567, N39568, N39569, N39570, N39571, N39572, N39573, N39574, N39575, N39576, N39578, N39579, N39581, N39582, N39584, N39586, N39587, N39588, N39589, N39591, N39592, N39593, N39595, N39596, N39598, N39602, N39603, N39606, N39608, N39609, N39610, N39611, N39613, N39615, N39616, N39617, N39618, N39621, N39622, N39623, N39624, N39625, N39626, N39627, N39628, N39629, N39631, N39633, N39634, N39635, N39636, N39637, N39638, N39642, N39643, N39645, N39646, N39647, N39649, N39653, N39654, N39656, N39658, N39661, N39662, N39663, N39664, N39666, N39669, N39672, N39674, N39679, N39680, N39681, N39682, N39685, N39686, N39687, N39692, N39695, N39697, N39698, N39699, N39700, N39701, N39702, N39703, N39704, N39706, N39707, N39708, N39709, N39711, N39713, N39714, N39715, N39717, N39718, N39720, N39721, N39722, N39724, N39725, N39726, N39727, N39729, N39730, N39731, N39733, N39734, N39736, N39737, N39740, N39741, N39743, N39745, N39748, N39751, N39754, N39755, N39756, N39757, N39758, N39759, N39760, N39761, N39763, N39765, N39766, N39768, N39770, N39771, N39773, N39776, N39778, N39779, N39781, N39782, N39783, N39786, N39787, N39788, N39789, N39790, N39791, N39792, N39793, N39794, N39795, N39797, N39798, N39800, N39801, N39803, N39804, N39805, N39806, N39808, N39809, N39810, N39811, N39813, N39814, N39815, N39816, N39817, N39818, N39820, N39821, N39822, N39823, N39825, N39827, N39828, N39830, N39831, N39833, N39834, N39837, N39838, N39839, N39841, N39842, N39843, N39846, N39847, N39848, N39849, N39850, N39851, N39852, N39853, N39854, N39855, N39856, N39860, N39862, N39863, N39864, N39865, N39866, N39867, N39868, N39870, N39871, N39872, N39875, N39876, N39877, N39879, N39880, N39882, N39883, N39884, N39885, N39886, N39889, N39890, N39892, N39894, N39895, N39896, N39897, N39899, N39901, N39902, N39904, N39905, N39906, N39907, N39910, N39912, N39913, N39914, N39915, N39917, N39918, N39920, N39921, N39922, N39923, N39924, N39925, N39926, N39927, N39928, N39929, N39930, N39931, N39933, N39935, N39936, N39939, N39940, N39942, N39944, N39946, N39948, N39950, N39951, N39952, N39954, N39955, N39956, N39957, N39959, N39960, N39961, N39962, N39963, N39965, N39966, N39968, N39969, N39972, N39973, N39974, N39975, N39976, N39977, N39978, N39980, N39982, N39984, N39985, N39987, N39988, N39990, N39991, N39992, N39993, N39994, N39995, N39996, N39999, N40001, N40003, N40005, N40006, N40007, N40008, N40009, N40011, N40013, N40014, N40016, N40017, N40019, N40023, N40024, N40027, N40028, N40031, N40032, N40036, N40037, N40038, N40039, N40044, N40046, N40047, N40048, N40051, N40052, N40053, N40054, N40055, N40056, N40057, N40058, N40061, N40062, N40063, N40064, N40066, N40068, N40069, N40070, N40071, N40073, N40074, N40076, N40077, N40078, N40080, N40081, N40082, N40083, N40084, N40085, N40088, N40089, N40090, N40091, N40092, N40094, N40096, N40099, N40101, N40102, N40103, N40104, N40106, N40107, N40108, N40109, N40111, N40112, N40114, N40115, N40116, N40118, N40119, N40120, N40121, N40124, N40125, N40126, N40127, N40128, N40129, N40133, N40134, N40136, N40137, N40138, N40139, N40142, N40143, N40144, N40145, N40147, N40148, N40152, N40153, N40154, N40155, N40156, N40157, N40158, N40159, N40160, N40161, N40164, N40166, N40168, N40169, N40170, N40171, N40172, N40173, N40174, N40176, N40177, N40178, N40179, N40180, N40181, N40188, N40191, N40192, N40196, N40199, N40200, N40201, N40202, N40204, N40205, N40206, N40207, N40208, N40209, N40210, N40211, N40212, N40213, N40214, N40216, N40217, N40218, N40220, N40221, N40222, N40223, N40225, N40227, N40229, N40230, N40231, N40232, N40233, N40234, N40236, N40237, N40238, N40239, N40240, N40242, N40244, N40245, N40247, N40248, N40249, N40250, N40252, N40253, N40254, N40258, N40259, N40260, N40261, N40263, N40267, N40268, N40270, N40272, N40274, N40275, N40276, N40278, N40279, N40280, N40281, N40282, N40284, N40287, N40288, N40289, N40291, N40294, N40296, N40299, N40300, N40301, N40302, N40303, N40306, N40307, N40308, N40309, N40311, N40313, N40314, N40315, N40316, N40318, N40319, N40320, N40321, N40322, N40324, N40325, N40326, N40329, N40330, N40331, N40332, N40333, N40334, N40335, N40336, N40338, N40339, N40341, N40342, N40344, N40345, N40346, N40347, N40348, N40349, N40350, N40351, N40352, N40353, N40354, N40355, N40357, N40358, N40360, N40361, N40362, N40363, N40364, N40365, N40367, N40369, N40370, N40371, N40372, N40373, N40375, N40376, N40377, N40379, N40381, N40382, N40384, N40385, N40386, N40389, N40390, N40392, N40393, N40394, N40396, N40397, N40398, N40399, N40400, N40404, N40405, N40406, N40408, N40409, N40410, N40412, N40413, N40415, N40416, N40417, N40418, N40420, N40421, N40422, N40423, N40424, N40425, N40427, N40428, N40433, N40434, N40435, N40436, N40437, N40438, N40439, N40441, N40443, N40444, N40445, N40446, N40447, N40450, N40452, N40454, N40455, N40456, N40457, N40458, N40459, N40461, N40462, N40464, N40465, N40466, N40467, N40468, N40469, N40470, N40472, N40474, N40477, N40478, N40479, N40481, N40483, N40484, N40486, N40488, N40489, N40490, N40491, N40492, N40493, N40494, N40495, N40497, N40498, N40499, N40500, N40502, N40505, N40506, N40507, N40509, N40510, N40511, N40513, N40514, N40516, N40517, N40518, N40522, N40523, N40525, N40526, N40527, N40528, N40530, N40531, N40533, N40535, N40537, N40542, N40544, N40545, N40546, N40547, N40549, N40550, N40551, N40552, N40553, N40554, N40557, N40558, N40560, N40561, N40562, N40563, N40564, N40565, N40566, N40567, N40568, N40571, N40573, N40574, N40575, N40577, N40578, N40579, N40583, N40585, N40587, N40589, N40590, N40591, N40592, N40594, N40595, N40596, N40598, N40599, N40601, N40602, N40604, N40605, N40607, N40608, N40610, N40612, N40613, N40614, N40615, N40616, N40617, N40618, N40619, N40620, N40621, N40626, N40627, N40630, N40631, N40632, N40633, N40634, N40636, N40637, N40640, N40642, N40645, N40647, N40648, N40649, N40650, N40654, N40655, N40657, N40658, N40659, N40661, N40662, N40664, N40665, N40668, N40670, N40671, N40673, N40675, N40676, N40677, N40678, N40680, N40681, N40682, N40683, N40684, N40685, N40686, N40687, N40688, N40691, N40693, N40694, N40695, N40696, N40697, N40698, N40699, N40700, N40701, N40702, N40708, N40709, N40710, N40711, N40712, N40713, N40714, N40715, N40716, N40719, N40720, N40721, N40722, N40723, N40724, N40728, N40729, N40731, N40732, N40733, N40735, N40736, N40738, N40739, N40740, N40742, N40744, N40746, N40747, N40748, N40749, N40750, N40756, N40757, N40758, N40760, N40761, N40762, N40763, N40766, N40767, N40768, N40769, N40770, N40771, N40772, N40773, N40775, N40776, N40778, N40779, N40780, N40786, N40787, N40788, N40789, N40790, N40791, N40793, N40794, N40795, N40797, N40798, N40801, N40804, N40805, N40809, N40810, N40811, N40813, N40816, N40822, N40823, N40826, N40827, N40828, N40829, N40830, N40831, N40832, N40833, N40834, N40836, N40837, N40838, N40839, N40840, N40841, N40843, N40844, N40845, N40846, N40849, N40850, N40852, N40854, N40855, N40856, N40857, N40858, N40859, N40860, N40861, N40862, N40863, N40865, N40866, N40868, N40869, N40870, N40871, N40872, N40875, N40876, N40878, N40879, N40880, N40886, N40888, N40892, N40893, N40896, N40899, N40902, N40903, N40904, N40905, N40906, N40907, N40908, N40909, N40910, N40911, N40913, N40915, N40917, N40919, N40920, N40922, N40923, N40924, N40926, N40929, N40930, N40931, N40933, N40934, N40935, N40936, N40937, N40939, N40940, N40942, N40944, N40945, N40946, N40947, N40949, N40950, N40954, N40955, N40956, N40957, N40959, N40960, N40961, N40962, N40963, N40965, N40969, N40971, N40973, N40974, N40978, N40979, N40981, N40983, N40984, N40986, N40987, N40989, N40990, N40991, N40993, N40994, N40995, N40997, N40998, N40999, N41000, N41003, N41006, N41008, N41010, N41012, N41013, N41017, N41018, N41020, N41021, N41022, N41023, N41024, N41026, N41027, N41028, N41029, N41031, N41032, N41033, N41034, N41035, N41036, N41037, N41038, N41039, N41041, N41043, N41045, N41046, N41047, N41048, N41049, N41050, N41052, N41053, N41054, N41055, N41057, N41059, N41060, N41062, N41063, N41064, N41065, N41066, N41067, N41068, N41069, N41070, N41071, N41072, N41073, N41074, N41075, N41076, N41078, N41079, N41080, N41081, N41083, N41084, N41085, N41088, N41093, N41094, N41095, N41096, N41097, N41098, N41100, N41101, N41103, N41104, N41105, N41106, N41107, N41108, N41110, N41111, N41114, N41115, N41117, N41119, N41120, N41121, N41122, N41123, N41124, N41127, N41128, N41129, N41130, N41131, N41132, N41134, N41135, N41136, N41138, N41139, N41144, N41145, N41146, N41147, N41148, N41149, N41150, N41151, N41152, N41153, N41154, N41159, N41160, N41161, N41162, N41165, N41166, N41167, N41168, N41170, N41171, N41172, N41173, N41174, N41176, N41178, N41179, N41181, N41182, N41183, N41184, N41185, N41186, N41187, N41189, N41190, N41193, N41194, N41195, N41196, N41199, N41200, N41201, N41202, N41204, N41208, N41209, N41210, N41211, N41212, N41213, N41214, N41215, N41216, N41219, N41220, N41223, N41224, N41225, N41226, N41227, N41228, N41229, N41232, N41234, N41235, N41236, N41237, N41239, N41240, N41242, N41244, N41246, N41247, N41248, N41249, N41250, N41252, N41253, N41255, N41256, N41257, N41259, N41260, N41262, N41263, N41265, N41266, N41267, N41271, N41273, N41276, N41278, N41279, N41280, N41282, N41283, N41284, N41285, N41286, N41287, N41289, N41290, N41293, N41294, N41295, N41296, N41297, N41299, N41300, N41302, N41303, N41304, N41305, N41306, N41309, N41310, N41311, N41312, N41313, N41315, N41316, N41318, N41319, N41321, N41322, N41323, N41324, N41325, N41329, N41330, N41331, N41333, N41334, N41336, N41337, N41339, N41341, N41342, N41343, N41344, N41348, N41349, N41350, N41352, N41353, N41354, N41355, N41356, N41357, N41359, N41360, N41362, N41363, N41364, N41367, N41368, N41369, N41371, N41372, N41373, N41374, N41375, N41376, N41377, N41378, N41379, N41380, N41381, N41382, N41384, N41386, N41387, N41388, N41389, N41390, N41391, N41392, N41393, N41394, N41395, N41397, N41399, N41400, N41401, N41403, N41404, N41405, N41406, N41407, N41409, N41410, N41412, N41414, N41415, N41417, N41418, N41419, N41421, N41424, N41425, N41426, N41428, N41430, N41431, N41432, N41433, N41434, N41435, N41437, N41438, N41439, N41440, N41441, N41443, N41445, N41446, N41450, N41452, N41453, N41456, N41457, N41458, N41459, N41460, N41461, N41462, N41464, N41466, N41467, N41470, N41471, N41473, N41474, N41476, N41479, N41481, N41483, N41484, N41486, N41489, N41490, N41491, N41493, N41494, N41495, N41496, N41497, N41499, N41500, N41504, N41505, N41506, N41511, N41512, N41513, N41514, N41515, N41518, N41519, N41520, N41521, N41522, N41525, N41526, N41527, N41528, N41529, N41530, N41531, N41532, N41536, N41537, N41540, N41541, N41542, N41543, N41544, N41545, N41547, N41549, N41550, N41551, N41552, N41553, N41554, N41555, N41556, N41558, N41559, N41560, N41561, N41562, N41564, N41565, N41566, N41567, N41568, N41569, N41570, N41571, N41572, N41573, N41574, N41575, N41576, N41577, N41578, N41579, N41580, N41582, N41583, N41584, N41586, N41587, N41588, N41589, N41590, N41591, N41593, N41595, N41596, N41597, N41598, N41600, N41601, N41603, N41604, N41606, N41607, N41608, N41609, N41612, N41613, N41616, N41619, N41621, N41622, N41623, N41628, N41632, N41633, N41636, N41638, N41639, N41640, N41642, N41643, N41645, N41646, N41649, N41650, N41651, N41652, N41654, N41655, N41657, N41658, N41659, N41660, N41661, N41662, N41664, N41665, N41666, N41667, N41668, N41669, N41670, N41671, N41673, N41674, N41675, N41679, N41680, N41681, N41685, N41687, N41692, N41695, N41697, N41698, N41699, N41700, N41701, N41707, N41708, N41709, N41710, N41712, N41714, N41715, N41716, N41717, N41720, N41724, N41725, N41726, N41727, N41728, N41731, N41732, N41733, N41736, N41737, N41741, N41743, N41745, N41749, N41750, N41751, N41752, N41753, N41754, N41758, N41759, N41760, N41761, N41763, N41764, N41765, N41766, N41767, N41768, N41769, N41770, N41775, N41776, N41777, N41778, N41781, N41783, N41786, N41787, N41788, N41792, N41793, N41795, N41796, N41797, N41798, N41800, N41802, N41803, N41804, N41805, N41806, N41807, N41810, N41811, N41812, N41813, N41814, N41815, N41818, N41820, N41822, N41823, N41827, N41829, N41830, N41831, N41832, N41833, N41835, N41836, N41837, N41838, N41839, N41840, N41842, N41843, N41844, N41845, N41846, N41848, N41849, N41851, N41856, N41859, N41860, N41861, N41862, N41865, N41866, N41867, N41869, N41871, N41873, N41874, N41875, N41876, N41877, N41878, N41880, N41881, N41882, N41883, N41885, N41887, N41888, N41889, N41890, N41891, N41892, N41893, N41894, N41895, N41896, N41897, N41898, N41899, N41900, N41901, N41902, N41903, N41904, N41906, N41907, N41908, N41910, N41911, N41912, N41915, N41916, N41917, N41918, N41919, N41920, N41921, N41923, N41924, N41927, N41929, N41931, N41932, N41933, N41935, N41936, N41937, N41938, N41941, N41942, N41943, N41944, N41945, N41947, N41948, N41950, N41951, N41952, N41953, N41956, N41957, N41958, N41959, N41960, N41962, N41964, N41965, N41966, N41968, N41969, N41970, N41972, N41973, N41975, N41977, N41979, N41980, N41982, N41983, N41984, N41985, N41986, N41988, N41990, N41991, N41992, N41993, N41994, N41995, N41996, N41998, N42000, N42001, N42002, N42003, N42004, N42005, N42006, N42008, N42011, N42012, N42013, N42014, N42015, N42016, N42018, N42019, N42020, N42022, N42024, N42025, N42026, N42028, N42029, N42030, N42031, N42033, N42035, N42039, N42040, N42041, N42045, N42047, N42051, N42054, N42055, N42056, N42059, N42061, N42062, N42064, N42066, N42068, N42069, N42070, N42071, N42072, N42074, N42076, N42078, N42080, N42082, N42084, N42085, N42086, N42087, N42088, N42089, N42091, N42092, N42094, N42095, N42096, N42097, N42100, N42101, N42103, N42104, N42105, N42106, N42107, N42108, N42109, N42110, N42113, N42114, N42115, N42116, N42118, N42125, N42127, N42128, N42129, N42131, N42132, N42133, N42136, N42138, N42140, N42141, N42142, N42144, N42145, N42146, N42149, N42150, N42151, N42152, N42153, N42154, N42156, N42158, N42160, N42162, N42164, N42168, N42169, N42170, N42174, N42175, N42176, N42177, N42178, N42180, N42181, N42182, N42185, N42186, N42187, N42188, N42189, N42191, N42192, N42194, N42195, N42197, N42198, N42199, N42200, N42201, N42203, N42204, N42206, N42207, N42208, N42209, N42210, N42211, N42212, N42213, N42214, N42217, N42218, N42219, N42220, N42221, N42222, N42224, N42225, N42227, N42229, N42230, N42232, N42233, N42234, N42235, N42237, N42238, N42240, N42241, N42242, N42243, N42245, N42246, N42247, N42248, N42249, N42250, N42252, N42254, N42255, N42256, N42257, N42258, N42259, N42260, N42262, N42263, N42264, N42265, N42267, N42269, N42270, N42271, N42272, N42273, N42276, N42279, N42280, N42281, N42283, N42284, N42286, N42287, N42288, N42290, N42292, N42294, N42295, N42296, N42297, N42299, N42300, N42301, N42302, N42303, N42304, N42305, N42306, N42308, N42310, N42311, N42313, N42315, N42317, N42318, N42320, N42322, N42323, N42326, N42327, N42328, N42330, N42331, N42332, N42336, N42337, N42342, N42343, N42344, N42345, N42350, N42351, N42352, N42353, N42354, N42355, N42356, N42357, N42360, N42362, N42363, N42364, N42365, N42367, N42368, N42369, N42370, N42376, N42378, N42381, N42382, N42384, N42385, N42386, N42388, N42389, N42390, N42392, N42393, N42395, N42397, N42398, N42399, N42400, N42404, N42406, N42407, N42410, N42411, N42412, N42413, N42414, N42415, N42417, N42418, N42420, N42421, N42422, N42423, N42426, N42427, N42428, N42430, N42431, N42432, N42433, N42434, N42436, N42438, N42439, N42440, N42441, N42446, N42448, N42449, N42450, N42451, N42453, N42457, N42458, N42459, N42460, N42461, N42462, N42463, N42464, N42465, N42466, N42468, N42469, N42470, N42471, N42472, N42473, N42475, N42476, N42477, N42480, N42482, N42483, N42484, N42487, N42488, N42491, N42492, N42493, N42494, N42496, N42498, N42499, N42500, N42502, N42503, N42505, N42508, N42512, N42513, N42515, N42516, N42517, N42519, N42522, N42523, N42524, N42527, N42528, N42529, N42531, N42532, N42534, N42535, N42541, N42542, N42545, N42547, N42548, N42549, N42551, N42552, N42553, N42554, N42556, N42559, N42561, N42562, N42563, N42564, N42565, N42569, N42571, N42572, N42573, N42575, N42577, N42578, N42579, N42581, N42582, N42584, N42585, N42586, N42587, N42588, N42589, N42590, N42591, N42592, N42596, N42599, N42601, N42602, N42603, N42605, N42606, N42607, N42609, N42610, N42611, N42612, N42614, N42615, N42616, N42619, N42620, N42622, N42624, N42628, N42629, N42630, N42631, N42632, N42635, N42636, N42638, N42639, N42642, N42645, N42646, N42649, N42650, N42651, N42653, N42655, N42657, N42659, N42662, N42664, N42665, N42667, N42671, N42672, N42673, N42679, N42681, N42682, N42683, N42684, N42685, N42686, N42687, N42688, N42691, N42693, N42698, N42699, N42700, N42701, N42702, N42703, N42704, N42708, N42710, N42711, N42713, N42714, N42717, N42718, N42719, N42721, N42723, N42724, N42725, N42726, N42727, N42729, N42730, N42731, N42732, N42733, N42734, N42737, N42739, N42740, N42741, N42742, N42745, N42746, N42747, N42748, N42753, N42754, N42755, N42756, N42757, N42758, N42760, N42763, N42764, N42765, N42766, N42768, N42769, N42771, N42773, N42774, N42775, N42776, N42777, N42778, N42779, N42780, N42781, N42782, N42784, N42785, N42786, N42787, N42789, N42791, N42794, N42795, N42796, N42797, N42799, N42801, N42802, N42803, N42804, N42805, N42808, N42809, N42810, N42811, N42813, N42814, N42815, N42816, N42817, N42818, N42820, N42821, N42822, N42823, N42824, N42825, N42826, N42830, N42831, N42833, N42837, N42838, N42842, N42843, N42845, N42846, N42847, N42848, N42849, N42850, N42852, N42853, N42854, N42855, N42857, N42859, N42860, N42863, N42864, N42866, N42868, N42869, N42871, N42872, N42874, N42875, N42876, N42880, N42882, N42884, N42885, N42887, N42888, N42889, N42892, N42893, N42894, N42896, N42897, N42898, N42900, N42902, N42903, N42904, N42905, N42906, N42908, N42909, N42910, N42911, N42912, N42913, N42914, N42915, N42917, N42918, N42919, N42920, N42921, N42922, N42923, N42924, N42925, N42926, N42927, N42928, N42929, N42932, N42936, N42938, N42939, N42940, N42941, N42942, N42944, N42946, N42947, N42949, N42950, N42951, N42952, N42953, N42956, N42957, N42958, N42959, N42963, N42964, N42965, N42966, N42969, N42971, N42972, N42973, N42974, N42977, N42979, N42983, N42984, N42985, N42986, N42987, N42988, N42989, N42990, N42991, N42993, N42994, N42995, N42996, N42997, N42999, N43001, N43002, N43003, N43004, N43005, N43006, N43008, N43009, N43010, N43011, N43012, N43013, N43014, N43016, N43018, N43019, N43020, N43021, N43022, N43024, N43026, N43027, N43028, N43029, N43030, N43031, N43033, N43034, N43035, N43036, N43037, N43038, N43039, N43040, N43041, N43042, N43043, N43044, N43047, N43048, N43049, N43050, N43051, N43052, N43054, N43057, N43058, N43059, N43060, N43061, N43062, N43063, N43064, N43065, N43066, N43068, N43069, N43070, N43071, N43072, N43075, N43079, N43080, N43081, N43082, N43083, N43084, N43088, N43089, N43091, N43093, N43094, N43095, N43098, N43105, N43106, N43107, N43108, N43110, N43111, N43112, N43113, N43114, N43115, N43116, N43117, N43118, N43119, N43121, N43122, N43123, N43124, N43125, N43126, N43127, N43130, N43131, N43132, N43134, N43135, N43137, N43139, N43140, N43141, N43142, N43143, N43144, N43145, N43146, N43147, N43148, N43150, N43151, N43152, N43153, N43154, N43156, N43157, N43158, N43159, N43161, N43162, N43163, N43164, N43165, N43166, N43168, N43169, N43170, N43173, N43174, N43175, N43179, N43180, N43181, N43183, N43187, N43188, N43189, N43190, N43191, N43192, N43193, N43194, N43196, N43197, N43200, N43203, N43204, N43206, N43207, N43210, N43211, N43212, N43214, N43215, N43216, N43219, N43222, N43223, N43225, N43226, N43230, N43232, N43233, N43234, N43236, N43237, N43238, N43240, N43241, N43242, N43243, N43244, N43245, N43246, N43247, N43248, N43250, N43252, N43253, N43255, N43256, N43258, N43259, N43260, N43262, N43263, N43266, N43267, N43270, N43274, N43275, N43277, N43279, N43280, N43281, N43283, N43284, N43285, N43287, N43288, N43289, N43290, N43294, N43295, N43297, N43298, N43299, N43300, N43301, N43302, N43305, N43306, N43307, N43308, N43310, N43313, N43316, N43317, N43318, N43319, N43320, N43321, N43322, N43323, N43328, N43332, N43334, N43335, N43336, N43337, N43338, N43339, N43340, N43341, N43342, N43343, N43345, N43348, N43349, N43350, N43351, N43352, N43353, N43354, N43355, N43356, N43357, N43361, N43362, N43364, N43365, N43368, N43369, N43372, N43373, N43374, N43376, N43377, N43378, N43379, N43380, N43381, N43382, N43383, N43384, N43386, N43387, N43388, N43390, N43391, N43392, N43393, N43394, N43397, N43399, N43400, N43401, N43402, N43403, N43404, N43407, N43409, N43411, N43412, N43413, N43414, N43416, N43417, N43418, N43420, N43421, N43422, N43423, N43424, N43425, N43426, N43428, N43430, N43431, N43432, N43433, N43434, N43437, N43438, N43439, N43440, N43442, N43443, N43444, N43446, N43447, N43448, N43449, N43450, N43452, N43455, N43456, N43457, N43458, N43459, N43460, N43461, N43462, N43463, N43465, N43466, N43467, N43468, N43469, N43470, N43472, N43473, N43474, N43476, N43477, N43478, N43479, N43480, N43481, N43482, N43483, N43484, N43485, N43486, N43487, N43488, N43489, N43490, N43491, N43492, N43493, N43494, N43495, N43496, N43497, N43498, N43499, N43500, N43501, N43502, N43503, N43504, N43505, N43506, N43507, N43508, N43509, N43510, N43511, N43512, N43513, N43514, N43515, N43516, N43517, N43518, N43519, N43520, N43521, N43522, N43524, N43525, N43526, N43527, N43528, N43529, N43530, N43531, N43532, N43533, N43535, N43536, N43537, N43538, N43540, N43541, N43542, N43544, N43545, N43546, N43547, N43548, N43549, N43550, N43551, N43552, N43553, N43555, N43556, N43558, N43560, N43562, N43563, N43565, N43566, N43567, N43568, N43569, N43570, N43571, N43572, N43573, N43574, N43576, N43577, N43578, N43579, N43580, N43581, N43583, N43584, N43586, N43587, N43588, N43589, N43590, N43591, N43592, N43594, N43595, N43596, N43597, N43598, N43599, N43600, N43601, N43602, N43603, N43604, N43605, N43606, N43607, N43608, N43609, N43610, N43611, N43612, N43613, N43614, N43615, N43616, N43617, N43618, N43619, N43621, N43622, N43623, N43624, N43625, N43626, N43628, N43629, N43630, N43632, N43634, N43635, N43636, N43637, N43638, N43639, N43640, N43641, N43642, N43644, N43645, N43646, N43647, N43648, N43649, N43650, N43651, N43652, N43653, N43654, N43655, N43656, N43657, N43658, N43659, N43660, N43661, N43662, N43663, N43664, N43665, N43666, N43667, N43668, N43669, N43670, N43671, N43672, N43673, N43674, N43676, N43677, N43678, N43679, N43680, N43681, N43682, N43683, N43684, N43685, N43686, N43687, N43688, N43689, N43691, N43692, N43693, N43694, N43695, N43696, N43697, N43698, N43699, N43700, N43701, N43702, N43704, N43705, N43706, N43707, N43708, N43709, N43710, N43711, N43712, N43713, N43714, N43715, N43716, N43717, N43718, N43719, N43720, N43721, N43722, N43723, N43724, N43725, N43726, N43727, N43728, N43730, N43731, N43732, N43733, N43734, N43735, N43736, N43737, N43738, N43739, N43740, N43741, N43742, N43743, N43744, N43745, N43746, N43748, N43749, N43750, N43751, N43752, N43753, N43754, N43755, N43756, N43757, N43758, N43759, N43761, N43763, N43765, N43766, N43767, N43768, N43769, N43772, N43773, N43774, N43775, N43777, N43778, N43779, N43780, N43781, N43782, N43783, N43784, N43785, N43786, N43787, N43788, N43789, N43790, N43791, N43792, N43793, N43794, N43795, N43797, N43798, N43799, N43800, N43801, N43802, N43804, N43805, N43806, N43807, N43808, N43809, N43810, N43811, N43812, N43813, N43814, N43815, N43816, N43817, N43818, N43819, N43820, N43821, N43822, N43823, N43824, N43825, N43826, N43827, N43828, N43829, N43830, N43831, N43832, N43833, N43834, N43835, N43836, N43837, N43838, N43839, N43840, N43841, N43842, N43843, N43845, N43846, N43847, N43848, N43849, N43850, N43851, N43852, N43853, N43854, N43855, N43856, N43857, N43859, N43860, N43861, N43862, N43863, N43864, N43865, N43866, N43867, N43868, N43869, N43870, N43871, N43872, N43873, N43874, N43875, N43876, N43877, N43879, N43880, N43881, N43882, N43883, N43884, N43885, N43886, N43887, N43888, N43889, N43891, N43892, N43893, N43894, N43895, N43896, N43897, N43898, N43900, N43901, N43902, N43903, N43904, N43905, N43906, N43907, N43908, N43909, N43910, N43911, N43912, N43913, N43914, N43915, N43916, N43917, N43918, N43919, N43921, N43922, N43923, N43924, N43925, N43926, N43927, N43928, N43929, N43930, N43931, N43932, N43934, N43935, N43936, N43937, N43938, N43939, N43942, N43943, N43944, N43945, N43946, N43947, N43948, N43949, N43950, N43951, N43952, N43953, N43955, N43956, N43957, N43958, N43959, N43960, N43961, N43962, N43964, N43965, N43966, N43967, N43968, N43969, N43970, N43971, N43972, N43973, N43974, N43975, N43976, N43977, N43978, N43979, N43980, N43981, N43982, N43983, N43984, N43985, N43986, N43987, N43988, N43989, N43990, N43991, N43992, N43994, N43995, N43996, N43997, N43999, N44000, N44001, N44002, N44003, N44004, N44005, N44007, N44008, N44009, N44010, N44011, N44012, N44013, N44014, N44015, N44016, N44017, N44018, N44019, N44020, N44021, N44022, N44023, N44024, N44025, N44026, N44027, N44028, N44029, N44030, N44031, N44032, N44033, N44034, N44035, N44036, N44037, N44038, N44039, N44040, N44041, N44042, N44043, N44044, N44045, N44046, N44047, N44048, N44049, N44050, N44051, N44052, N44053, N44055, N44056, N44057, N44058, N44059, N44060, N44061, N44062, N44063, N44064, N44065, N44066, N44067, N44069, N44070, N44071, N44072, N44073, N44074, N44075, N44076, N44077, N44078, N44079, N44080, N44081, N44082, N44083, N44084, N44085, N44086, N44087, N44088, N44089, N44090, N44091, N44092, N44093, N44094, N44095, N44097, N44098, N44099, N44100, N44101, N44102, N44103, N44105, N44106, N44107, N44108, N44109, N44110, N44111, N44112, N44113, N44114, N44115, N44116, N44117, N44118, N44119, N44121, N44122, N44123, N44124, N44125, N44126, N44127, N44128, N44129, N44130, N44131, N44132, N44133, N44135, N44136, N44137, N44139, N44141, N44142, N44143, N44144, N44145, N44146, N44147, N44148, N44149, N44150, N44151, N44152, N44153, N44154, N44155, N44156, N44158, N44159, N44160, N44161, N44162, N44163, N44164, N44165, N44166, N44167, N44168, N44169, N44171, N44172, N44174, N44175, N44177, N44178, N44181, N44182, N44183, N44184, N44185, N44186, N44187, N44188, N44189, N44190, N44191, N44192, N44193, N44194, N44195, N44196, N44197, N44198, N44199, N44200, N44201, N44202, N44203, N44204, N44205, N44206, N44207, N44208, N44209, N44210, N44212, N44213, N44215, N44216, N44217, N44218, N44219, N44220, N44221, N44222, N44224, N44225, N44226, N44227, N44229, N44230, N44232, N44233, N44234, N44235, N44236, N44237, N44238, N44239, N44240, N44241, N44242, N44243, N44244, N44246, N44248, N44249, N44250, N44251, N44252, N44254, N44255, N44256, N44257, N44258, N44259, N44261, N44262, N44263, N44264, N44265, N44266, N44267, N44268, N44269, N44271, N44272, N44273, N44274, N44275, N44276, N44277, N44278, N44279, N44281, N44282, N44283, N44284, N44285, N44286, N44288, N44289, N44290, N44291, N44292, N44293, N44294, N44295, N44296, N44297, N44298, N44299, N44300, N44301, N44302, N44303, N44304, N44305, N44306, N44307, N44308, N44309, N44310, N44311, N44312, N44313, N44314, N44316, N44317, N44318, N44319, N44320, N44321, N44322, N44323, N44324, N44325, N44326, N44327, N44328, N44329, N44330, N44331, N44332, N44333, N44334, N44335, N44338, N44339, N44341, N44342, N44343, N44345, N44346, N44347, N44348, N44349, N44350, N44352, N44353, N44354, N44355, N44356, N44357, N44359, N44360, N44363, N44364, N44365, N44366, N44367, N44368, N44369, N44370, N44371, N44372, N44373, N44375, N44376, N44377, N44378, N44379, N44380, N44381, N44384, N44385, N44386, N44387, N44388, N44389, N44390, N44391, N44392, N44393, N44394, N44395, N44396, N44397, N44399, N44400, N44401, N44402, N44403, N44404, N44405, N44406, N44407, N44408, N44409, N44410, N44411, N44412, N44413, N44414, N44415, N44416, N44417, N44418, N44419, N44420, N44421, N44422, N44423, N44424, N44425, N44426, N44427, N44428, N44429, N44430, N44431, N44432, N44433, N44434, N44435, N44436, N44437, N44438, N44440, N44441, N44442, N44443, N44444, N44445, N44446, N44447, N44448, N44450, N44451, N44452, N44453, N44456, N44457, N44458, N44459, N44461, N44462, N44463, N44464, N44465, N44466, N44467, N44469, N44470, N44471, N44472, N44473, N44474, N44475, N44476, N44478, N44479, N44480, N44481, N44482, N44483, N44484, N44486, N44488, N44489, N44491, N44492, N44493, N44494, N44495, N44496, N44497, N44498, N44499, N44500, N44502, N44503, N44504, N44505, N44506, N44507, N44508, N44509, N44510, N44511, N44512, N44513, N44514, N44515, N44516, N44517, N44518, N44519, N44520, N44521, N44522, N44523, N44525, N44526, N44527, N44528, N44529, N44530, N44531, N44532, N44533, N44534, N44536, N44537, N44538, N44539, N44540, N44541, N44543, N44544, N44545, N44547, N44548, N44549, N44550, N44551, N44552, N44553, N44554, N44555, N44556, N44557, N44558, N44559, N44560, N44561, N44562, N44563, N44564, N44566, N44567, N44568, N44569, N44570, N44572, N44573, N44574, N44575, N44576, N44577, N44578, N44579, N44580, N44581, N44582, N44583, N44585, N44586, N44587, N44588, N44589, N44590, N44592, N44593, N44594, N44595, N44596, N44597, N44598, N44599, N44600, N44601, N44602, N44604, N44605, N44606, N44607, N44608, N44609, N44610, N44611, N44612, N44613, N44614, N44615, N44616, N44617, N44618, N44619, N44620, N44621, N44622, N44625, N44626, N44627, N44628, N44629, N44630, N44631, N44632, N44633, N44634, N44635, N44636, N44637, N44638, N44639, N44641, N44643, N44644, N44645, N44646, N44647, N44648, N44649, N44650, N44651, N44652, N44653, N44654, N44655, N44656, N44657, N44658, N44659, N44660, N44661, N44662, N44664, N44666, N44667, N44668, N44669, N44670, N44671, N44672, N44673, N44674, N44675, N44676, N44677, N44678, N44679, N44680, N44681, N44682, N44683, N44684, N44685, N44686, N44687, N44688, N44689, N44690, N44691, N44692, N44693, N44694, N44695, N44696, N44698, N44699, N44700, N44701, N44702, N44704, N44705, N44706, N44707, N44709, N44711, N44712, N44713, N44714, N44715, N44716, N44717, N44718, N44719, N44722, N44723, N44724, N44725, N44726, N44728, N44729, N44730, N44732, N44733, N44734, N44735, N44736, N44737, N44738, N44739, N44740, N44741, N44742, N44743, N44744, N44745, N44746, N44748, N44749, N44750, N44751, N44752, N44753, N44754, N44755, N44756, N44757, N44758, N44759, N44760, N44761, N44762, N44763, N44764, N44768, N44769, N44770, N44771, N44772, N44773, N44774, N44775, N44776, N44777, N44778, N44779, N44780, N44781, N44782, N44783, N44784, N44785, N44786, N44787, N44788, N44789, N44791, N44792, N44793, N44795, N44797, N44798, N44799, N44801, N44802, N44803, N44804, N44805, N44806, N44807, N44808, N44809, N44810, N44811, N44812, N44813, N44814, N44815, N44816, N44817, N44818, N44819, N44820, N44821, N44823, N44824, N44825, N44826, N44827, N44828, N44829, N44830, N44831, N44832, N44833, N44835, N44836, N44837, N44838, N44839, N44840, N44841, N44842, N44843, N44844, N44845, N44846, N44847, N44848, N44850, N44851, N44852, N44853, N44854, N44855, N44856, N44857, N44858, N44859, N44860, N44861, N44862, N44863, N44864, N44865, N44866, N44867, N44868, N44869, N44870, N44871, N44872, N44873, N44874, N44875, N44876, N44877, N44878, N44879, N44880, N44881, N44882, N44883, N44884, N44885, N44886, N44888, N44889, N44890, N44891, N44893, N44894, N44896, N44897, N44898, N44899, N44900, N44901, N44902, N44903, N44904, N44905, N44906, N44907, N44908, N44909, N44910, N44911, N44912, N44913, N44914, N44915, N44916, N44917, N44918, N44919, N44920, N44921, N44922, N44923, N44924, N44925, N44926, N44927, N44928, N44929, N44930, N44931, N44932, N44933, N44934, N44935, N44936, N44938, N44939, N44940, N44941, N44942, N44943, N44945, N44946, N44947, N44948, N44949, N44950, N44952, N44953, N44954, N44955, N44956, N44957, N44958, N44959, N44960, N44961, N44962, N44963, N44964, N44965, N44966, N44968, N44969, N44971, N44972, N44973, N44974, N44976, N44977, N44978, N44979, N44980, N44981, N44982, N44983, N44984, N44985, N44986, N44989, N44990, N44991, N44992, N44993, N44994, N44995, N44996, N44997, N44998, N44999, N45000, N45001, N45002, N45003, N45004, N45005, N45006, N45007, N45008, N45009, N45010, N45011, N45012, N45013, N45014, N45015, N45016, N45017, N45018, N45020, N45021, N45022, N45023, N45024, N45025, N45026, N45027, N45028, N45029, N45030, N45031, N45032, N45033, N45034, N45036, N45037, N45038, N45039, N45040, N45041, N45042, N45043, N45044, N45045, N45046, N45047, N45048, N45050, N45051, N45052, N45053, N45054, N45055, N45056, N45057, N45058, N45059, N45060, N45061, N45063, N45064, N45065, N45066, N45067, N45068, N45069, N45070, N45071, N45072, N45073, N45074, N45075, N45076, N45078, N45079, N45080, N45081, N45082, N45084, N45085, N45086, N45087, N45088, N45089, N45090, N45091, N45092, N45093, N45094, N45095, N45096, N45097, N45098, N45099, N45100, N45101, N45102, N45103, N45105, N45106, N45107, N45108, N45109, N45110, N45111, N45113, N45114, N45115, N45116, N45117, N45118, N45119, N45120, N45121, N45122, N45123, N45124, N45125, N45127, N45128, N45129, N45130, N45131, N45132, N45133, N45135, N45136, N45138, N45139, N45142, N45143, N45144, N45145, N45146, N45147, N45148, N45149, N45150, N45151, N45153, N45154, N45155, N45157, N45158, N45159, N45160, N45161, N45162, N45163, N45164, N45165, N45166, N45167, N45168, N45169, N45170, N45171, N45172, N45173, N45174, N45175, N45176, N45178, N45179, N45180, N45181, N45182, N45183, N45185, N45186, N45187, N45188, N45189, N45190, N45191, N45192, N45193, N45194, N45195, N45196, N45197, N45198, N45199, N45200, N45201, N45202, N45203, N45205, N45206, N45208, N45209, N45210, N45212, N45213, N45214, N45215, N45216, N45217, N45219, N45220, N45221, N45222, N45223, N45224, N45225, N45227, N45228, N45229, N45230, N45231, N45232, N45233, N45234, N45235, N45236, N45237, N45238, N45242, N45243, N45244, N45245, N45246, N45247, N45248, N45249, N45250, N45251, N45252, N45253, N45254, N45255, N45256, N45257, N45258, N45259, N45260, N45261, N45262, N45263, N45267, N45269, N45270, N45271, N45272, N45273, N45274, N45275, N45276, N45277, N45278, N45279, N45280, N45281, N45282, N45283, N45284, N45285, N45286, N45287, N45288, N45289, N45290, N45291, N45292, N45293, N45294, N45295, N45296, N45297, N45298, N45299, N45300, N45301, N45303, N45304, N45305, N45307, N45308, N45309, N45310, N45311, N45312, N45313, N45314, N45316, N45317, N45318, N45319, N45320, N45321, N45322, N45323, N45324, N45325, N45326, N45327, N45328, N45329, N45330, N45331, N45332, N45333, N45335, N45336, N45337, N45338, N45339, N45340, N45341, N45342, N45343, N45344, N45345, N45346, N45347, N45348, N45349, N45352, N45353, N45354, N45355, N45356, N45357, N45358, N45359, N45360, N45361, N45362, N45363, N45364, N45365, N45366, N45367, N45369, N45370, N45372, N45373, N45374, N45375, N45376, N45377, N45378, N45379, N45380, N45381, N45382, N45383, N45384, N45385, N45386, N45387, N45388, N45389, N45390, N45391, N45393, N45394, N45395, N45396, N45397, N45398, N45399, N45402, N45403, N45405, N45406, N45407, N45408, N45409, N45410, N45411, N45412, N45413, N45414, N45415, N45416, N45417, N45418, N45419, N45420, N45421, N45422, N45423, N45424, N45425, N45426, N45427, N45429, N45430, N45431, N45433, N45434, N45435, N45436, N45438, N45439, N45440, N45441, N45442, N45443, N45444, N45445, N45447, N45448, N45449, N45450, N45451, N45452, N45458, N45459, N45460, N45461, N45462, N45464, N45465, N45466, N45467, N45468, N45469, N45471, N45472, N45473, N45474, N45475, N45476, N45477, N45478, N45479, N45480, N45481, N45483, N45484, N45485, N45486, N45487, N45488, N45489, N45490, N45491, N45492, N45493, N45494, N45495, N45496, N45497, N45498, N45499, N45500, N45501, N45502, N45503, N45504, N45505, N45506, N45507, N45508, N45509, N45511, N45513, N45514, N45515, N45516, N45517, N45518, N45519, N45520, N45521, N45522, N45523, N45524, N45525, N45526, N45527, N45530, N45531, N45532, N45533, N45535, N45536, N45537, N45538, N45539, N45540, N45541, N45542, N45543, N45544, N45545, N45547, N45548, N45549, N45550, N45551, N45552, N45553, N45554, N45555, N45556, N45557, N45558, N45559, N45561, N45562, N45563, N45564, N45566, N45567, N45568, N45569, N45570, N45571, N45572, N45573, N45574, N45575, N45576, N45577, N45578, N45579, N45580, N45581, N45584, N45585, N45586, N45587, N45588, N45589, N45590, N45592, N45593, N45595, N45597, N45599, N45600, N45601, N45602, N45603, N45605, N45606, N45607, N45608, N45609, N45610, N45611, N45612, N45613, N45614, N45615, N45616, N45617, N45618, N45619, N45620, N45621, N45622, N45623, N45625, N45627, N45628, N45629, N45630, N45631, N45633, N45634, N45635, N45636, N45637, N45638, N45639, N45640, N45641, N45642, N45643, N45646, N45647, N45648, N45649, N45650, N45652, N45653, N45654, N45655, N45656, N45657, N45658, N45659, N45660, N45661, N45662, N45663, N45664, N45665, N45666, N45667, N45669, N45671, N45673, N45674, N45676, N45677, N45678, N45679, N45680, N45681, N45682, N45683, N45685, N45686, N45687, N45688, N45689, N45690, N45691, N45692, N45693, N45694, N45695, N45696, N45697, N45698, N45699, N45701, N45702, N45703, N45705, N45706, N45707, N45708, N45709, N45710, N45711, N45712, N45713, N45714, N45716, N45717, N45718, N45719, N45720, N45721, N45722, N45723, N45724, N45725, N45726, N45727, N45728, N45729, N45730, N45732, N45733, N45735, N45736, N45737, N45739, N45740, N45741, N45742, N45743, N45744, N45745, N45746, N45747, N45748, N45749, N45750, N45751, N45752, N45753, N45754, N45756, N45757, N45758, N45759, N45760, N45761, N45762, N45763, N45764, N45765, N45766, N45768, N45769, N45770, N45771, N45772, N45773, N45774, N45775, N45776, N45778, N45779, N45780, N45782, N45783, N45784, N45786, N45787, N45789, N45790, N45791, N45792, N45793, N45795, N45796, N45797, N45798, N45799, N45800, N45801, N45802, N45803, N45804, N45805, N45806, N45807, N45808, N45809, N45810, N45811, N45812, N45813, N45814, N45815, N45816, N45817, N45818, N45819, N45820, N45821, N45822, N45823, N45824, N45825, N45826, N45827, N45828, N45829, N45830, N45831, N45833, N45834, N45835, N45836, N45837, N45838, N45839, N45840, N45841, N45842, N45843, N45844, N45845, N45846, N45847, N45848, N45849, N45850, N45851, N45852, N45853, N45854, N45855, N45856, N45857, N45858, N45859, N45860, N45861, N45862, N45863, N45865, N45866, N45867, N45868, N45869, N45870, N45871, N45872, N45873, N45874, N45875, N45876, N45877, N45878, N45879, N45880, N45881, N45882, N45883, N45884, N45885, N45886, N45887, N45888, N45889, N45890, N45891, N45892, N45893, N45894, N45895, N45896, N45897, N45898, N45899, N45901, N45902, N45903, N45904, N45905, N45906, N45907, N45908, N45909, N45910, N45911, N45912, N45913, N45914, N45915, N45916, N45917, N45918, N45919, N45920, N45921, N45922, N45923, N45924, N45925, N45926, N45927, N45928, N45929, N45930, N45931, N45932, N45933, N45934, N45935, N45936, N45938, N45939, N45940, N45941, N45942, N45944, N45945, N45946, N45947, N45948, N45949, N45950, N45951, N45952, N45953, N45954, N45955, N45956, N45957, N45958, N45960, N45961, N45962, N45963, N45964, N45965, N45966, N45967, N45968, N45969, N45971, N45972, N45973, N45974, N45975, N45976, N45979, N45980, N45981, N45983, N45984, N45985, N45986, N45987, N45988, N45989, N45990, N45991, N45992, N45993, N45994, N45995, N45996, N45997, N45999, N46000, N46002, N46003, N46004, N46005, N46006, N46007, N46008, N46011, N46012, N46013, N46014, N46015, N46016, N46017, N46018, N46019, N46020, N46021, N46022, N46023, N46024, N46025, N46026, N46027, N46028, N46029, N46030, N46031, N46032, N46034, N46035, N46036, N46037, N46038, N46039, N46040, N46041, N46042, N46043, N46044, N46045, N46047, N46048, N46049, N46051, N46052, N46053, N46054, N46056, N46057, N46058, N46059, N46060, N46061, N46063, N46064, N46065, N46066, N46067, N46068, N46069, N46070, N46071, N46072, N46073, N46074, N46075, N46077, N46078, N46079, N46080, N46081, N46082, N46085, N46086, N46087, N46089, N46090, N46091, N46092, N46093, N46094, N46095, N46096, N46097, N46098, N46099, N46100, N46101, N46102, N46103, N46104, N46105, N46106, N46107, N46108, N46109, N46110, N46111, N46112, N46113, N46114, N46115, N46116, N46117, N46118, N46121, N46122, N46123, N46124, N46125, N46126, N46127, N46128, N46129, N46131, N46132, N46133, N46134, N46135, N46136, N46137, N46139, N46140, N46141, N46142, N46143, N46144, N46145, N46146, N46147, N46148, N46149, N46150, N46151, N46152, N46153, N46154, N46155, N46156, N46157, N46158, N46159, N46160, N46161, N46162, N46163, N46164, N46166, N46167, N46168, N46169, N46170, N46171, N46172, N46173, N46174, N46175, N46176, N46177, N46178, N46179, N46180, N46181, N46182, N46183, N46184, N46185, N46186, N46187, N46188, N46190, N46191, N46192, N46193, N46194, N46195, N46196, N46197, N46198, N46200, N46201, N46202, N46203, N46204, N46205, N46206, N46207, N46208, N46209, N46210, N46211, N46212, N46213, N46214, N46215, N46216, N46217, N46218, N46219, N46220, N46221, N46222, N46223, N46226, N46227, N46228, N46229, N46230, N46231, N46232, N46233, N46234, N46235, N46236, N46237, N46238, N46239, N46241, N46242, N46243, N46244, N46245, N46246, N46247, N46248, N46249, N46251, N46252, N46253, N46254, N46255, N46256, N46257, N46258, N46260, N46261, N46262, N46263, N46264, N46265, N46267, N46268, N46269, N46270, N46271, N46272, N46273, N46274, N46275, N46276, N46277, N46278, N46280, N46281, N46282, N46283, N46284, N46285, N46286, N46288, N46289, N46290, N46291, N46292, N46293, N46295, N46296, N46297, N46298, N46299, N46302, N46303, N46304, N46305, N46306, N46307, N46309, N46310, N46311, N46312, N46314, N46315, N46316, N46317, N46318, N46319, N46320, N46321, N46322, N46323, N46324, N46325, N46326, N46327, N46328, N46329, N46330, N46331, N46332, N46333, N46336, N46337, N46338, N46339, N46340, N46341, N46342, N46343, N46344, N46345, N46346, N46347, N46348, N46349, N46350, N46351, N46352, N46353, N46354, N46355, N46356, N46357, N46358, N46359, N46360, N46361, N46362, N46365, N46366, N46367, N46368, N46369, N46370, N46371, N46372, N46373, N46374, N46375, N46376, N46377, N46378, N46379, N46380, N46381, N46382, N46384, N46385, N46387, N46388, N46389, N46391, N46393, N46394, N46395, N46396, N46397, N46398, N46399, N46400, N46401, N46402, N46403, N46404, N46405, N46406, N46407, N46408, N46409, N46410, N46411, N46412, N46413, N46414, N46415, N46416, N46417, N46419, N46420, N46421, N46422, N46423, N46424, N46425, N46426, N46428, N46429, N46430, N46431, N46432, N46433, N46434, N46435, N46436, N46437, N46438, N46439, N46440, N46441, N46442, N46443, N46444, N46445, N46446, N46447, N46448, N46449, N46450, N46451, N46452, N46453, N46454, N46455, N46456, N46457, N46459, N46460, N46461, N46462, N46463, N46464, N46465, N46466, N46467, N46468, N46469, N46470, N46471, N46472, N46473, N46474, N46475, N46476, N46477, N46478, N46479, N46480, N46481, N46483, N46484, N46485, N46486, N46487, N46489, N46490, N46491, N46492, N46493, N46494, N46495, N46496, N46497, N46498, N46499, N46500, N46501, N46503, N46505, N46506, N46507, N46508, N46509, N46510, N46511, N46512, N46513, N46514, N46515, N46517, N46518, N46519, N46520, N46521, N46523, N46524, N46525, N46526, N46527, N46528, N46529, N46530, N46531, N46532, N46533, N46534, N46536, N46537, N46538, N46539, N46540, N46541, N46542, N46543, N46544, N46545, N46546, N46547, N46548, N46549, N46550, N46551, N46552, N46553, N46554, N46555, N46556, N46557, N46558, N46559, N46560, N46561, N46562, N46563, N46564, N46565, N46566, N46567, N46568, N46569, N46570, N46571, N46572, N46573, N46574, N46575, N46576, N46577, N46578, N46579, N46580, N46581, N46582, N46583, N46584, N46585, N46586, N46587, N46588, N46589, N46590, N46591, N46592, N46593, N46594, N46596, N46597, N46598, N46599, N46601, N46602, N46603, N46604, N46605, N46606, N46608, N46609, N46610, N46611, N46612, N46613, N46614, N46615, N46616, N46617, N46618, N46619, N46620, N46621, N46622, N46623, N46624, N46625, N46626, N46627, N46628, N46629, N46631, N46632, N46633, N46634, N46635, N46636, N46637, N46638, N46639, N46640, N46641, N46642, N46643, N46644, N46645, N46646, N46647, N46648, N46649, N46650, N46651, N46653, N46654, N46655, N46656, N46657, N46658, N46659, N46660, N46661, N46662, N46664, N46665, N46666, N46667, N46668, N46669, N46671, N46672, N46673, N46674, N46675, N46676, N46677, N46678, N46679, N46680, N46681, N46682, N46683, N46684, N46685, N46686, N46687, N46688, N46689, N46690, N46691, N46692, N46693, N46694, N46695, N46696, N46697, N46699, N46700, N46701, N46702, N46703, N46704, N46705, N46707, N46708, N46709, N46710, N46712, N46713, N46714, N46715, N46716, N46717, N46718, N46719, N46720, N46721, N46722, N46723, N46725, N46726, N46727, N46728, N46729, N46730, N46731, N46732, N46733, N46734, N46735, N46736, N46737, N46738, N46740, N46741, N46742, N46743, N46744, N46745, N46746, N46747, N46748, N46749, N46750, N46751, N46752, N46753, N46754, N46756, N46757, N46758, N46759, N46760, N46761, N46762, N46763, N46764, N46765, N46766, N46767, N46768, N46769, N46772, N46773, N46774, N46775, N46776, N46777, N46778, N46779, N46780, N46781, N46782, N46783, N46784, N46785, N46786, N46787, N46788, N46790, N46791, N46792, N46793, N46794, N46795, N46796, N46797, N46798, N46799, N46800, N46801, N46802, N46803, N46804, N46805, N46806, N46807, N46808, N46809, N46810, N46812, N46813, N46814, N46815, N46816, N46817, N46818, N46819, N46820, N46821, N46822, N46823, N46824, N46825, N46826, N46827, N46828, N46829, N46830, N46832, N46833, N46834, N46835, N46836, N46837, N46838, N46839, N46840, N46841, N46843, N46844, N46845, N46846, N46847, N46848, N46850, N46851, N46852, N46853, N46854, N46855, N46856, N46857, N46859, N46860, N46862, N46863, N46864, N46865, N46866, N46867, N46868, N46869, N46870, N46871, N46872, N46873, N46874, N46875, N46876, N46877, N46878, N46879, N46880, N46881, N46882, N46883, N46884, N46885, N46886, N46887, N46888, N46889, N46890, N46891, N46892, N46893, N46894, N46895, N46896, N46897, N46898, N46899, N46900, N46902, N46903, N46904, N46905, N46906, N46907, N46908, N46909, N46910, N46911, N46912, N46913, N46914, N46915, N46916, N46917, N46918, N46919, N46920, N46921, N46922, N46923, N46924, N46925, N46926, N46928, N46929, N46931, N46932, N46933, N46934, N46935, N46936, N46937, N46939, N46940, N46941, N46942, N46945, N46946, N46947, N46948, N46949, N46950, N46951, N46952, N46953, N46954, N46955, N46956, N46957, N46958, N46959, N46960, N46961, N46962, N46963, N46964, N46965, N46966, N46967, N46968, N46969, N46970, N46971, N46972, N46973, N46975, N46976, N46977, N46978, N46979, N46980, N46981, N46982, N46983, N46984, N46985, N46987, N46988, N46989, N46990, N46991, N46992, N46993, N46994, N46995, N46997, N46998, N46999, N47001, N47002, N47003, N47004, N47005, N47006, N47007, N47008, N47009, N47010, N47011, N47012, N47013, N47014, N47015, N47016, N47017, N47018, N47019, N47020, N47021, N47023, N47024, N47025, N47026, N47027, N47028, N47029, N47030, N47031, N47032, N47034, N47035, N47036, N47037, N47038, N47039, N47040, N47041, N47042, N47043, N47044, N47045, N47046, N47047, N47048, N47049, N47050, N47051, N47052, N47053, N47054, N47055, N47056, N47058, N47059, N47060, N47061, N47062, N47063, N47064, N47065, N47066, N47067, N47068, N47069, N47070, N47071, N47072, N47073, N47074, N47075, N47076, N47077, N47078, N47079, N47080, N47081, N47082, N47083, N47084, N47086, N47087, N47088, N47089, N47090, N47091, N47092, N47093, N47094, N47095, N47096, N47097, N47098, N47099, N47100, N47101, N47102, N47103, N47104, N47105, N47106, N47107, N47108, N47109, N47110, N47111, N47112, N47113, N47115, N47116, N47118, N47119, N47120, N47121, N47122, N47123, N47124, N47125, N47127, N47128, N47129, N47130, N47131, N47133, N47134, N47135, N47136, N47137, N47138, N47139, N47141, N47142, N47143, N47145, N47146, N47147, N47148, N47149, N47150, N47151, N47152, N47153, N47155, N47156, N47157, N47158, N47159, N47160, N47161, N47162, N47163, N47164, N47165, N47166, N47167, N47168, N47170, N47171, N47172, N47173, N47174, N47175, N47176, N47177, N47178, N47179, N47180, N47181, N47182, N47184, N47185, N47186, N47187, N47188, N47189, N47190, N47191, N47192, N47193, N47196, N47197, N47198, N47199, N47200, N47201, N47202, N47203, N47204, N47205, N47206, N47207, N47208, N47209, N47210, N47211, N47212, N47213, N47214, N47215, N47216, N47217, N47219, N47220, N47221, N47222, N47223, N47224, N47225, N47226, N47227, N47228, N47229, N47230, N47231, N47232, N47234, N47235, N47236, N47237, N47238, N47239, N47240, N47241, N47242, N47243, N47244, N47246, N47247, N47248, N47249, N47250, N47251, N47252, N47253, N47254, N47255, N47256, N47257, N47258, N47259, N47260, N47261, N47262, N47263, N47264, N47266, N47267, N47268, N47269, N47270, N47271, N47272, N47273, N47274, N47275, N47276, N47277, N47278, N47279, N47280, N47281, N47282, N47283, N47284, N47285, N47286, N47287, N47288, N47289, N47290, N47291, N47292, N47293, N47294, N47295, N47296, N47297, N47298, N47299, N47300, N47301, N47302, N47303, N47304, N47305, N47306, N47307, N47308, N47309, N47310, N47311, N47312, N47313, N47314, N47315, N47316, N47317, N47318, N47319, N47320, N47321, N47322, N47323, N47324, N47325, N47326, N47327, N47328, N47329, N47330, N47331, N47332, N47335, N47336, N47337, N47338, N47339, N47340, N47341, N47342, N47343, N47344, N47345, N47346, N47347, N47348, N47349, N47350, N47351, N47352, N47353, N47354, N47355, N47356, N47357, N47358, N47359, N47360, N47361, N47362, N47363, N47364, N47365, N47366, N47367, N47368, N47369, N47370, N47371, N47372, N47373, N47374, N47376, N47378, N47379, N47380, N47381, N47382, N47383, N47384, N47385, N47386, N47387, N47388, N47389, N47390, N47391, N47392, N47393, N47394, N47395, N47396, N47397, N47398, N47399, N47400, N47401, N47402, N47403, N47404, N47405, N47406, N47407, N47408, N47409, N47410, N47411, N47412, N47413, N47414, N47415, N47416, N47417, N47418, N47420, N47421, N47422, N47423, N47424, N47425, N47426, N47427, N47428, N47429, N47430, N47432, N47433, N47434, N47435, N47436, N47437, N47438, N47439, N47440, N47441, N47442, N47443, N47444, N47445, N47446, N47447, N47448, N47449, N47450, N47452, N47453, N47455, N47456, N47457, N47458, N47459, N47460, N47461, N47462, N47463, N47464, N47465, N47466, N47467, N47468, N47469, N47470, N47472, N47473, N47474, N47476, N47477, N47478, N47479, N47480, N47481, N47482, N47483, N47484, N47485, N47486, N47487, N47488, N47489, N47490, N47491, N47492, N47493, N47494, N47496, N47497, N47498, N47500, N47501, N47502, N47503, N47504, N47505, N47506, N47507, N47508, N47510, N47511, N47512, N47513, N47515, N47517, N47518, N47519, N47520, N47521, N47522, N47523, N47524, N47525, N47526, N47527, N47528, N47529, N47530, N47531, N47532, N47533, N47534, N47536, N47537, N47538, N47539, N47540, N47541, N47542, N47543, N47544, N47545, N47547, N47548, N47549, N47550, N47551, N47552, N47553, N47554, N47555, N47556, N47557, N47558, N47559, N47560, N47561, N47562, N47563, N47564, N47565, N47566, N47567, N47568, N47569, N47570, N47571, N47572, N47573, N47574, N47575, N47576, N47577, N47578, N47579, N47580, N47581, N47582, N47583, N47584, N47585, N47586, N47587, N47588, N47589, N47590, N47591, N47592, N47593, N47594, N47595, N47596, N47597, N47598, N47599, N47600, N47601, N47602, N47603, N47604, N47605, N47606, N47607, N47608, N47609, N47610, N47612, N47613, N47614, N47615, N47616, N47617, N47618, N47619, N47620, N47622, N47623, N47624, N47625, N47626, N47627, N47628, N47630, N47631, N47632, N47633, N47634, N47636, N47639, N47641, N47642, N47643, N47644, N47646, N47647, N47648, N47649, N47650, N47651, N47652, N47653, N47654, N47655, N47656, N47657, N47658, N47659, N47660, N47662, N47664, N47665, N47666, N47667, N47668, N47670, N47671, N47672, N47674, N47675, N47676, N47677, N47678, N47679, N47680, N47681, N47682, N47683, N47684, N47685, N47686, N47687, N47688, N47689, N47690, N47691, N47692, N47693, N47694, N47695, N47696, N47697, N47698, N47699, N47700, N47701, N47702, N47703, N47704, N47705, N47706, N47707, N47708, N47709, N47710, N47711, N47712, N47713, N47714, N47716, N47718, N47719, N47720, N47721, N47722, N47723, N47724, N47725, N47726, N47728, N47729, N47730, N47731, N47732, N47733, N47734, N47735, N47736, N47737, N47738, N47739, N47741, N47742, N47743, N47744, N47745, N47746, N47747, N47748, N47749, N47750, N47751, N47753, N47754, N47755, N47756, N47757, N47759, N47760, N47761, N47762, N47763, N47764, N47765, N47766, N47767, N47768, N47769, N47770, N47772, N47773, N47774, N47775, N47776, N47777, N47778, N47779, N47780, N47781, N47782, N47783, N47784, N47785, N47786, N47787, N47788, N47789, N47790, N47791, N47792, N47793, N47794, N47795, N47796, N47797, N47798, N47799, N47800, N47801, N47802, N47803, N47804, N47805, N47806, N47807, N47808, N47810, N47811, N47812, N47813, N47814, N47815, N47816, N47817, N47818, N47819, N47820, N47821, N47822, N47823, N47824, N47825, N47826, N47827, N47828, N47829, N47830, N47831, N47832, N47833, N47834, N47835, N47836, N47837, N47839, N47840, N47841, N47842, N47843, N47845, N47846, N47847, N47848, N47849, N47850, N47851, N47852, N47853, N47854, N47855, N47856, N47857, N47858, N47859, N47860, N47861, N47862, N47863, N47864, N47865, N47866, N47867, N47868, N47869, N47870, N47871, N47872, N47874, N47875, N47876, N47877, N47878, N47880, N47881, N47882, N47883, N47884, N47885, N47886, N47887, N47888, N47889, N47890, N47891, N47892, N47893, N47894, N47895, N47896, N47897, N47898, N47899, N47900, N47901, N47903, N47904, N47905, N47906, N47907, N47908, N47909, N47910, N47911, N47912, N47913, N47914, N47915, N47916, N47917, N47918, N47919, N47920, N47922, N47923, N47925, N47926, N47927, N47928, N47929, N47930, N47931, N47932, N47933, N47934, N47935, N47936, N47937, N47938, N47939, N47940, N47941, N47942, N47943, N47944, N47945, N47946, N47948, N47949, N47950, N47951, N47952, N47953, N47954, N47955, N47957, N47958, N47959, N47960, N47961, N47962, N47963, N47964, N47965, N47966, N47967, N47968, N47969, N47970, N47971, N47972, N47973, N47974, N47975, N47976, N47977, N47978, N47979, N47980, N47981, N47982, N47983, N47984, N47985, N47986, N47987, N47988, N47989, N47990, N47991, N47992, N47993, N47994, N47995, N47996, N47997, N47998, N47999, N48000, N48001, N48002, N48003, N48004, N48005, N48006, N48007, N48008, N48009, N48010, N48011, N48012, N48013, N48014, N48015, N48016, N48017, N48018, N48019, N48020, N48021, N48022, N48023, N48024, N48025, N48026, N48027, N48029, N48030, N48031, N48032, N48033, N48034, N48035, N48036, N48037, N48038, N48040, N48041, N48042, N48043, N48044, N48045, N48046, N48047, N48049, N48050, N48051, N48052, N48053, N48054, N48055, N48056, N48058, N48059, N48061, N48062, N48063, N48064, N48065, N48066, N48067, N48068, N48069, N48070, N48071, N48072, N48073, N48074, N48075, N48076, N48077, N48078, N48079, N48080, N48081, N48082, N48083, N48084, N48085, N48087, N48088, N48089, N48090, N48091, N48092, N48093, N48094, N48095, N48096, N48097, N48098, N48099, N48100, N48102, N48103, N48104, N48105, N48106, N48107, N48108, N48109, N48110, N48111, N48113, N48115, N48116, N48117, N48118, N48119, N48120, N48121, N48122, N48123, N48124, N48125, N48126, N48127, N48129, N48130, N48131, N48132, N48133, N48135, N48137, N48138, N48139, N48140, N48141, N48142, N48143, N48145, N48147, N48148, N48149, N48150, N48152, N48153, N48154, N48155, N48156, N48157, N48158, N48159, N48160, N48161, N48162, N48164, N48165, N48167, N48168, N48169, N48170, N48171, N48172, N48173, N48174, N48175, N48176, N48177, N48178, N48179, N48180, N48181, N48182, N48183, N48184, N48185, N48187, N48188, N48189, N48190, N48191, N48192, N48193, N48194, N48195, N48196, N48197, N48198, N48199, N48200, N48201, N48202, N48203, N48204, N48205, N48206, N48207, N48208, N48210, N48211, N48212, N48213, N48214, N48216, N48217, N48219, N48220, N48221, N48222, N48223, N48224, N48225, N48226, N48227, N48228, N48229, N48230, N48231, N48233, N48234, N48235, N48236, N48237, N48238, N48240, N48241, N48242, N48243, N48244, N48245, N48246, N48248, N48249, N48250, N48251, N48252, N48253, N48254, N48255, N48256, N48257, N48258, N48259, N48260, N48262, N48263, N48264, N48265, N48267, N48268, N48269, N48270, N48271, N48272, N48273, N48274, N48275, N48277, N48278, N48279, N48280, N48281, N48282, N48283, N48284, N48286, N48287, N48288, N48289, N48290, N48291, N48292, N48293, N48294, N48295, N48296, N48297, N48298, N48299, N48300, N48302, N48303, N48306, N48307, N48308, N48309, N48311, N48312, N48313, N48314, N48315, N48316, N48317, N48318, N48319, N48320, N48321, N48323, N48325, N48326, N48327, N48328, N48329, N48331, N48332, N48333, N48334, N48335, N48336, N48337, N48338, N48339, N48340, N48341, N48342, N48343, N48344, N48345, N48346, N48347, N48349, N48350, N48351, N48352, N48353, N48354, N48356, N48357, N48358, N48359, N48360, N48362, N48363, N48364, N48365, N48366, N48367, N48368, N48369, N48370, N48371, N48372, N48374, N48375, N48377, N48379, N48380, N48382, N48383, N48384, N48385, N48386, N48387, N48388, N48389, N48390, N48391, N48392, N48393, N48394, N48395, N48396, N48397, N48398, N48399, N48400, N48401, N48404, N48405, N48406, N48407, N48408, N48409, N48410, N48411, N48412, N48413, N48414, N48415, N48416, N48417, N48418, N48419, N48420, N48421, N48422, N48423, N48424, N48425, N48426, N48427, N48428, N48429, N48430, N48431, N48432, N48433, N48435, N48436, N48437, N48438, N48439, N48440, N48441, N48442, N48443, N48444, N48445, N48446, N48447, N48448, N48449, N48450, N48451, N48452, N48454, N48455, N48456, N48457, N48459, N48461, N48462, N48463, N48464, N48465, N48466, N48468, N48469, N48470, N48471, N48472, N48473, N48474, N48475, N48476, N48477, N48478, N48479, N48480, N48481, N48482, N48483, N48484, N48485, N48486, N48488, N48489, N48490, N48491, N48492, N48493, N48494, N48495, N48496, N48497, N48498, N48499, N48500, N48501, N48502, N48503, N48504, N48505, N48506, N48507, N48508, N48511, N48512, N48513, N48515, N48516, N48517, N48518, N48519, N48521, N48523, N48524, N48525, N48526, N48527, N48528, N48529, N48530, N48531, N48532, N48533, N48534, N48535, N48536, N48537, N48538, N48539, N48540, N48541, N48542, N48543, N48545, N48546, N48547, N48549, N48550, N48551, N48552, N48553, N48555, N48557, N48558, N48559, N48560, N48561, N48562, N48563, N48564, N48565, N48566, N48567, N48568, N48569, N48570, N48571, N48572, N48573, N48574, N48575, N48576, N48578, N48579, N48581, N48582, N48583, N48584, N48585, N48586, N48587, N48588, N48589, N48590, N48591, N48592, N48593, N48594, N48595, N48596, N48597, N48598, N48600, N48601, N48602, N48603, N48604, N48605, N48606, N48607, N48609, N48610, N48611, N48612, N48613, N48614, N48615, N48616, N48617, N48618, N48619, N48620, N48621, N48622, N48623, N48624, N48625, N48626, N48627, N48628, N48629, N48630, N48631, N48632, N48633, N48634, N48635, N48636, N48637, N48638, N48639, N48641, N48642, N48643, N48644, N48645, N48646, N48647, N48649, N48650, N48651, N48652, N48653, N48654, N48655, N48656, N48657, N48658, N48659, N48660, N48661, N48662, N48663, N48664, N48665, N48666, N48667, N48668, N48669, N48670, N48671, N48672, N48673, N48674, N48675, N48676, N48677, N48679, N48680, N48681, N48682, N48683, N48684, N48685, N48686, N48687, N48688, N48689, N48690, N48691, N48692, N48693, N48694, N48695, N48696, N48697, N48698, N48699, N48700, N48701, N48702, N48704, N48705, N48706, N48707, N48708, N48709, N48710, N48711, N48712, N48713, N48714, N48715, N48716, N48718, N48720, N48721, N48722, N48723, N48724, N48725, N48726, N48727, N48728, N48729, N48730, N48731, N48732, N48734, N48735, N48736, N48737, N48738, N48739, N48740, N48741, N48742, N48744, N48745, N48746, N48747, N48748, N48749, N48750, N48751, N48752, N48753, N48754, N48755, N48756, N48757, N48758, N48759, N48760, N48762, N48763, N48764, N48765, N48766, N48767, N48768, N48769, N48770, N48771, N48772, N48773, N48774, N48775, N48776, N48777, N48778, N48779, N48780, N48781, N48782, N48783, N48784, N48785, N48786, N48787, N48788, N48789, N48790, N48791, N48792, N48793, N48794, N48795, N48796, N48797, N48798, N48799, N48800, N48801, N48802, N48803, N48804, N48805, N48806, N48807, N48808, N48809, N48810, N48811, N48812, N48813, N48814, N48815, N48817, N48818, N48819, N48820, N48821, N48822, N48823, N48824, N48825, N48826, N48828, N48829, N48830, N48832, N48833, N48835, N48836, N48837, N48838, N48839, N48840, N48841, N48842, N48843, N48844, N48845, N48846, N48847, N48848, N48849, N48850, N48851, N48852, N48853, N48854, N48855, N48856, N48857, N48858, N48859, N48860, N48861, N48862, N48863, N48864, N48865, N48866, N48867, N48868, N48869, N48870, N48871, N48872, N48873, N48874, N48875, N48876, N48877, N48878, N48879, N48880, N48881, N48882, N48883, N48884, N48885, N48886, N48887, N48888, N48889, N48890, N48892, N48894, N48895, N48897, N48898, N48899, N48900, N48901, N48902, N48903, N48904, N48905, N48906, N48907, N48909, N48910, N48911, N48912, N48913, N48914, N48915, N48916, N48917, N48918, N48919, N48920, N48921, N48922, N48923, N48924, N48925, N48926, N48927, N48928, N48929, N48930, N48932, N48933, N48934, N48935, N48936, N48937, N48938, N48939, N48940, N48941, N48943, N48944, N48945, N48946, N48947, N48948, N48949, N48950, N48951, N48952, N48954, N48955, N48956, N48957, N48958, N48959, N48960, N48961, N48962, N48963, N48964, N48965, N48966, N48967, N48969, N48971, N48972, N48973, N48974, N48975, N48977, N48978, N48979, N48980, N48981, N48982, N48983, N48984, N48985, N48986, N48988, N48989, N48990, N48991, N48992, N48994, N48995, N48996, N48997, N48998, N48999, N49000, N49001, N49002, N49003, N49004, N49005, N49006, N49007, N49008, N49009, N49011, N49012, N49013, N49014, N49015, N49016, N49017, N49018, N49019, N49020, N49021, N49022, N49023, N49024, N49025, N49026, N49028, N49030, N49033, N49034, N49035, N49036, N49037, N49038, N49039, N49040, N49041, N49042, N49043, N49044, N49045, N49046, N49048, N49049, N49050, N49051, N49052, N49053, N49054, N49055, N49056, N49057, N49058, N49059, N49060, N49061, N49062, N49063, N49064, N49065, N49066, N49068, N49069, N49070, N49071, N49072, N49073, N49074, N49075, N49076, N49077, N49078, N49079, N49080, N49081, N49082, N49083, N49084, N49085, N49086, N49087, N49088, N49090, N49091, N49092, N49093, N49094, N49095, N49097, N49098, N49099, N49100, N49101, N49102, N49103, N49104, N49105, N49107, N49108, N49109, N49110, N49111, N49112, N49113, N49114, N49115, N49118, N49119, N49120, N49121, N49123, N49124, N49125, N49126, N49127, N49128, N49130, N49131, N49132, N49133, N49135, N49136, N49137, N49138, N49139, N49140, N49141, N49142, N49143, N49144, N49145, N49146, N49147, N49148, N49149, N49150, N49151, N49153, N49154, N49155, N49156, N49157, N49158, N49159, N49160, N49161, N49162, N49163, N49164, N49165, N49166, N49167, N49168, N49169, N49170, N49171, N49172, N49173, N49174, N49175, N49176, N49177, N49178, N49180, N49181, N49182, N49183, N49185, N49186, N49187, N49188, N49189, N49190, N49191, N49192, N49193, N49195, N49196, N49197, N49198, N49199, N49200, N49201, N49202, N49204, N49205, N49206, N49207, N49208, N49209, N49210, N49211, N49212, N49213, N49214, N49215, N49216, N49217, N49218, N49220, N49222, N49223, N49224, N49225, N49226, N49227, N49228, N49229, N49230, N49231, N49232, N49233, N49234, N49235, N49236, N49237, N49239, N49240, N49241, N49242, N49243, N49244, N49245, N49246, N49247, N49248, N49249, N49250, N49251, N49252, N49253, N49254, N49255, N49256, N49257, N49258, N49259, N49260, N49261, N49262, N49263, N49265, N49266, N49267, N49268, N49269, N49270, N49271, N49272, N49274, N49275, N49276, N49277, N49279, N49280, N49281, N49282, N49284, N49285, N49286, N49287, N49288, N49289, N49290, N49291, N49292, N49293, N49294, N49295, N49296, N49297, N49298, N49300, N49301, N49302, N49303, N49304, N49305, N49306, N49308, N49309, N49310, N49311, N49312, N49313, N49314, N49315, N49317, N49318, N49319, N49320, N49321, N49322, N49323, N49324, N49325, N49326, N49327, N49328, N49330, N49331, N49333, N49334, N49335, N49336, N49338, N49339, N49340, N49341, N49342, N49343, N49344, N49345, N49346, N49347, N49348, N49349, N49350, N49351, N49352, N49353, N49354, N49355, N49356, N49357, N49358, N49359, N49360, N49363, N49364, N49366, N49367, N49368, N49369, N49370, N49371, N49372, N49373, N49374, N49375, N49377, N49378, N49380, N49381, N49382, N49383, N49384, N49385, N49386, N49387, N49388, N49389, N49390, N49391, N49392, N49393, N49394, N49395, N49396, N49397, N49398, N49399, N49400, N49401, N49402, N49403, N49404, N49405, N49406, N49407, N49408, N49409, N49410, N49411, N49412, N49413, N49414, N49415, N49416, N49417, N49418, N49419, N49420, N49422, N49423, N49424, N49425, N49426, N49428, N49429, N49430, N49431, N49432, N49433, N49434, N49435, N49436, N49437, N49438, N49439, N49441, N49442, N49443, N49444, N49445, N49446, N49447, N49448, N49449, N49450, N49451, N49452, N49453, N49454, N49456, N49457, N49459, N49460, N49461, N49462, N49463, N49464, N49465, N49467, N49468, N49469, N49470, N49471, N49473, N49474, N49475, N49476, N49477, N49478, N49479, N49480, N49481, N49483, N49484, N49485, N49486, N49487, N49488, N49489, N49490, N49491, N49492, N49493, N49494, N49495, N49496, N49497, N49498, N49499, N49500, N49501, N49502, N49503, N49504, N49506, N49507, N49508, N49509, N49510, N49511, N49512, N49513, N49514, N49515, N49516, N49517, N49518, N49519, N49520, N49521, N49522, N49523, N49524, N49525, N49526, N49527, N49528, N49529, N49530, N49531, N49532, N49533, N49534, N49535, N49536, N49537, N49538, N49539, N49540, N49541, N49542, N49543, N49544, N49545, N49546, N49547, N49548, N49549, N49550, N49551, N49552, N49555, N49556, N49557, N49558, N49559, N49560, N49562, N49563, N49564, N49565, N49566, N49567, N49568, N49569, N49570, N49571, N49572, N49573, N49574, N49575, N49576, N49577, N49578, N49579, N49580, N49581, N49582, N49583, N49584, N49585, N49586, N49587, N49589, N49590, N49591, N49592, N49593, N49594, N49595, N49596, N49597, N49598, N49599, N49600, N49601, N49602, N49603, N49604, N49605, N49606, N49607, N49608, N49609, N49610, N49611, N49612, N49613, N49614, N49616, N49617, N49618, N49619, N49620, N49622, N49624, N49625, N49626, N49628, N49629, N49630, N49631, N49632, N49633, N49634, N49635, N49636, N49637, N49638, N49639, N49640, N49641, N49643, N49644, N49645, N49646, N49647, N49648, N49649, N49650, N49651, N49652, N49653, N49655, N49656, N49657, N49658, N49660, N49661, N49662, N49663, N49664, N49665, N49666, N49667, N49668, N49669, N49670, N49672, N49673, N49674, N49675, N49676, N49677, N49678, N49679, N49680, N49681, N49682, N49683, N49684, N49685, N49687, N49688, N49689, N49690, N49691, N49692, N49693, N49694, N49695, N49696, N49697, N49698, N49699, N49700, N49701, N49702, N49703, N49705, N49706, N49707, N49708, N49709, N49710, N49711, N49712, N49713, N49714, N49715, N49716, N49717, N49718, N49719, N49720, N49721, N49722, N49723, N49724, N49725, N49726, N49727, N49728, N49729, N49730, N49731, N49732, N49733, N49734, N49735, N49736, N49737, N49739, N49740, N49741, N49742, N49743, N49744, N49745, N49746, N49747, N49748, N49749, N49750, N49751, N49752, N49753, N49754, N49755, N49756, N49757, N49758, N49759, N49760, N49761, N49763, N49765, N49767, N49768, N49769, N49770, N49771, N49772, N49773, N49774, N49776, N49777, N49778, N49779, N49780, N49781, N49782, N49783, N49784, N49785, N49787, N49788, N49789, N49790, N49791, N49792, N49794, N49795, N49796, N49797, N49798, N49799, N49800, N49801, N49802, N49803, N49804, N49805, N49806, N49807, N49808, N49809, N49810, N49811, N49812, N49813, N49814, N49815, N49816, N49817, N49818, N49819, N49820, N49821, N49822, N49823, N49824, N49825, N49826, N49827, N49828, N49829, N49830, N49831, N49832, N49835, N49836, N49837, N49838, N49839, N49840, N49841, N49842, N49843, N49844, N49845, N49846, N49847, N49848, N49849, N49850, N49851, N49852, N49853, N49854, N49855, N49856, N49857, N49858, N49860, N49861, N49862, N49863, N49864, N49865, N49866, N49867, N49868, N49869, N49870, N49871, N49872, N49873, N49874, N49875, N49876, N49877, N49878, N49879, N49880, N49881, N49882, N49883, N49884, N49885, N49886, N49887, N49888, N49889, N49890, N49891, N49892, N49894, N49895, N49896, N49898, N49899, N49901, N49903, N49904, N49905, N49906, N49907, N49908, N49909, N49910, N49911, N49912, N49913, N49914, N49915, N49917, N49918, N49919, N49920, N49921, N49923, N49924, N49925, N49926, N49927, N49928, N49929, N49930, N49931, N49932, N49933, N49934, N49935, N49936, N49937, N49938, N49939, N49940, N49941, N49942, N49943, N49944, N49945, N49946, N49947, N49948, N49949, N49950, N49951, N49952, N49953, N49954, N49955, N49956, N49957, N49958, N49959, N49960, N49961, N49962, N49963, N49964, N49965, N49966, N49967, N49969, N49970, N49972, N49973, N49974, N49975, N49976, N49977, N49979, N49980, N49981, N49982, N49983, N49985, N49986, N49987, N49988, N49989, N49991, N49992, N49993, N49994, N49995, N49996, N49997, N49998, N49999, N50000, N50001, N50003, N50004, N50005, N50006, N50007, N50008, N50009, N50010, N50011, N50012, N50013, N50014, N50015, N50016, N50017, N50018, N50019, N50020, N50021, N50022, N50023, N50024, N50025, N50026, N50027, N50028, N50030, N50031, N50032, N50033, N50034, N50035, N50036, N50037, N50038, N50039, N50040, N50041, N50042, N50043, N50044, N50045, N50046, N50047, N50048, N50049, N50050, N50051, N50053, N50054, N50055, N50056, N50057, N50058, N50059, N50060, N50061, N50062, N50063, N50064, N50065, N50066, N50067, N50068, N50069, N50070, N50071, N50072, N50073, N50074, N50075, N50076, N50077, N50078, N50079, N50080, N50081, N50082, N50084, N50085, N50086, N50087, N50089, N50090, N50091, N50092, N50093, N50094, N50095, N50096, N50098, N50099, N50100, N50101, N50102, N50103, N50104, N50105, N50106, N50108, N50109, N50110, N50111, N50113, N50115, N50116, N50117, N50119, N50120, N50121, N50122, N50123, N50124, N50125, N50126, N50129, N50130, N50131, N50132, N50133, N50134, N50135, N50136, N50137, N50138, N50139, N50140, N50142, N50143, N50144, N50145, N50146, N50147, N50148, N50149, N50150, N50151, N50152, N50153, N50154, N50157, N50158, N50159, N50160, N50161, N50162, N50163, N50164, N50165, N50166, N50167, N50168, N50169, N50170, N50171, N50172, N50173, N50174, N50175, N50177, N50179, N50180, N50181, N50182, N50183, N50185, N50186, N50187, N50188, N50189, N50190, N50191, N50192, N50193, N50194, N50195, N50196, N50197, N50200, N50201, N50203, N50204, N50205, N50206, N50208, N50209, N50210, N50211, N50212, N50213, N50214, N50215, N50216, N50217, N50218, N50220, N50221, N50222, N50223, N50224, N50225, N50226, N50227, N50229, N50230, N50231, N50232, N50234, N50235, N50236, N50237, N50238, N50239, N50240, N50241, N50242, N50243, N50244, N50246, N50247, N50248, N50249, N50250, N50251, N50252, N50253, N50254, N50255, N50256, N50258, N50259, N50260, N50262, N50263, N50264, N50265, N50266, N50267, N50268, N50270, N50272, N50273, N50274, N50276, N50277, N50278, N50279, N50280, N50281, N50282, N50283, N50284, N50285, N50286, N50287, N50288, N50289, N50290, N50291, N50292, N50293, N50294, N50295, N50296, N50297, N50298, N50299, N50300, N50301, N50302, N50303, N50304, N50305, N50306, N50307, N50308, N50309, N50310, N50312, N50313, N50315, N50316, N50317, N50318, N50319, N50320, N50321, N50323, N50324, N50325, N50326, N50327, N50328, N50329, N50330, N50331, N50332, N50333, N50334, N50335, N50336, N50337, N50338, N50339, N50340, N50341, N50342, N50343, N50344, N50345, N50346, N50347, N50349, N50350, N50351, N50352, N50353, N50354, N50355, N50356, N50357, N50358, N50359, N50360, N50361, N50362, N50363, N50364, N50366, N50367, N50368, N50369, N50370, N50371, N50372, N50373, N50374, N50375, N50376, N50377, N50378, N50379, N50380, N50381, N50382, N50383, N50384, N50385, N50386, N50387, N50388, N50389, N50390, N50391, N50392, N50393, N50396, N50397, N50398, N50399, N50400, N50401, N50402, N50403, N50404, N50405, N50406, N50407, N50408, N50409, N50410, N50411, N50412, N50413, N50414, N50415, N50416, N50417, N50418, N50419, N50420, N50421, N50422, N50424, N50425, N50426, N50427, N50428, N50429, N50430, N50432, N50433, N50434, N50435, N50436, N50437, N50438, N50439, N50440, N50441, N50442, N50443, N50444, N50445, N50446, N50447, N50448, N50449, N50450, N50451, N50452, N50453, N50454, N50456, N50457, N50458, N50459, N50461, N50462, N50463, N50464, N50465, N50466, N50467, N50468, N50469, N50470, N50471, N50472, N50473, N50474, N50475, N50476, N50477, N50478, N50479, N50480, N50481, N50482, N50483, N50484, N50485, N50486, N50487, N50488, N50489, N50490, N50491, N50492, N50493, N50494, N50495, N50496, N50497, N50498, N50499, N50500, N50501, N50502, N50503, N50504, N50506, N50507, N50508, N50509, N50510, N50512, N50513, N50514, N50515, N50516, N50517, N50518, N50519, N50520, N50521, N50522, N50523, N50524, N50525, N50526, N50527, N50528, N50529, N50530, N50531, N50532, N50533, N50535, N50536, N50537, N50538, N50539, N50540, N50541, N50542, N50543, N50544, N50545, N50546, N50547, N50548, N50549, N50550, N50551, N50552, N50553, N50554, N50555, N50556, N50557, N50558, N50559, N50560, N50561, N50562, N50563, N50564, N50565, N50566, N50567, N50569, N50570, N50571, N50572, N50573, N50574, N50575, N50576, N50577, N50578, N50579, N50580, N50581, N50582, N50583, N50584, N50585, N50586, N50588, N50589, N50590, N50592, N50593, N50596, N50598, N50599, N50600, N50601, N50603, N50604, N50605, N50606, N50607, N50608, N50609, N50610, N50611, N50612, N50613, N50614, N50615, N50616, N50617, N50618, N50619, N50620, N50621, N50622, N50623, N50624, N50625, N50627, N50628, N50629, N50630, N50631, N50632, N50633, N50635, N50636, N50637, N50638, N50639, N50640, N50641, N50642, N50643, N50644, N50645, N50646, N50648, N50649, N50650, N50651, N50652, N50653, N50654, N50655, N50656, N50657, N50658, N50659, N50660, N50661, N50662, N50663, N50664, N50665, N50667, N50668, N50669, N50670, N50671, N50672, N50673, N50674, N50675, N50676, N50677, N50678, N50679, N50680, N50681, N50682, N50683, N50684, N50685, N50687, N50688, N50689, N50690, N50691, N50693, N50694, N50695, N50696, N50697, N50698, N50699, N50700, N50701, N50702, N50703, N50705, N50706, N50707, N50708, N50709, N50710, N50711, N50712, N50713, N50714, N50715, N50716, N50717, N50718, N50719, N50720, N50721, N50722, N50723, N50724, N50725, N50726, N50728, N50729, N50730, N50731, N50732, N50733, N50734, N50735, N50736, N50737, N50738, N50739, N50741, N50742, N50743, N50744, N50745, N50746, N50747, N50748, N50749, N50750, N50751, N50752, N50753, N50754, N50755, N50756, N50757, N50758, N50759, N50760, N50761, N50762, N50763, N50764, N50765, N50766, N50767, N50768, N50769, N50770, N50771, N50772, N50773, N50774, N50775, N50776, N50777, N50778, N50779, N50780, N50781, N50782, N50783, N50784, N50785, N50786, N50787, N50788, N50789, N50790, N50791, N50792, N50793, N50794, N50795, N50796, N50797, N50798, N50799, N50800, N50801, N50802, N50803, N50804, N50805, N50806, N50807, N50808, N50809, N50810, N50811, N50812, N50813, N50814, N50815, N50816, N50817, N50818, N50819, N50820, N50821, N50822, N50824, N50825, N50826, N50827, N50828, N50829, N50830, N50831, N50832, N50833, N50834, N50835, N50836, N50837, N50838, N50839, N50840, N50841, N50842, N50843, N50844, N50845, N50846, N50847, N50848, N50849, N50850, N50851, N50852, N50853, N50855, N50856, N50857, N50858, N50859, N50860, N50862, N50864, N50865, N50866, N50867, N50868, N50869, N50870, N50871, N50872, N50873, N50874, N50875, N50876, N50878, N50879, N50880, N50881, N50882, N50883, N50884, N50885, N50886, N50887, N50888, N50891, N50892, N50893, N50894, N50895, N50896, N50898, N50899, N50900, N50901, N50902, N50903, N50904, N50905, N50906, N50908, N50910, N50911, N50912, N50913, N50914, N50915, N50916, N50918, N50919, N50920, N50921, N50922, N50923, N50924, N50925, N50926, N50927, N50928, N50929, N50930, N50932, N50933, N50934, N50936, N50937, N50939, N50941, N50942, N50944, N50945, N50946, N50949, N50950, N50952, N50953, N50954, N50955, N50956, N50957, N50958, N50959, N50960, N50961, N50962, N50963, N50964, N50965, N50966, N50968, N50969, N50970, N50971, N50972, N50973, N50975, N50976, N50978, N50979, N50980, N50981, N50982, N50983, N50984, N50985, N50986, N50988, N50989, N50990, N50991, N50992, N50993, N50994, N50995, N50996, N50997, N50998, N50999, N51000, N51001, N51002, N51003, N51004, N51005, N51006, N51007, N51008, N51009, N51010, N51011, N51012, N51013, N51014, N51015, N51016, N51017, N51018, N51019, N51020, N51021, N51022, N51023, N51026, N51027, N51028, N51029, N51030, N51031, N51032, N51033, N51034, N51036, N51037, N51039, N51040, N51041, N51043, N51044, N51045, N51047, N51048, N51049, N51050, N51052, N51053, N51054, N51055, N51056, N51057, N51058, N51059, N51060, N51061, N51062, N51064, N51065, N51066, N51067, N51068, N51069, N51070, N51071, N51072, N51073, N51074, N51075, N51076, N51077, N51078, N51079, N51080, N51081, N51082, N51083, N51084, N51085, N51086, N51087, N51089, N51090, N51091, N51093, N51094, N51095, N51096, N51097, N51098, N51101, N51102, N51103, N51105, N51106, N51107, N51108, N51110, N51111, N51112, N51113, N51114, N51115, N51116, N51117, N51118, N51119, N51120, N51121, N51122, N51123, N51124, N51125, N51126, N51127, N51128, N51129, N51130, N51131, N51132, N51133, N51134, N51135, N51136, N51137, N51139, N51140, N51141, N51142, N51143, N51144, N51145, N51146, N51147, N51148, N51150, N51151, N51152, N51153, N51154, N51155, N51156, N51157, N51159, N51160, N51161, N51162, N51163, N51164, N51165, N51166, N51167, N51168, N51169, N51170, N51171, N51172, N51173, N51174, N51175, N51176, N51177, N51178, N51179, N51180, N51181, N51182, N51183, N51184, N51185, N51186, N51187, N51188, N51189, N51190, N51191, N51193, N51194, N51195, N51197, N51198, N51200, N51201, N51202, N51203, N51204, N51205, N51206, N51207, N51208, N51209, N51210, N51211, N51212, N51213, N51214, N51215, N51216, N51217, N51219, N51220, N51221, N51222, N51223, N51224, N51225, N51226, N51228, N51229, N51230, N51231, N51232, N51233, N51234, N51235, N51236, N51237, N51238, N51239, N51240, N51242, N51244, N51245, N51246, N51248, N51249, N51250, N51251, N51252, N51253, N51254, N51255, N51256, N51257, N51258, N51259, N51260, N51261, N51262, N51263, N51265, N51266, N51267, N51268, N51269, N51270, N51271, N51272, N51273, N51274, N51276, N51277, N51278, N51279, N51280, N51281, N51282, N51283, N51284, N51285, N51286, N51287, N51288, N51289, N51290, N51291, N51292, N51294, N51295, N51296, N51297, N51298, N51299, N51300, N51301, N51302, N51303, N51304, N51305, N51306, N51308, N51309, N51310, N51311, N51312, N51313, N51314, N51315, N51316, N51317, N51318, N51319, N51320, N51321, N51322, N51324, N51325, N51326, N51327, N51328, N51329, N51331, N51332, N51333, N51334, N51335, N51336, N51338, N51340, N51341, N51342, N51343, N51344, N51345, N51346, N51347, N51348, N51349, N51350, N51351, N51352, N51353, N51355, N51357, N51358, N51359, N51360, N51361, N51362, N51363, N51364, N51365, N51366, N51367, N51368, N51369, N51371, N51372, N51374, N51375, N51376, N51377, N51378, N51379, N51381, N51382, N51383, N51384, N51385, N51386, N51387, N51388, N51389, N51390, N51392, N51394, N51395, N51396, N51397, N51398, N51399, N51400, N51401, N51402, N51403, N51405, N51406, N51407, N51408, N51409, N51410, N51411, N51412, N51413, N51414, N51415, N51416, N51417, N51418, N51419, N51420, N51421, N51422, N51423, N51424, N51425, N51426, N51427, N51428, N51430, N51431, N51432, N51433, N51434, N51435, N51436, N51437, N51438, N51439, N51440, N51441, N51442, N51443, N51444, N51445, N51446, N51447, N51448, N51449, N51450, N51452, N51453, N51454, N51455, N51456, N51457, N51458, N51459, N51460, N51461, N51463, N51464, N51465, N51466, N51467, N51468, N51469, N51470, N51471, N51473, N51474, N51475, N51476, N51477, N51478, N51479, N51480, N51481, N51482, N51483, N51484, N51485, N51486, N51487, N51488, N51489, N51490, N51491, N51492, N51493, N51494, N51495, N51496, N51497, N51499, N51500, N51502, N51504, N51505, N51506, N51507, N51508, N51509, N51510, N51511, N51512, N51513, N51514, N51515, N51517, N51518, N51519, N51520, N51522, N51523, N51524, N51525, N51526, N51527, N51528, N51529, N51530, N51531, N51533, N51534, N51537, N51538, N51539, N51541, N51542, N51543, N51544, N51545, N51546, N51547, N51548, N51550, N51551, N51552, N51553, N51554, N51555, N51556, N51557, N51558, N51559, N51560, N51561, N51562, N51563, N51564, N51565, N51566, N51567, N51568, N51569, N51570, N51572, N51573, N51574, N51575, N51576, N51577, N51578, N51579, N51580, N51581, N51582, N51583, N51584, N51586, N51587, N51588, N51589, N51590, N51591, N51592, N51593, N51594, N51595, N51596, N51597, N51598, N51599, N51600, N51601, N51602, N51603, N51604, N51605, N51606, N51607, N51608, N51609, N51610, N51612, N51613, N51614, N51615, N51616, N51617, N51618, N51619, N51620, N51621, N51622, N51623, N51624, N51625, N51626, N51627, N51628, N51629, N51630, N51631, N51632, N51633, N51634, N51635, N51636, N51637, N51638, N51639, N51640, N51641, N51642, N51643, N51644, N51645, N51646, N51647, N51648, N51649, N51650, N51651, N51652, N51653, N51654, N51655, N51656, N51657, N51658, N51659, N51660, N51661, N51662, N51663, N51664, N51665, N51666, N51667, N51668, N51669, N51670, N51671, N51672, N51673, N51674, N51675, N51676, N51677, N51678, N51679, N51680, N51681, N51682, N51683, N51684, N51685, N51686, N51687, N51688, N51689, N51690, N51691, N51692, N51693, N51694, N51695, N51696, N51697, N51698, N51699, N51700, N51701, N51702, N51703, N51704, N51705, N51706, N51707, N51708, N51709, N51710, N51711, N51712, N51713, N51714, N51715, N51716, N51717, N51718, N51719, N51720, N51721, N51722, N51723, N51724, N51725, N51726, N51727, N51728, N51729, N51730, N51731, N51732, N51733, N51735, N51736, N51737, N51738, N51739, N51740, N51741, N51742, N51743, N51745, N51746, N51747, N51748, N51749, N51750, N51751, N51752, N51754, N51755, N51756, N51757, N51758, N51759, N51760, N51761, N51762, N51763, N51764, N51765, N51766, N51767, N51768, N51769, N51770, N51771, N51772, N51773, N51774, N51775, N51776, N51777, N51778, N51779, N51780, N51781, N51782, N51783, N51784, N51785, N51786, N51787, N51788, N51789, N51790, N51791, N51792, N51793, N51794, N51795, N51796, N51797, N51798, N51799, N51800, N51801, N51802, N51803, N51804, N51805, N51806, N51807, N51808, N51809, N51810, N51811, N51812, N51813, N51814, N51815, N51816, N51817, N51818, N51819, N51820, N51821, N51822, N51823, N51824, N51825, N51826, N51827, N51828, N51829, N51830, N51831, N51832, N51833, N51834, N51835, N51836, N51837, N51838, N51839, N51840, N51841, N51842, N51844, N51845, N51846, N51847, N51848, N51849, N51850, N51851, N51852, N51853, N51854, N51855, N51856, N51857, N51858, N51859, N51860, N51861, N51862, N51863, N51864, N51865, N51867, N51868, N51869, N51870, N51871, N51872, N51873, N51874, N51875, N51876, N51877, N51878, N51879, N51880, N51881, N51882, N51883, N51884, N51885, N51886, N51887, N51888, N51889, N51890, N51891, N51892, N51893, N51894, N51896, N51897, N51898, N51899, N51900, N51901, N51902, N51903, N51904, N51905, N51906, N51907, N51908, N51909, N51910, N51911, N51912, N51913, N51914, N51915, N51916, N51917, N51918, N51919, N51920, N51921, N51922, N51923, N51924, N51926, N51927, N51928, N51929, N51930, N51931, N51932, N51933, N51934, N51935, N51937, N51938, N51939, N51940, N51941, N51942, N51943, N51944, N51945, N51946, N51947, N51948, N51949, N51950, N51951, N51952, N51953, N51954, N51955, N51956, N51957, N51958, N51959, N51960, N51961, N51962, N51963, N51964, N51965, N51966, N51967, N51968, N51969, N51970, N51971, N51973, N51974, N51975, N51976, N51977, N51978, N51979, N51980, N51981, N51982, N51983, N51984, N51985, N51986, N51987, N51988, N51989, N51990, N51991, N51992, N51993, N51994, N51995, N51996, N51997, N51998, N51999, N52000, N52001, N52002, N52003, N52004, N52005, N52006, N52007, N52008, N52009, N52011, N52012, N52013, N52014, N52015, N52016, N52017, N52018, N52019, N52020, N52021, N52022, N52023, N52025, N52026, N52027, N52028, N52029, N52030, N52031, N52032, N52033, N52034, N52035, N52036, N52037, N52038, N52039, N52040, N52041, N52042, N52043, N52044, N52045, N52046, N52047, N52048, N52049, N52050, N52051, N52052, N52053, N52054, N52055, N52056, N52057, N52058, N52059, N52060, N52061, N52062, N52063, N52064, N52065, N52066, N52067, N52069, N52070, N52071, N52072, N52073, N52074, N52075, N52076, N52077, N52078, N52079, N52080, N52081, N52082, N52083, N52085, N52086, N52087, N52089, N52090, N52091, N52092, N52094, N52095, N52096, N52097, N52098, N52099, N52100, N52101, N52102, N52103, N52105, N52106, N52107, N52108, N52109, N52110, N52111, N52112, N52113, N52114, N52115, N52116, N52117, N52118, N52119, N52120, N52121, N52122, N52123, N52124, N52125, N52126, N52127, N52128, N52129, N52130, N52131, N52132, N52133, N52134, N52135, N52136, N52137, N52138, N52139, N52140, N52141, N52142, N52143, N52144, N52145, N52146, N52147, N52148, N52149, N52150, N52151, N52152, N52153, N52154, N52155, N52156, N52157, N52158, N52159, N52160, N52161, N52162, N52163, N52164, N52165, N52166, N52167, N52168, N52169, N52170, N52171, N52172, N52173, N52174, N52175, N52176, N52177, N52178, N52179, N52180, N52182, N52183, N52184, N52185, N52186, N52187, N52188, N52189, N52190, N52191, N52192, N52193, N52194, N52195, N52196, N52197, N52198, N52199, N52200, N52201, N52202, N52203, N52204, N52205, N52207, N52208, N52209, N52210, N52211, N52212, N52213, N52214, N52215, N52216, N52217, N52218, N52219, N52220, N52221, N52222, N52223, N52224, N52225, N52226, N52227, N52228, N52229, N52230, N52231, N52232, N52233, N52234, N52235, N52236, N52237, N52239, N52240, N52241, N52242, N52243, N52244, N52245, N52246, N52247, N52248, N52249, N52250, N52251, N52252, N52253, N52254, N52255, N52256, N52257, N52258, N52259, N52260, N52261, N52262, N52263, N52264, N52265, N52266, N52267, N52268, N52269, N52270, N52271, N52272, N52273, N52274, N52275, N52276, N52277, N52278, N52279, N52280, N52281, N52282, N52283, N52284, N52285, N52286, N52287, N52288, N52289, N52290, N52291, N52292, N52293, N52294, N52295, N52296, N52297, N52298, N52299, N52300, N52301, N52302, N52303, N52304, N52305, N52306, N52307, N52308, N52309, N52310, N52311, N52312, N52313, N52314, N52315, N52316, N52317, N52318, N52319, N52320, N52321, N52322, N52323, N52324, N52325, N52327, N52329, N52330, N52331, N52332, N52333, N52334, N52335, N52336, N52337, N52338, N52339, N52340, N52341, N52342, N52343, N52344, N52345, N52346, N52347, N52348, N52349, N52350, N52351, N52352, N52353, N52354, N52355, N52356, N52357, N52358, N52359, N52360, N52361, N52362, N52363, N52364, N52365, N52366, N52367, N52368, N52369, N52370, N52371, N52372, N52373, N52374, N52375, N52376, N52377, N52378, N52379, N52380, N52381, N52382, N52383, N52384, N52385, N52386, N52387, N52388, N52389, N52390, N52391, N52392, N52393, N52394, N52395, N52396, N52397, N52398, N52399, N52400, N52401, N52402, N52403, N52404, N52405, N52406, N52407, N52408, N52409, N52410, N52411, N52412, N52413, N52414, N52415, N52416, N52417, N52418, N52419, N52420, N52421, N52422, N52423, N52424, N52425, N52426, N52427, N52428, N52429, N52431, N52432, N52433, N52434, N52435, N52436, N52437, N52438, N52439, N52440, N52441, N52442, N52443, N52444, N52445, N52446, N52447, N52448, N52449, N52450, N52451, N52452, N52453, N52455, N52456, N52457, N52458, N52459, N52460, N52461, N52462, N52463, N52464, N52465, N52466, N52467, N52468, N52469, N52470, N52471, N52472, N52473, N52474, N52475, N52476, N52477, N52478, N52479, N52480, N52481, N52482, N52483, N52484, N52485, N52486, N52487, N52488, N52489, N52490, N52491, N52492, N52493, N52494, N52495, N52496, N52497, N52498, N52499, N52500, N52501, N52502, N52503, N52504, N52505, N52506, N52507, N52508, N52509, N52510, N52511, N52512, N52513, N52514, N52515, N52516, N52517, N52519, N52520, N52521, N52522, N52523, N52524, N52525, N52526, N52527, N52528, N52529, N52530, N52531, N52532, N52533, N52534, N52535, N52536, N52537, N52538, N52539, N52540, N52541, N52542, N52543, N52544, N52546, N52547, N52548, N52549, N52550, N52551, N52552, N52553, N52554, N52555, N52556, N52557, N52558, N52559, N52560, N52561, N52562, N52563, N52564, N52565, N52566, N52567, N52568, N52569, N52570, N52571, N52572, N52573, N52574, N52575, N52576, N52578, N52579, N52580, N52581, N52582, N52583, N52584, N52585, N52586, N52587, N52588, N52589, N52590, N52591, N52592, N52593, N52594, N52595, N52596, N52597, N52598, N52599, N52600, N52601, N52602, N52603, N52604, N52606, N52608, N52609, N52610, N52611, N52613, N52614, N52615, N52616, N52617, N52618, N52619, N52620, N52621, N52622, N52623, N52624, N52625, N52626, N52627, N52628, N52629, N52630, N52631, N52632, N52633, N52634, N52636, N52637, N52638, N52639, N52640, N52641, N52642, N52643, N52644, N52645, N52646, N52647, N52648, N52649, N52650, N52651, N52652, N52653, N52654, N52655, N52656, N52657, N52658, N52659, N52661, N52662, N52663, N52664, N52665, N52666, N52667, N52668, N52669, N52670, N52671, N52672, N52673, N52674, N52675, N52676, N52677, N52678, N52679, N52680, N52681, N52682, N52683, N52684, N52685, N52686, N52687, N52688, N52689, N52690, N52691, N52692, N52693, N52694, N52695, N52696, N52697, N52698, N52699, N52700, N52701, N52702, N52703, N52704, N52705, N52706, N52707, N52708, N52709, N52710, N52711, N52712, N52713, N52714, N52715, N52716, N52717, N52718, N52719, N52720, N52721, N52722, N52723, N52724, N52725, N52726, N52727, N52728, N52729, N52730, N52731, N52732, N52733, N52734, N52735, N52736, N52737, N52738, N52739, N52740, N52741, N52742, N52743, N52744, N52745, N52746, N52747, N52748, N52749, N52750, N52751, N52752, N52753, N52754, N52755, N52756, N52757, N52758, N52759, N52760, N52761, N52762, N52763, N52764, N52765, N52766, N52767, N52768, N52769, N52770, N52771, N52772, N52773, N52774, N52775, N52776, N52777, N52778, N52779, N52780, N52781, N52782, N52783, N52784, N52785, N52786, N52787, N52788, N52789, N52790, N52791, N52792, N52793, N52794, N52795, N52796, N52797, N52798, N52800, N52801, N52802, N52803, N52804, N52805, N52806, N52807, N52808, N52809, N52810, N52811, N52812, N52814, N52815, N52816, N52817, N52818, N52819, N52820, N52821, N52822, N52823, N52824, N52825, N52826, N52827, N52828, N52829, N52830, N52831, N52832, N52833, N52834, N52835, N52836, N52838, N52839, N52840, N52841, N52842, N52843, N52844, N52845, N52846, N52847, N52848, N52849, N52850, N52851, N52852, N52853, N52854, N52855, N52856, N52857, N52858, N52859, N52860, N52861, N52862, N52863, N52864, N52865, N52866, N52867, N52868, N52869, N52870, N52871, N52872, N52873, N52874, N52875, N52876, N52877, N52878, N52879, N52880, N52882, N52883, N52884, N52885, N52886, N52887, N52888, N52889, N52890, N52891, N52892, N52893, N52894, N52895, N52896, N52897, N52898, N52899, N52900, N52901, N52902, N52903, N52904, N52905, N52906, N52907, N52908, N52909, N52910, N52911, N52912, N52913, N52914, N52915, N52916, N52917, N52918, N52919, N52920, N52921, N52922, N52923, N52924, N52925, N52926, N52927, N52928, N52929, N52930, N52931, N52932, N52933, N52934, N52935, N52936, N52937, N52938, N52940, N52941, N52942, N52943, N52944, N52945, N52946, N52947, N52948, N52949, N52950, N52951, N52952, N52953, N52954, N52955, N52956, N52957, N52958, N52959, N52960, N52961, N52962, N52963, N52964, N52965, N52967, N52968, N52969, N52970, N52971, N52972, N52973, N52974, N52975, N52976, N52977, N52978, N52979, N52980, N52981, N52982, N52983, N52984, N52985, N52986, N52987, N52988, N52989, N52990, N52991, N52992, N52993, N52994, N52995, N52996, N52997, N52998, N52999, N53000, N53001, N53002, N53003, N53004, N53005, N53006, N53007, N53008, N53009, N53010, N53011, N53012, N53013, N53014, N53015, N53016, N53017, N53018, N53019, N53020, N53021, N53022, N53024, N53025, N53026, N53028, N53029, N53030, N53031, N53032, N53033, N53034, N53035, N53036, N53037, N53038, N53039, N53040, N53041, N53042, N53043, N53044, N53045, N53046, N53047, N53048, N53049, N53050, N53051, N53052, N53053, N53054, N53055, N53056, N53057, N53058, N53059, N53060, N53061, N53062, N53063, N53064, N53066, N53067, N53068, N53069, N53070, N53071, N53072, N53073, N53074, N53075, N53077, N53078, N53079, N53080, N53081, N53082, N53083, N53084, N53085, N53086, N53087, N53088, N53089, N53090, N53091, N53092, N53093, N53094, N53095, N53096, N53097, N53098, N53099, N53100, N53101, N53102, N53103, N53104, N53105, N53106, N53107, N53108, N53109, N53110, N53111, N53112, N53113, N53114, N53115, N53116, N53117, N53118, N53119, N53120, N53121, N53122, N53123, N53124, N53125, N53126, N53127, N53128, N53129, N53130, N53131, N53132, N53133, N53134, N53135, N53136, N53137, N53138, N53139, N53140, N53141, N53142, N53143, N53144, N53145, N53146, N53147, N53148, N53149, N53150, N53151, N53152, N53153, N53154, N53155, N53156, N53157, N53158, N53159, N53160, N53161, N53162, N53163, N53164, N53165, N53166, N53167, N53168, N53169, N53170, N53171, N53172, N53173, N53174, N53175, N53176, N53177, N53178, N53179, N53180, N53181, N53182, N53183, N53184, N53185, N53186, N53187, N53188, N53189, N53190, N53191, N53192, N53193, N53194, N53195, N53196, N53197, N53198, N53199, N53200, N53201, N53202, N53204, N53205, N53206, N53207, N53208, N53209, N53210, N53211, N53212, N53213, N53214, N53215, N53216, N53217, N53218, N53219, N53220, N53221, N53222, N53223, N53224, N53225, N53226, N53227, N53228, N53229, N53230, N53231, N53233, N53234, N53235, N53236, N53237, N53238, N53239, N53240, N53241, N53242, N53243, N53244, N53245, N53246, N53247, N53248, N53249, N53250, N53251, N53252, N53253, N53254, N53255, N53256, N53257, N53258, N53259, N53260, N53261, N53262, N53263, N53264, N53265, N53266, N53267, N53268, N53269, N53270, N53271, N53272, N53273, N53274, N53275, N53276, N53277, N53278, N53279, N53280, N53281, N53282, N53283, N53284, N53285, N53286, N53287, N53288, N53289, N53290, N53291, N53292, N53293, N53294, N53295, N53296, N53297, N53298, N53299, N53300, N53301, N53302, N53303, N53304, N53305, N53306, N53307, N53308, N53309, N53310, N53311, N53312, N53313, N53314, N53315, N53316, N53317, N53318, N53319, N53320, N53321, N53322, N53323, N53325, N53326, N53327, N53328, N53329, N53330, N53331, N53332, N53333, N53334, N53335, N53336, N53337, N53338, N53339, N53340, N53341, N53342, N53343, N53344, N53345, N53346, N53347, N53348, N53349, N53350, N53351, N53353, N53354, N53355, N53356, N53357, N53358, N53359, N53360, N53361, N53363, N53364, N53366, N53367, N53368, N53369, N53370, N53371, N53372, N53373, N53374, N53375, N53376, N53377, N53378, N53379, N53380, N53381, N53382, N53383, N53384, N53385, N53386, N53387, N53388, N53389, N53390, N53391, N53393, N53394, N53395, N53396, N53397, N53398, N53399, N53400, N53401, N53402, N53403, N53404, N53405, N53406, N53407, N53408, N53409, N53410, N53411, N53412, N53413, N53414, N53415, N53416, N53417, N53418, N53419, N53420, N53421, N53422, N53423, N53424, N53425, N53426, N53427, N53428, N53429, N53430, N53431, N53432, N53433, N53434, N53435, N53436, N53437, N53438, N53439, N53440, N53441, N53442, N53443, N53444, N53445, N53446, N53447, N53448, N53449, N53450, N53451, N53452, N53454, N53455, N53456, N53457, N53458, N53459, N53460, N53461, N53462, N53463, N53464, N53465, N53466, N53467, N53468, N53469, N53470, N53471, N53472, N53473, N53474, N53475, N53476, N53477, N53478, N53479, N53480, N53481, N53482, N53483, N53484, N53485, N53486, N53487, N53488, N53489, N53490, N53491, N53492, N53493, N53494, N53495, N53496, N53497, N53498, N53499, N53500, N53501, N53502, N53503, N53504, N53505, N53506, N53507, N53508, N53509, N53510, N53511, N53512, N53513, N53514, N53515, N53516, N53517, N53518, N53519, N53520, N53521, N53522, N53523, N53524, N53525, N53526, N53527, N53528, N53529, N53530, N53531, N53532, N53533, N53534, N53535, N53536, N53537, N53538, N53539, N53540, N53541, N53542, N53543, N53544, N53545, N53546, N53547, N53548, N53549, N53550, N53551, N53552, N53553, N53554, N53555, N53556, N53557, N53558, N53559, N53560, N53561, N53562, N53563, N53564, N53565, N53566, N53567, N53568, N53569, N53570, N53571, N53572, N53573, N53574, N53575, N53576, N53577, N53578, N53579, N53580, N53581, N53582, N53583, N53584, N53585, N53586, N53587, N53588, N53589, N53590, N53591, N53592, N53593, N53594, N53595, N53596, N53597, N53598, N53599, N53601, N53602, N53603, N53604, N53605, N53606, N53607, N53608, N53609, N53610, N53611, N53612, N53613, N53614, N53615, N53616, N53617, N53618, N53619, N53620, N53621, N53622, N53623, N53624, N53625, N53626, N53627, N53628, N53629, N53630, N53632, N53633, N53634, N53635, N53636, N53637, N53638, N53639, N53640, N53641, N53642, N53643, N53644, N53645, N53646, N53647, N53648, N53649, N53650, N53651, N53652, N53653, N53654, N53655, N53656, N53657, N53658, N53659, N53660, N53661, N53662, N53663, N53664, N53665, N53666, N53667, N53668, N53669, N53670, N53671, N53672, N53673, N53674, N53675, N53676, N53677, N53678, N53679, N53680, N53681, N53682, N53683, N53684, N53685, N53686, N53687, N53688, N53689, N53690, N53691, N53692, N53693, N53694, N53695, N53696, N53697, N53698, N53699, N53700, N53701, N53702, N53703, N53704, N53705, N53706, N53707, N53708, N53709, N53710, N53711, N53712, N53713, N53714, N53715, N53716, N53717, N53718, N53719, N53720, N53721, N53722, N53723, N53724, N53725, N53726, N53727, N53728, N53729, N53730, N53731, N53732, N53733, N53734, N53735, N53736, N53737, N53738, N53739, N53740, N53741, N53742, N53743, N53744, N53745, N53746, N53747, N53748, N53749, N53750, N53751, N53752, N53753, N53754, N53755, N53756, N53757, N53758, N53759, N53760, N53761, N53762, N53763, N53764, N53765, N53766, N53767, N53768, N53769, N53770, N53771, N53772, N53773, N53774, N53775, N53776, N53777, N53778, N53779, N53780, N53781, N53782, N53783, N53784, N53785, N53786, N53787, N53788, N53789, N53790, N53791, N53792, N53793, N53794, N53795, N53796, N53797, N53798, N53800, N53801, N53802, N53803, N53804, N53805, N53806, N53807, N53808, N53809, N53810, N53811, N53812, N53813, N53814, N53815, N53816, N53817, N53818, N53819, N53820, N53821, N53822, N53823, N53824, N53825, N53826, N53827, N53828, N53829, N53830, N53831, N53832, N53833, N53834, N53835, N53836, N53837, N53838, N53839, N53840, N53841, N53842, N53843, N53844, N53845, N53846, N53847, N53848, N53849, N53850, N53851, N53852, N53853, N53854, N53855, N53856, N53857, N53858, N53859, N53860, N53861, N53863, N53864, N53865, N53866, N53867, N53868, N53869, N53870, N53871, N53872, N53873, N53874, N53875, N53876, N53877, N53878, N53879, N53880, N53881, N53882, N53883, N53884, N53885, N53886, N53887, N53888, N53889, N53890, N53891, N53892, N53893, N53894, N53895, N53896, N53897, N53898, N53899, N53900, N53901, N53902, N53903, N53904, N53905, N53906, N53907, N53908, N53909, N53910, N53911, N53912, N53913, N53914, N53915, N53916, N53917, N53918, N53919, N53920, N53921, N53922, N53923, N53924, N53925, N53926, N53927, N53928, N53929, N53930, N53931, N53932, N53933, N53934, N53935, N53936, N53937, N53938, N53939, N53940, N53941, N53942, N53943, N53944, N53945, N53946, N53947, N53948, N53949, N53950, N53951, N53952, N53953, N53954, N53955, N53956, N53957, N53958, N53959, N53960, N53961, N53962, N53963, N53964, N53965, N53966, N53967, N53968, N53969, N53970, N53971, N53972, N53973, N53974, N53975, N53976, N53977, N53978, N53979, N53980, N53981, N53982, N53983, N53984, N53985, N53986, N53987, N53988, N53989, N53990, N53991, N53992, N53993, N53994, N53996, N53997, N53998, N53999, N54000, N54001, N54002, N54003, N54004, N54005, N54006, N54007, N54008, N54009, N54010, N54011, N54012, N54013, N54014, N54015, N54016, N54017, N54018, N54019, N54020, N54021, N54022, N54023, N54024, N54025, N54026, N54027, N54028, N54029, N54030, N54031, N54032, N54033, N54034, N54035, N54036, N54037, N54038, N54039, N54040, N54041, N54042, N54043, N54044, N54045, N54046, N54047, N54048, N54049, N54050, N54051, N54052, N54053, N54054, N54055, N54056, N54057, N54058, N54059, N54060, N54061, N54062, N54063, N54064, N54065, N54066, N54067, N54068, N54069, N54071, N54072, N54073, N54074, N54075, N54076, N54077, N54078, N54079, N54080, N54081, N54082, N54083, N54084, N54085, N54086, N54087, N54088, N54089, N54090, N54091, N54092, N54093, N54094, N54095, N54096, N54097, N54098, N54099, N54100, N54101, N54102, N54103, N54104, N54105, N54106, N54107, N54108, N54109, N54110, N54111, N54112, N54113, N54114, N54115, N54116, N54117, N54118, N54119, N54120, N54121, N54122, N54123, N54124, N54125, N54126, N54127, N54128, N54129, N54130, N54131, N54132, N54133, N54134, N54135, N54136, N54137, N54138, N54139, N54140, N54141, N54142, N54143, N54144, N54145, N54146, N54147, N54148, N54149, N54150, N54151, N54152, N54153, N54154, N54155, N54156, N54157, N54158, N54159, N54160, N54161, N54162, N54163, N54164, N54165, N54166, N54167, N54168, N54169, N54170, N54171, N54172, N54173, N54174, N54175, N54176, N54177, N54178, N54179, N54180, N54181, N54182, N54183, N54184, N54185, N54186, N54187, N54188, N54189, N54190, N54191, N54192, N54193, N54194, N54195, N54196, N54197, N54198, N54199, N54200, N54201, N54202, N54203, N54204, N54205, N54206, N54207, N54208, N54209, N54210, N54211, N54212, N54213, N54214, N54215, N54216, N54217, N54218, N54219, N54220, N54221, N54222, N54223, N54224, N54225, N54226, N54227, N54228, N54229, N54230, N54231, N54232, N54233, N54234, N54235, N54236, N54237, N54238, N54239, N54240, N54241, N54242, N54243, N54244, N54245, N54246, N54247, N54248, N54249, N54250, N54251, N54252, N54253, N54254, N54255, N54256, N54257, N54258, N54259, N54260, N54261, N54262, N54263, N54264, N54265, N54266, N54267, N54268, N54269, N54270, N54271, N54272, N54273, N54274, N54275, N54276, N54277, N54278, N54279, N54280, N54281, N54282, N54283, N54284, N54285, N54286, N54287, N54288, N54289, N54290, N54291, N54292, N54293, N54294, N54295, N54296, N54297, N54298, N54299, N54300, N54301, N54302, N54303, N54304, N54305, N54306, N54307, N54308, N54309, N54310, N54311, N54312, N54313, N54314, N54315, N54316, N54317, N54318, N54319, N54320, N54321;
    wire n12873, n12875, n12876, n12878, n12879, n12880, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12893, n12894, n12895, n12896, n12898, n12900, n12901, n12902, n12903, n12904, n12906, n12907, n12909, n12910, n12912, n12913, n12914, n12915, n12917, n12919, n12921, n12922, n12923, n12926, n12927, n12928, n12929, n12930, n12932, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12944, n12945, n12946, n12947, n12948, n12950, n12951, n12953, n12954, n12955, n12956, n12957, n12959, n12960, n12961, n12962, n12963, n12964, n12966, n12967, n12968, n12970, n12971, n12972, n12974, n12975, n12976, n12977, n12978, n12979, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12992, n12993, n12994, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13009, n13010, n13011, n13012, n13013, n13014, n13016, n13017, n13018, n13019, n13020, n13022, n13025, n13026, n13027, n13029, n13030, n13031, n13032, n13034, n13036, n13037, n13038, n13039, n13041, n13042, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13066, n13067, n13068, n13069, n13070, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13119, n13121, n13122, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13155, n13156, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13166, n13167, n13169, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13183, n13184, n13185, n13186, n13187, n13188, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13201, n13202, n13203, n13204, n13205, n13207, n13208, n13209, n13210, n13212, n13213, n13214, n13215, n13216, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13226, n13227, n13229, n13230, n13231, n13232, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13251, n13252, n13253, n13254, n13255, n13256, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13278, n13279, n13280, n13281, n13282, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13308, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13328, n13329, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13340, n13341, n13343, n13344, n13345, n13346, n13347, n13349, n13350, n13351, n13352, n13354, n13355, n13356, n13357, n13358, n13359, n13363, n13364, n13365, n13366, n13367, n13368, n13370, n13371, n13372, n13374, n13375, n13378, n13379, n13380, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13409, n13411, n13412, n13413, n13414, n13416, n13417, n13418, n13419, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13432, n13433, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13445, n13447, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13459, n13460, n13461, n13462, n13463, n13464, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13484, n13485, n13486, n13487, n13488, n13489, n13491, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13506, n13507, n13508, n13509, n13510, n13511, n13513, n13515, n13516, n13518, n13519, n13520, n13521, n13522, n13523, n13525, n13526, n13528, n13529, n13530, n13531, n13532, n13534, n13535, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13549, n13550, n13552, n13553, n13554, n13555, n13557, n13558, n13559, n13560, n13561, n13562, n13564, n13565, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13590, n13591, n13592, n13593, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13609, n13613, n13614, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13629, n13630, n13631, n13632, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13648, n13649, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13664, n13665, n13667, n13668, n13669, n13670, n13671, n13672, n13675, n13676, n13677, n13678, n13680, n13682, n13683, n13685, n13687, n13688, n13689, n13690, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13701, n13702, n13703, n13704, n13705, n13706, n13708, n13709, n13710, n13712, n13713, n13714, n13715, n13716, n13717, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13735, n13736, n13738, n13739, n13740, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13762, n13763, n13764, n13765, n13766, n13768, n13769, n13771, n13772, n13773, n13774, n13777, n13778, n13779, n13780, n13782, n13783, n13784, n13786, n13787, n13788, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13804, n13805, n13807, n13808, n13810, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13839, n13840, n13841, n13843, n13845, n13846, n13848, n13849, n13850, n13851, n13853, n13854, n13855, n13856, n13857, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13868, n13871, n13872, n13874, n13875, n13876, n13877, n13878, n13879, n13881, n13882, n13883, n13884, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13894, n13895, n13897, n13898, n13899, n13900, n13902, n13903, n13904, n13907, n13908, n13909, n13911, n13912, n13913, n13914, n13916, n13917, n13918, n13919, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13930, n13931, n13933, n13935, n13936, n13937, n13938, n13939, n13940, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13957, n13958, n13960, n13961, n13962, n13963, n13964, n13966, n13967, n13968, n13970, n13971, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14001, n14002, n14003, n14004, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14035, n14036, n14038, n14039, n14041, n14042, n14043, n14044, n14046, n14047, n14048, n14049, n14050, n14051, n14053, n14054, n14055, n14057, n14058, n14059, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14080, n14081, n14082, n14083, n14085, n14086, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14102, n14103, n14105, n14106, n14108, n14109, n14110, n14111, n14112, n14114, n14115, n14116, n14117, n14118, n14120, n14121, n14122, n14123, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14148, n14149, n14150, n14152, n14153, n14154, n14155, n14156, n14157, n14160, n14162, n14163, n14164, n14166, n14167, n14168, n14169, n14170, n14172, n14173, n14175, n14176, n14177, n14178, n14179, n14181, n14182, n14183, n14184, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14204, n14206, n14209, n14210, n14211, n14213, n14218, n14220, n14221, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14270, n14271, n14272, n14273, n14276, n14277, n14278, n14279, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14290, n14292, n14293, n14294, n14295, n14297, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14312, n14313, n14314, n14315, n14316, n14317, n14319, n14320, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14348, n14349, n14350, n14351, n14353, n14356, n14357, n14358, n14360, n14362, n14363, n14364, n14365, n14366, n14367, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14383, n14384, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14418, n14419, n14420, n14421, n14422, n14423, n14425, n14426, n14427, n14430, n14431, n14432, n14434, n14435, n14437, n14438, n14439, n14440, n14442, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14454, n14456, n14457, n14458, n14459, n14460, n14461, n14463, n14464, n14465, n14466, n14467, n14468, n14470, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14500, n14501, n14503, n14504, n14505, n14506, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14516, n14517, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14547, n14548, n14549, n14550, n14551, n14552, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14564, n14565, n14566, n14567, n14569, n14571, n14572, n14573, n14574, n14575, n14576, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14595, n14596, n14597, n14598, n14599, n14601, n14602, n14605, n14607, n14609, n14610, n14611, n14612, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14664, n14665, n14667, n14668, n14669, n14670, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14681, n14682, n14683, n14684, n14686, n14687, n14688, n14689, n14690, n14692, n14693, n14695, n14696, n14697, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14710, n14711, n14712, n14713, n14714, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14734, n14735, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14753, n14754, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14784, n14786, n14787, n14788, n14789, n14790, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14825, n14827, n14828, n14829, n14830, n14832, n14833, n14834, n14835, n14836, n14838, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14864, n14865, n14866, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14877, n14878, n14879, n14880, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14921, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14932, n14933, n14934, n14935, n14937, n14938, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14948, n14949, n14950, n14951, n14952, n14954, n14955, n14956, n14957, n14959, n14960, n14962, n14963, n14964, n14965, n14966, n14967, n14970, n14972, n14973, n14974, n14975, n14976, n14977, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15003, n15004, n15007, n15008, n15009, n15010, n15011, n15012, n15014, n15016, n15017, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15033, n15034, n15036, n15037, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15072, n15073, n15074, n15076, n15077, n15079, n15080, n15081, n15082, n15083, n15084, n15086, n15087, n15088, n15089, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15102, n15103, n15106, n15108, n15109, n15112, n15113, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15145, n15146, n15147, n15149, n15150, n15151, n15153, n15154, n15155, n15157, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15172, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15184, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15200, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15210, n15211, n15212, n15213, n15215, n15216, n15218, n15219, n15220, n15221, n15222, n15223, n15225, n15226, n15227, n15229, n15230, n15231, n15232, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15250, n15251, n15252, n15253, n15256, n15258, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15275, n15276, n15277, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15292, n15293, n15295, n15297, n15298, n15299, n15300, n15301, n15302, n15305, n15306, n15309, n15311, n15312, n15314, n15315, n15316, n15318, n15320, n15321, n15322, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15347, n15348, n15349, n15350, n15351, n15352, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15363, n15364, n15365, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15404, n15405, n15406, n15407, n15408, n15409, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15443, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15454, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15470, n15471, n15472, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15486, n15487, n15488, n15490, n15491, n15492, n15493, n15495, n15498, n15499, n15502, n15503, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15514, n15515, n15517, n15518, n15521, n15523, n15524, n15525, n15526, n15527, n15528, n15530, n15531, n15533, n15535, n15536, n15538, n15539, n15542, n15544, n15546, n15547, n15548, n15549, n15551, n15552, n15553, n15554, n15555, n15557, n15558, n15559, n15560, n15562, n15563, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15573, n15574, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15639, n15640, n15641, n15642, n15644, n15645, n15647, n15648, n15649, n15650, n15651, n15652, n15654, n15655, n15656, n15657, n15658, n15659, n15661, n15662, n15663, n15665, n15666, n15667, n15668, n15669, n15671, n15672, n15674, n15675, n15676, n15679, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15692, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15706, n15707, n15710, n15712, n15713, n15714, n15716, n15717, n15718, n15720, n15721, n15723, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15739, n15742, n15743, n15744, n15745, n15746, n15747, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15757, n15758, n15759, n15760, n15762, n15763, n15764, n15765, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15789, n15790, n15791, n15792, n15794, n15796, n15797, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15820, n15821, n15822, n15824, n15825, n15826, n15827, n15829, n15830, n15832, n15833, n15834, n15838, n15839, n15840, n15841, n15842, n15843, n15845, n15846, n15848, n15849, n15850, n15851, n15853, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15891, n15892, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15909, n15911, n15912, n15913, n15914, n15915, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15930, n15931, n15932, n15933, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15949, n15950, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15964, n15965, n15966, n15967, n15968, n15971, n15972, n15973, n15974, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15985, n15986, n15987, n15988, n15989, n15990, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16011, n16013, n16015, n16016, n16017, n16018, n16019, n16021, n16023, n16024, n16025, n16027, n16028, n16030, n16031, n16032, n16033, n16034, n16037, n16038, n16039, n16040, n16041, n16043, n16044, n16045, n16047, n16048, n16049, n16051, n16052, n16053, n16054, n16055, n16056, n16059, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16080, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16114, n16115, n16117, n16119, n16120, n16122, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16134, n16135, n16136, n16137, n16139, n16140, n16141, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16155, n16156, n16157, n16158, n16159, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16171, n16172, n16173, n16174, n16175, n16176, n16178, n16179, n16180, n16181, n16182, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16192, n16194, n16195, n16196, n16199, n16200, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16211, n16212, n16213, n16214, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16232, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16275, n16276, n16277, n16279, n16280, n16281, n16284, n16285, n16286, n16287, n16288, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16302, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16324, n16325, n16327, n16329, n16331, n16333, n16335, n16336, n16337, n16338, n16339, n16340, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16365, n16366, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16380, n16381, n16382, n16383, n16384, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16395, n16396, n16397, n16399, n16401, n16404, n16405, n16406, n16407, n16408, n16410, n16411, n16412, n16413, n16414, n16415, n16418, n16419, n16420, n16422, n16423, n16424, n16425, n16426, n16427, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16451, n16452, n16454, n16455, n16456, n16459, n16460, n16461, n16463, n16464, n16465, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16475, n16476, n16477, n16478, n16479, n16481, n16482, n16483, n16484, n16485, n16486, n16488, n16489, n16490, n16491, n16492, n16493, n16495, n16496, n16497, n16498, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16517, n16518, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16528, n16530, n16531, n16532, n16534, n16535, n16536, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16552, n16553, n16554, n16555, n16557, n16558, n16559, n16561, n16562, n16563, n16564, n16566, n16567, n16568, n16569, n16570, n16572, n16573, n16574, n16575, n16577, n16579, n16580, n16581, n16583, n16584, n16585, n16587, n16588, n16589, n16590, n16593, n16594, n16595, n16596, n16597, n16599, n16600, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16630, n16633, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16643, n16644, n16646, n16647, n16648, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16668, n16669, n16670, n16671, n16672, n16673, n16675, n16676, n16678, n16679, n16680, n16681, n16683, n16685, n16686, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16726, n16727, n16728, n16729, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16739, n16740, n16741, n16743, n16744, n16745, n16746, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16761, n16762, n16763, n16764, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16798, n16799, n16800, n16802, n16804, n16805, n16807, n16808, n16810, n16811, n16812, n16813, n16815, n16816, n16817, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16829, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16840, n16842, n16843, n16844, n16845, n16849, n16850, n16851, n16852, n16853, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16868, n16869, n16870, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16880, n16881, n16882, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16907, n16908, n16909, n16910, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16921, n16922, n16923, n16924, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16941, n16943, n16944, n16945, n16946, n16947, n16948, n16950, n16951, n16952, n16953, n16955, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16982, n16983, n16985, n16986, n16987, n16988, n16989, n16991, n16992, n16993, n16994, n16995, n16997, n16998, n17000, n17001, n17003, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17020, n17021, n17022, n17023, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17042, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17064, n17065, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17077, n17078, n17079, n17080, n17081, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17092, n17093, n17094, n17096, n17097, n17099, n17100, n17101, n17103, n17104, n17105, n17108, n17109, n17111, n17112, n17113, n17114, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17125, n17126, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17142, n17143, n17144, n17145, n17146, n17147, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17184, n17185, n17186, n17187, n17189, n17190, n17192, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17204, n17205, n17206, n17207, n17208, n17211, n17212, n17213, n17215, n17217, n17218, n17220, n17222, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17237, n17238, n17239, n17240, n17241, n17242, n17244, n17245, n17246, n17247, n17248, n17249, n17253, n17254, n17256, n17257, n17258, n17259, n17261, n17262, n17263, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17275, n17276, n17277, n17279, n17280, n17281, n17282, n17283, n17284, n17286, n17287, n17288, n17289, n17290, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17302, n17303, n17305, n17306, n17307, n17308, n17309, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17319, n17320, n17321, n17322, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17336, n17338, n17339, n17340, n17341, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17361, n17363, n17364, n17365, n17366, n17368, n17370, n17371, n17372, n17373, n17374, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17394, n17395, n17396, n17398, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17426, n17427, n17429, n17430, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17447, n17448, n17449, n17450, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17461, n17462, n17463, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17481, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17522, n17524, n17525, n17527, n17528, n17530, n17531, n17532, n17533, n17534, n17535, n17538, n17539, n17540, n17541, n17543, n17545, n17546, n17547, n17549, n17551, n17552, n17553, n17554, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17572, n17573, n17574, n17575, n17576, n17577, n17580, n17581, n17583, n17584, n17585, n17587, n17588, n17589, n17592, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17602, n17603, n17605, n17606, n17607, n17608, n17610, n17611, n17613, n17615, n17616, n17617, n17618, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17643, n17644, n17645, n17646, n17647, n17648, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17663, n17664, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17702, n17703, n17704, n17705, n17706, n17708, n17710, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17720, n17721, n17722, n17724, n17725, n17726, n17729, n17730, n17731, n17732, n17733, n17734, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17746, n17747, n17748, n17750, n17751, n17752, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17767, n17768, n17769, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17795, n17796, n17797, n17798, n17799, n17801, n17802, n17803, n17805, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17833, n17834, n17835, n17836, n17837, n17839, n17840, n17841, n17842, n17844, n17845, n17846, n17848, n17849, n17850, n17851, n17853, n17854, n17855, n17856, n17857, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17886, n17887, n17889, n17890, n17891, n17892, n17893, n17896, n17898, n17899, n17900, n17901, n17902, n17904, n17906, n17907, n17909, n17910, n17913, n17914, n17915, n17916, n17919, n17920, n17921, n17923, n17924, n17926, n17928, n17929, n17930, n17932, n17933, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17946, n17947, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17967, n17968, n17969, n17970, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17994, n17995, n17996, n17998, n18000, n18001, n18002, n18003, n18004, n18006, n18008, n18009, n18011, n18012, n18013, n18014, n18015, n18017, n18018, n18019, n18020, n18021, n18023, n18024, n18025, n18026, n18028, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18055, n18056, n18057, n18059, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18098, n18099, n18100, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18111, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18121, n18122, n18123, n18124, n18125, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18139, n18140, n18141, n18142, n18143, n18145, n18146, n18147, n18148, n18150, n18151, n18152, n18154, n18155, n18156, n18158, n18160, n18161, n18162, n18163, n18164, n18165, n18167, n18168, n18169, n18170, n18171, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18202, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18235, n18236, n18237, n18238, n18239, n18241, n18242, n18243, n18244, n18246, n18247, n18248, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18262, n18263, n18265, n18266, n18268, n18269, n18270, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18280, n18282, n18283, n18284, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18304, n18305, n18306, n18307, n18308, n18309, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18352, n18353, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18363, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18373, n18374, n18376, n18377, n18378, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18417, n18418, n18419, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18431, n18432, n18433, n18434, n18435, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18462, n18463, n18465, n18466, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18485, n18486, n18487, n18489, n18490, n18491, n18492, n18494, n18496, n18497, n18498, n18499, n18500, n18501, n18503, n18504, n18505, n18507, n18508, n18509, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18520, n18521, n18522, n18523, n18525, n18527, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18545, n18546, n18547, n18548, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18562, n18564, n18565, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18577, n18579, n18580, n18581, n18582, n18584, n18585, n18586, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18620, n18621, n18623, n18624, n18625, n18626, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18666, n18667, n18669, n18670, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18686, n18687, n18689, n18690, n18691, n18692, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18725, n18726, n18727, n18728, n18729, n18731, n18732, n18733, n18734, n18735, n18736, n18738, n18740, n18742, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18752, n18753, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18777, n18778, n18779, n18780, n18782, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18800, n18801, n18802, n18803, n18804, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18821, n18823, n18824, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18835, n18836, n18837, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18849, n18851, n18852, n18853, n18854, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18882, n18885, n18886, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18908, n18909, n18910, n18911, n18913, n18914, n18915, n18916, n18917, n18918, n18920, n18922, n18923, n18925, n18926, n18927, n18928, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18938, n18940, n18941, n18942, n18943, n18945, n18946, n18947, n18948, n18950, n18951, n18952, n18953, n18954, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18982, n18985, n18986, n18987, n18989, n18990, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19009, n19010, n19012, n19013, n19014, n19015, n19016, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19034, n19035, n19036, n19037, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19049, n19050, n19052, n19053, n19054, n19055, n19059, n19060, n19061, n19062, n19064, n19065, n19067, n19069, n19071, n19072, n19073, n19074, n19075, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19089, n19090, n19091, n19092, n19093, n19094, n19096, n19098, n19099, n19101, n19102, n19103, n19106, n19107, n19110, n19111, n19114, n19115, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19176, n19177, n19179, n19180, n19181, n19183, n19184, n19185, n19186, n19188, n19189, n19191, n19192, n19193, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19208, n19210, n19211, n19214, n19216, n19217, n19218, n19219, n19221, n19222, n19223, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19243, n19244, n19245, n19249, n19250, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19275, n19276, n19278, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19297, n19298, n19299, n19300, n19301, n19302, n19304, n19305, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19325, n19327, n19328, n19330, n19331, n19332, n19333, n19335, n19336, n19337, n19338, n19339, n19342, n19343, n19344, n19345, n19348, n19349, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19376, n19377, n19378, n19379, n19381, n19382, n19383, n19384, n19385, n19387, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19400, n19401, n19403, n19404, n19405, n19406, n19407, n19408, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19446, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19458, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19475, n19476, n19477, n19478, n19479, n19480, n19483, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19494, n19495, n19496, n19497, n19498, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19525, n19526, n19528, n19529, n19530, n19533, n19535, n19538, n19539, n19540, n19541, n19542, n19544, n19545, n19546, n19547, n19548, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19562, n19563, n19565, n19566, n19569, n19571, n19572, n19573, n19574, n19575, n19576, n19578, n19579, n19580, n19581, n19582, n19584, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19594, n19595, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19618, n19619, n19620, n19621, n19624, n19625, n19626, n19627, n19628, n19629, n19631, n19632, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19669, n19671, n19672, n19674, n19675, n19677, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19687, n19688, n19689, n19690, n19691, n19692, n19694, n19695, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19745, n19749, n19750, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19781, n19782, n19783, n19784, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19817, n19818, n19820, n19821, n19825, n19826, n19827, n19828, n19830, n19831, n19833, n19834, n19835, n19836, n19837, n19838, n19840, n19841, n19842, n19843, n19845, n19846, n19847, n19848, n19849, n19850, n19853, n19854, n19855, n19856, n19857, n19858, n19860, n19861, n19862, n19863, n19865, n19866, n19867, n19868, n19869, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19894, n19895, n19896, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19906, n19907, n19908, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19919, n19922, n19923, n19924, n19925, n19926, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19940, n19941, n19943, n19944, n19945, n19946, n19947, n19949, n19950, n19952, n19954, n19955, n19956, n19957, n19958, n19959, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19987, n19989, n19990, n19991, n19992, n19993, n19994, n19996, n19997, n19999, n20000, n20001, n20004, n20005, n20006, n20008, n20009, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20037, n20038, n20039, n20040, n20041, n20043, n20044, n20045, n20046, n20049, n20050, n20051, n20052, n20053, n20054, n20056, n20058, n20061, n20062, n20063, n20064, n20065, n20067, n20070, n20071, n20073, n20075, n20076, n20078, n20079, n20080, n20081, n20083, n20084, n20085, n20086, n20088, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20100, n20101, n20102, n20103, n20104, n20106, n20107, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20120, n20121, n20122, n20124, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20136, n20137, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20155, n20156, n20157, n20159, n20160, n20161, n20162, n20163, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20187, n20188, n20193, n20194, n20195, n20196, n20198, n20200, n20201, n20202, n20204, n20205, n20206, n20207, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20271, n20272, n20273, n20274, n20275, n20276, n20280, n20282, n20283, n20285, n20288, n20289, n20290, n20293, n20294, n20296, n20297, n20298, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20310, n20311, n20312, n20313, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20355, n20356, n20357, n20358, n20361, n20362, n20363, n20364, n20365, n20366, n20368, n20370, n20371, n20372, n20373, n20374, n20375, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20395, n20397, n20398, n20399, n20400, n20401, n20402, n20405, n20406, n20410, n20412, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20423, n20424, n20426, n20427, n20428, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20456, n20457, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20480, n20481, n20482, n20483, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20494, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20509, n20510, n20511, n20512, n20513, n20514, n20516, n20517, n20518, n20519, n20520, n20521, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20535, n20537, n20538, n20539, n20540, n20542, n20543, n20544, n20546, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20587, n20589, n20590, n20591, n20592, n20593, n20595, n20596, n20597, n20599, n20600, n20603, n20605, n20608, n20609, n20611, n20612, n20614, n20615, n20616, n20617, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20639, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20651, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20662, n20664, n20665, n20666, n20667, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20681, n20682, n20683, n20684, n20686, n20687, n20688, n20689, n20690, n20691, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20704, n20705, n20706, n20707, n20708, n20709, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20745, n20746, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20772, n20774, n20775, n20777, n20778, n20779, n20780, n20781, n20782, n20784, n20785, n20786, n20788, n20789, n20790, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20800, n20801, n20802, n20804, n20805, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20817, n20819, n20820, n20821, n20822, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20865, n20866, n20867, n20868, n20869, n20871, n20872, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20889, n20890, n20891, n20892, n20894, n20895, n20896, n20897, n20898, n20899, n20901, n20903, n20904, n20905, n20907, n20908, n20909, n20910, n20912, n20913, n20914, n20915, n20917, n20918, n20919, n20920, n20922, n20923, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20934, n20936, n20937, n20939, n20940, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20953, n20954, n20955, n20956, n20957, n20959, n20960, n20961, n20962, n20964, n20965, n20966, n20967, n20968, n20969, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21020, n21021, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21039, n21040, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21117, n21118, n21120, n21121, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21135, n21136, n21137, n21138, n21139, n21141, n21142, n21143, n21144, n21146, n21147, n21148, n21149, n21151, n21152, n21153, n21154, n21155, n21156, n21158, n21159, n21160, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21204, n21205, n21207, n21208, n21209, n21210, n21212, n21215, n21216, n21218, n21220, n21221, n21222, n21223, n21224, n21225, n21229, n21230, n21232, n21233, n21234, n21236, n21237, n21239, n21240, n21242, n21243, n21244, n21245, n21246, n21247, n21249, n21250, n21253, n21255, n21256, n21258, n21259, n21260, n21262, n21263, n21265, n21266, n21267, n21268, n21269, n21271, n21272, n21273, n21275, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21286, n21288, n21289, n21290, n21293, n21294, n21295, n21297, n21298, n21299, n21300, n21301, n21303, n21305, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21317, n21318, n21319, n21320, n21321, n21322, n21324, n21326, n21328, n21329, n21335, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21351, n21353, n21355, n21358, n21359, n21360, n21361, n21363, n21364, n21365, n21366, n21367, n21369, n21370, n21373, n21374, n21375, n21376, n21378, n21379, n21380, n21381, n21383, n21384, n21385, n21387, n21389, n21390, n21391, n21392, n21393, n21394, n21396, n21398, n21400, n21401, n21403, n21405, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21417, n21418, n21419, n21420, n21422, n21423, n21424, n21425, n21427, n21428, n21429, n21430, n21431, n21434, n21435, n21436, n21437, n21439, n21440, n21441, n21442, n21443, n21444, n21446, n21447, n21448, n21449, n21451, n21453, n21454, n21455, n21456, n21458, n21460, n21461, n21462, n21463, n21464, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21482, n21484, n21486, n21487, n21488, n21489, n21490, n21492, n21493, n21494, n21495, n21496, n21497, n21499, n21500, n21501, n21502, n21504, n21505, n21506, n21507, n21508, n21510, n21511, n21512, n21513, n21514, n21515, n21517, n21519, n21520, n21522, n21524, n21525, n21526, n21528, n21529, n21531, n21532, n21533, n21534, n21535, n21536, n21539, n21541, n21542, n21543, n21544, n21545, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21556, n21557, n21558, n21559, n21560, n21563, n21564, n21565, n21568, n21570, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21583, n21587, n21588, n21589, n21592, n21593, n21594, n21595, n21596, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21608, n21612, n21614, n21615, n21616, n21618, n21619, n21620, n21621, n21623, n21625, n21626, n21627, n21628, n21630, n21632, n21633, n21634, n21635, n21638, n21639, n21640, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21670, n21671, n21673, n21674, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21689, n21690, n21691, n21693, n21695, n21696, n21697, n21699, n21700, n21701, n21702, n21703, n21704, n21706, n21707, n21708, n21709, n21710, n21711, n21713, n21714, n21716, n21718, n21720, n21722, n21723, n21724, n21725, n21726, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21740, n21743, n21744, n21747, n21748, n21749, n21750, n21751, n21752, n21754, n21755, n21756, n21757, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21771, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21782, n21783, n21784, n21785, n21787, n21789, n21790, n21791, n21792, n21793, n21794, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21834, n21836, n21837, n21838, n21839, n21840, n21841, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21853, n21854, n21855, n21856, n21858, n21859, n21861, n21863, n21865, n21866, n21867, n21870, n21872, n21873, n21874, n21875, n21877, n21878, n21879, n21880, n21881, n21883, n21884, n21886, n21887, n21888, n21890, n21892, n21893, n21894, n21895, n21896, n21897, n21899, n21900, n21901, n21903, n21904, n21905, n21906, n21907, n21910, n21911, n21912, n21913, n21915, n21917, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21931, n21932, n21933, n21934, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21955, n21956, n21960, n21961, n21962, n21963, n21965, n21967, n21968, n21969, n21970, n21972, n21973, n21974, n21975, n21976, n21977, n21979, n21980, n21981, n21984, n21985, n21986, n21988, n21990, n21992, n21993, n21997, n22000, n22001, n22002, n22004, n22005, n22006, n22007, n22009, n22010, n22011, n22012, n22013, n22015, n22016, n22017, n22020, n22021, n22022, n22025, n22027, n22028, n22030, n22031, n22033, n22034, n22035, n22036, n22038, n22039, n22041, n22042, n22044, n22045, n22046, n22047, n22048, n22050, n22051, n22054, n22055, n22056, n22057, n22061, n22062, n22063, n22065, n22072, n22074, n22075, n22078, n22079, n22082, n22083, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22101, n22103, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22118, n22119, n22120, n22122, n22124, n22125, n22127, n22128, n22129, n22130, n22131, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22141, n22143, n22144, n22146, n22148, n22149, n22151, n22152, n22153, n22154, n22155, n22156, n22158, n22159, n22160, n22162, n22163, n22164, n22165, n22166, n22168, n22169, n22170, n22171, n22172, n22174, n22175, n22176, n22178, n22179, n22180, n22181, n22182, n22184, n22187, n22189, n22190, n22192, n22193, n22194, n22195, n22196, n22198, n22200, n22201, n22202, n22203, n22205, n22207, n22208, n22209, n22210, n22211, n22212, n22214, n22216, n22219, n22220, n22224, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22236, n22238, n22239, n22242, n22245, n22246, n22247, n22250, n22252, n22253, n22254, n22255, n22256, n22258, n22259, n22260, n22261, n22264, n22265, n22267, n22268, n22269, n22270, n22271, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22285, n22286, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22304, n22305, n22306, n22308, n22309, n22310, n22313, n22314, n22316, n22318, n22319, n22320, n22321, n22322, n22323, n22325, n22326, n22328, n22331, n22333, n22335, n22336, n22337, n22338, n22339, n22345, n22346, n22347, n22348, n22349, n22351, n22352, n22353, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22364, n22366, n22367, n22369, n22370, n22371, n22373, n22374, n22375, n22376, n22378, n22379, n22381, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22392, n22393, n22394, n22395, n22396, n22399, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22421, n22422, n22423, n22425, n22426, n22427, n22428, n22429, n22431, n22433, n22434, n22436, n22437, n22438, n22441, n22442, n22443, n22444, n22445, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22455, n22456, n22457, n22458, n22459, n22461, n22462, n22463, n22464, n22465, n22466, n22468, n22469, n22471, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22491, n22492, n22493, n22494, n22496, n22497, n22499, n22500, n22501, n22502, n22504, n22505, n22506, n22507, n22508, n22509, n22513, n22514, n22515, n22518, n22519, n22522, n22524, n22525, n22526, n22527, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22538, n22539, n22540, n22542, n22543, n22544, n22545, n22546, n22548, n22550, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22562, n22564, n22565, n22566, n22567, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22590, n22591, n22592, n22593, n22594, n22596, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22619, n22620, n22623, n22624, n22625, n22626, n22627, n22628, n22630, n22632, n22633, n22635, n22636, n22637, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22649, n22651, n22652, n22653, n22654, n22655, n22657, n22658, n22660, n22661, n22662, n22663, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22678, n22679, n22680, n22681, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22695, n22696, n22697, n22698, n22700, n22701, n22702, n22703, n22707, n22708, n22710, n22711, n22712, n22713, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22725, n22726, n22728, n22729, n22731, n22732, n22733, n22734, n22735, n22736, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22762, n22763, n22765, n22766, n22767, n22768, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22781, n22784, n22785, n22786, n22787, n22788, n22789, n22791, n22793, n22795, n22796, n22798, n22799, n22800, n22801, n22802, n22803, n22805, n22807, n22808, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22820, n22825, n22826, n22828, n22830, n22832, n22833, n22835, n22836, n22837, n22838, n22839, n22841, n22843, n22844, n22845, n22847, n22848, n22849, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22874, n22875, n22877, n22878, n22879, n22881, n22882, n22883, n22885, n22886, n22887, n22889, n22890, n22891, n22892, n22894, n22896, n22897, n22898, n22899, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22912, n22913, n22915, n22917, n22919, n22921, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22935, n22936, n22937, n22938, n22939, n22940, n22943, n22944, n22945, n22946, n22948, n22949, n22950, n22952, n22953, n22954, n22956, n22957, n22958, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22979, n22981, n22982, n22983, n22985, n22986, n22987, n22988, n22989, n22990, n22992, n22993, n22995, n22996, n22999, n23002, n23003, n23004, n23005, n23006, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23020, n23021, n23022, n23023, n23024, n23025, n23027, n23030, n23031, n23033, n23034, n23035, n23036, n23037, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23055, n23060, n23061, n23062, n23063, n23065, n23066, n23067, n23069, n23070, n23071, n23073, n23074, n23075, n23077, n23078, n23079, n23080, n23082, n23083, n23084, n23085, n23088, n23089, n23091, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23113, n23115, n23118, n23119, n23120, n23122, n23123, n23124, n23125, n23127, n23128, n23130, n23131, n23132, n23134, n23136, n23138, n23139, n23140, n23143, n23144, n23145, n23146, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23158, n23160, n23161, n23162, n23163, n23164, n23166, n23167, n23168, n23169, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23187, n23189, n23190, n23191, n23192, n23193, n23195, n23200, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23215, n23216, n23219, n23220, n23226, n23227, n23229, n23230, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23242, n23243, n23248, n23249, n23250, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23260, n23263, n23264, n23265, n23266, n23267, n23268, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23278, n23279, n23281, n23282, n23284, n23285, n23286, n23288, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23298, n23299, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23313, n23314, n23317, n23318, n23319, n23321, n23322, n23323, n23325, n23326, n23327, n23328, n23329, n23330, n23332, n23333, n23334, n23335, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23350, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23360, n23361, n23362, n23363, n23364, n23368, n23371, n23372, n23373, n23375, n23377, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23393, n23394, n23396, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23407, n23408, n23409, n23410, n23411, n23412, n23414, n23416, n23417, n23418, n23419, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23434, n23435, n23436, n23437, n23438, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23469, n23470, n23471, n23472, n23473, n23474, n23476, n23477, n23479, n23480, n23483, n23484, n23485, n23487, n23488, n23490, n23491, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23507, n23509, n23510, n23511, n23512, n23513, n23514, n23516, n23518, n23519, n23520, n23523, n23524, n23525, n23526, n23527, n23529, n23530, n23531, n23532, n23533, n23534, n23536, n23538, n23539, n23541, n23542, n23543, n23544, n23545, n23546, n23548, n23549, n23550, n23551, n23552, n23553, n23555, n23556, n23557, n23561, n23562, n23564, n23565, n23566, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23576, n23577, n23578, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23589, n23591, n23593, n23595, n23596, n23598, n23599, n23601, n23603, n23604, n23605, n23606, n23608, n23609, n23612, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23631, n23632, n23633, n23635, n23637, n23638, n23639, n23640, n23642, n23643, n23644, n23645, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23657, n23658, n23659, n23662, n23663, n23664, n23665, n23666, n23668, n23669, n23670, n23672, n23673, n23674, n23676, n23677, n23678, n23679, n23681, n23682, n23683, n23684, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23694, n23695, n23696, n23697, n23698, n23703, n23704, n23706, n23707, n23709, n23710, n23711, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23733, n23734, n23735, n23736, n23737, n23740, n23741, n23742, n23743, n23744, n23745, n23747, n23748, n23750, n23751, n23752, n23753, n23754, n23756, n23757, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23773, n23775, n23776, n23777, n23779, n23780, n23781, n23782, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23792, n23793, n23794, n23796, n23797, n23798, n23799, n23801, n23802, n23804, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23816, n23818, n23820, n23821, n23822, n23823, n23825, n23826, n23827, n23828, n23829, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23849, n23850, n23851, n23854, n23855, n23856, n23857, n23859, n23860, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23871, n23873, n23875, n23876, n23877, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23890, n23892, n23893, n23895, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23906, n23907, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23923, n23924, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23943, n23945, n23946, n23948, n23949, n23950, n23952, n23953, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23964, n23965, n23966, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23976, n23977, n23979, n23980, n23982, n23984, n23985, n23986, n23987, n23989, n23990, n23992, n23993, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24025, n24026, n24029, n24030, n24031, n24032, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24042, n24044, n24045, n24046, n24048, n24049, n24050, n24051, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24063, n24064, n24067, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24082, n24083, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24093, n24094, n24095, n24096, n24099, n24100, n24101, n24102, n24103, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24116, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24132, n24135, n24136, n24141, n24142, n24145, n24146, n24147, n24148, n24149, n24150, n24152, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24163, n24165, n24166, n24167, n24169, n24170, n24171, n24174, n24175, n24176, n24177, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24189, n24190, n24191, n24193, n24194, n24195, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24215, n24216, n24217, n24218, n24219, n24220, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24231, n24232, n24233, n24235, n24236, n24237, n24239, n24240, n24242, n24243, n24245, n24247, n24248, n24250, n24251, n24252, n24253, n24255, n24256, n24257, n24258, n24260, n24261, n24262, n24263, n24264, n24265, n24267, n24268, n24269, n24270, n24271, n24272, n24275, n24276, n24278, n24280, n24281, n24282, n24284, n24285, n24287, n24288, n24289, n24291, n24292, n24293, n24294, n24296, n24300, n24301, n24303, n24304, n24306, n24307, n24308, n24310, n24311, n24313, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24326, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24343, n24344, n24345, n24346, n24348, n24349, n24350, n24351, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24361, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24373, n24375, n24376, n24377, n24378, n24379, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24394, n24395, n24396, n24397, n24398, n24400, n24401, n24402, n24405, n24406, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24421, n24422, n24423, n24424, n24425, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24437, n24438, n24439, n24441, n24442, n24444, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24455, n24456, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24467, n24469, n24470, n24471, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24484, n24485, n24487, n24488, n24490, n24491, n24492, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24507, n24508, n24509, n24510, n24511, n24513, n24514, n24517, n24518, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24528, n24529, n24532, n24533, n24536, n24537, n24538, n24540, n24541, n24542, n24543, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24553, n24554, n24556, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24575, n24576, n24577, n24579, n24580, n24581, n24583, n24585, n24586, n24587, n24588, n24589, n24591, n24594, n24595, n24596, n24597, n24600, n24601, n24602, n24604, n24605, n24606, n24608, n24610, n24611, n24612, n24614, n24616, n24617, n24618, n24620, n24623, n24625, n24626, n24627, n24629, n24630, n24631, n24632, n24634, n24635, n24636, n24637, n24639, n24640, n24641, n24643, n24645, n24648, n24649, n24652, n24653, n24654, n24655, n24656, n24658, n24659, n24660, n24661, n24662, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24707, n24708, n24709, n24710, n24712, n24713, n24714, n24716, n24718, n24719, n24720, n24721, n24722, n24723, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24733, n24734, n24735, n24737, n24738, n24740, n24741, n24743, n24744, n24745, n24746, n24748, n24750, n24751, n24753, n24754, n24755, n24756, n24758, n24759, n24760, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24778, n24779, n24780, n24781, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24808, n24809, n24810, n24811, n24812, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24825, n24827, n24828, n24831, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24841, n24842, n24843, n24845, n24846, n24849, n24850, n24851, n24852, n24853, n24854, n24857, n24860, n24861, n24862, n24863, n24865, n24866, n24867, n24868, n24873, n24874, n24875, n24876, n24878, n24879, n24880, n24881, n24882, n24883, n24886, n24888, n24889, n24891, n24892, n24893, n24897, n24898, n24899, n24900, n24901, n24902, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24918, n24919, n24920, n24921, n24923, n24924, n24925, n24926, n24928, n24930, n24931, n24932, n24934, n24935, n24936, n24940, n24942, n24944, n24947, n24948, n24949, n24951, n24952, n24953, n24955, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24965, n24966, n24967, n24970, n24971, n24972, n24974, n24976, n24977, n24980, n24981, n24982, n24984, n24985, n24986, n24987, n24988, n24989, n24991, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25004, n25005, n25007, n25008, n25009, n25010, n25011, n25013, n25014, n25015, n25018, n25019, n25020, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25043, n25044, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25055, n25056, n25058, n25059, n25060, n25061, n25063, n25065, n25068, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25089, n25090, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25116, n25117, n25119, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25133, n25134, n25137, n25138, n25139, n25140, n25141, n25142, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25159, n25160, n25161, n25162, n25163, n25164, n25166, n25167, n25168, n25169, n25173, n25174, n25175, n25176, n25177, n25178, n25180, n25182, n25183, n25184, n25185, n25187, n25188, n25189, n25191, n25194, n25195, n25196, n25197, n25198, n25201, n25202, n25203, n25204, n25205, n25206, n25208, n25209, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25230, n25231, n25232, n25234, n25236, n25241, n25242, n25243, n25244, n25245, n25246, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25258, n25259, n25261, n25262, n25263, n25264, n25269, n25270, n25271, n25273, n25274, n25275, n25276, n25277, n25279, n25280, n25283, n25284, n25286, n25287, n25289, n25290, n25291, n25292, n25293, n25294, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25311, n25312, n25314, n25315, n25317, n25320, n25321, n25322, n25323, n25325, n25326, n25327, n25328, n25329, n25331, n25332, n25333, n25334, n25335, n25336, n25338, n25341, n25342, n25343, n25344, n25346, n25348, n25349, n25351, n25352, n25353, n25354, n25355, n25357, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25369, n25370, n25371, n25372, n25374, n25377, n25378, n25379, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25391, n25392, n25393, n25394, n25395, n25398, n25402, n25403, n25404, n25405, n25406, n25408, n25409, n25410, n25411, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25421, n25422, n25423, n25424, n25427, n25428, n25432, n25433, n25435, n25436, n25438, n25440, n25441, n25442, n25444, n25445, n25446, n25447, n25449, n25450, n25453, n25454, n25455, n25457, n25459, n25460, n25462, n25463, n25465, n25466, n25467, n25469, n25471, n25474, n25475, n25476, n25477, n25478, n25479, n25481, n25482, n25484, n25485, n25486, n25487, n25488, n25490, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25502, n25503, n25504, n25507, n25508, n25509, n25510, n25511, n25513, n25515, n25516, n25517, n25518, n25519, n25522, n25524, n25525, n25526, n25528, n25529, n25531, n25532, n25533, n25534, n25536, n25537, n25539, n25544, n25546, n25547, n25548, n25550, n25551, n25553, n25555, n25557, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25579, n25580, n25581, n25582, n25583, n25584, n25586, n25588, n25590, n25591, n25592, n25593, n25594, n25597, n25598, n25600, n25601, n25602, n25603, n25604, n25605, n25607, n25608, n25613, n25614, n25615, n25619, n25621, n25624, n25625, n25626, n25627, n25630, n25631, n25632, n25633, n25635, n25636, n25638, n25639, n25640, n25641, n25642, n25644, n25649, n25650, n25651, n25653, n25654, n25656, n25657, n25658, n25660, n25661, n25662, n25663, n25664, n25665, n25668, n25669, n25671, n25672, n25676, n25677, n25679, n25680, n25681, n25683, n25685, n25689, n25691, n25692, n25693, n25694, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25706, n25707, n25708, n25710, n25712, n25716, n25717, n25718, n25719, n25720, n25721, n25723, n25725, n25728, n25730, n25731, n25732, n25734, n25738, n25741, n25743, n25745, n25747, n25748, n25750, n25751, n25753, n25754, n25756, n25758, n25759, n25760, n25764, n25765, n25766, n25768, n25771, n25773, n25774, n25775, n25776, n25777, n25778, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25792, n25794, n25795, n25796, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25808, n25810, n25813, n25814, n25815, n25816, n25817, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25829, n25830, n25831, n25832, n25833, n25834, n25836, n25837, n25839, n25841, n25842, n25844, n25845, n25846, n25847, n25849, n25850, n25852, n25856, n25857, n25858, n25860, n25862, n25863, n25864, n25865, n25866, n25868, n25869, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25889, n25890, n25891, n25893, n25894, n25895, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25909, n25911, n25912, n25915, n25916, n25917, n25919, n25920, n25921, n25922, n25924, n25925, n25926, n25927, n25929, n25930, n25931, n25932, n25933, n25934, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25945, n25947, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25969, n25973, n25974, n25975, n25977, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26001, n26003, n26004, n26007, n26008, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26021, n26022, n26025, n26026, n26027, n26030, n26031, n26033, n26035, n26036, n26037, n26038, n26040, n26041, n26043, n26044, n26045, n26046, n26047, n26049, n26051, n26054, n26057, n26059, n26060, n26061, n26063, n26064, n26066, n26067, n26068, n26069, n26070, n26071, n26074, n26075, n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26092, n26093, n26095, n26098, n26099, n26101, n26102, n26105, n26107, n26108, n26109, n26110, n26111, n26114, n26115, n26117, n26119, n26121, n26122, n26125, n26126, n26127, n26128, n26129, n26130, n26133, n26135, n26136, n26140, n26142, n26143, n26144, n26145, n26147, n26148, n26149, n26150, n26151, n26155, n26156, n26157, n26158, n26159, n26160, n26164, n26165, n26167, n26168, n26169, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26182, n26184, n26185, n26186, n26187, n26190, n26193, n26194, n26195, n26196, n26198, n26202, n26203, n26205, n26207, n26209, n26210, n26211, n26212, n26213, n26216, n26217, n26218, n26220, n26222, n26224, n26225, n26226, n26229, n26232, n26233, n26239, n26240, n26241, n26242, n26243, n26245, n26248, n26250, n26252, n26253, n26255, n26256, n26257, n26258, n26260, n26262, n26263, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26275, n26278, n26280, n26281, n26282, n26283, n26287, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26299, n26300, n26301, n26302, n26303, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26318, n26319, n26320, n26321, n26323, n26324, n26325, n26327, n26328, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26338, n26340, n26341, n26342, n26343, n26344, n26345, n26348, n26350, n26352, n26355, n26356, n26357, n26360, n26362, n26364, n26366, n26368, n26370, n26371, n26373, n26376, n26377, n26379, n26380, n26381, n26382, n26383, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26398, n26401, n26404, n26405, n26407, n26411, n26412, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26430, n26431, n26433, n26437, n26438, n26439, n26441, n26443, n26444, n26445, n26447, n26448, n26449, n26450, n26451, n26455, n26456, n26457, n26458, n26459, n26460, n26462, n26463, n26464, n26465, n26466, n26468, n26469, n26471, n26472, n26473, n26474, n26476, n26479, n26481, n26482, n26484, n26485, n26486, n26487, n26488, n26489, n26491, n26493, n26495, n26497, n26498, n26501, n26502, n26504, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26516, n26517, n26519, n26520, n26525, n26526, n26527, n26530, n26532, n26533, n26536, n26538, n26539, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26552, n26554, n26555, n26556, n26557, n26559, n26560, n26561, n26564, n26565, n26566, n26567, n26568, n26569, n26572, n26576, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26604, n26605, n26606, n26607, n26608, n26610, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26621, n26622, n26623, n26624, n26626, n26627, n26628, n26632, n26633, n26634, n26635, n26636, n26638, n26639, n26641, n26642, n26643, n26645, n26646, n26647, n26648, n26650, n26651, n26652, n26653, n26654, n26655, n26657, n26658, n26661, n26663, n26664, n26665, n26666, n26667, n26669, n26670, n26671, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26693, n26694, n26695, n26696, n26697, n26700, n26703, n26704, n26707, n26708, n26709, n26711, n26713, n26715, n26716, n26719, n26720, n26722, n26723, n26724, n26725, n26727, n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26737, n26738, n26740, n26742, n26744, n26746, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26758, n26759, n26761, n26762, n26763, n26764, n26767, n26768, n26769, n26770, n26772, n26773, n26774, n26775, n26778, n26779, n26780, n26782, n26783, n26786, n26788, n26791, n26792, n26793, n26795, n26796, n26797, n26801, n26802, n26804, n26805, n26806, n26807, n26808, n26810, n26811, n26812, n26813, n26814, n26815, n26817, n26818, n26819, n26824, n26826, n26827, n26829, n26831, n26833, n26834, n26835, n26836, n26838, n26839, n26840, n26841, n26842, n26843, n26846, n26847, n26848, n26849, n26850, n26852, n26853, n26856, n26858, n26859, n26860, n26861, n26862, n26863, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26881, n26882, n26883, n26884, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26897, n26898, n26900, n26901, n26902, n26906, n26908, n26910, n26911, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26922, n26925, n26926, n26927, n26928, n26929, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26941, n26943, n26944, n26946, n26947, n26948, n26949, n26951, n26952, n26953, n26956, n26958, n26959, n26960, n26962, n26963, n26965, n26966, n26967, n26968, n26969, n26970, n26972, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26985, n26990, n26994, n26995, n26996, n26998, n27000, n27003, n27005, n27006, n27007, n27008, n27009, n27011, n27012, n27015, n27017, n27018, n27019, n27020, n27022, n27026, n27028, n27029, n27030, n27031, n27032, n27033, n27037, n27039, n27043, n27044, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27059, n27060, n27062, n27064, n27066, n27067, n27068, n27069, n27070, n27072, n27076, n27077, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27089, n27092, n27093, n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27115, n27116, n27117, n27119, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27131, n27132, n27137, n27138, n27139, n27140, n27141, n27143, n27144, n27145, n27146, n27147, n27149, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27160, n27161, n27162, n27163, n27164, n27165, n27167, n27168, n27170, n27171, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27181, n27182, n27183, n27184, n27185, n27186, n27190, n27191, n27196, n27197, n27199, n27201, n27205, n27206, n27207, n27209, n27210, n27211, n27213, n27214, n27215, n27217, n27218, n27219, n27220, n27221, n27223, n27225, n27226, n27229, n27231, n27232, n27234, n27235, n27236, n27237, n27239, n27240, n27241, n27245, n27247, n27249, n27250, n27252, n27255, n27256, n27257, n27259, n27260, n27261, n27262, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27274, n27275, n27276, n27278, n27279, n27280, n27281, n27282, n27283, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27293, n27294, n27296, n27297, n27298, n27300, n27301, n27303, n27304, n27305, n27308, n27309, n27310, n27314, n27316, n27317, n27318, n27319, n27320, n27321, n27324, n27325, n27327, n27328, n27329, n27331, n27332, n27334, n27336, n27337, n27339, n27340, n27342, n27346, n27347, n27349, n27353, n27354, n27355, n27357, n27358, n27360, n27361, n27362, n27365, n27366, n27368, n27369, n27370, n27373, n27374, n27376, n27377, n27378, n27379, n27380, n27382, n27384, n27387, n27389, n27391, n27392, n27393, n27394, n27396, n27397, n27399, n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27411, n27412, n27413, n27416, n27417, n27419, n27420, n27421, n27422, n27423, n27425, n27426, n27427, n27428, n27429, n27431, n27433, n27434, n27436, n27438, n27439, n27440, n27442, n27444, n27445, n27448, n27449, n27452, n27453, n27454, n27455, n27456, n27459, n27462, n27463, n27464, n27465, n27467, n27472, n27473, n27474, n27477, n27478, n27479, n27480, n27482, n27483, n27484, n27486, n27488, n27489, n27492, n27496, n27498, n27499, n27500, n27501, n27503, n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27540, n27541, n27543, n27544, n27545, n27546, n27547, n27549, n27552, n27553, n27554, n27556, n27557, n27558, n27560, n27561, n27562, n27564, n27565, n27566, n27567, n27571, n27572, n27573, n27574, n27575, n27577, n27578, n27581, n27582, n27583, n27584, n27585, n27588, n27589, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27615, n27616, n27617, n27619, n27620, n27621, n27623, n27624, n27625, n27631, n27634, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27651, n27652, n27656, n27657, n27658, n27659, n27661, n27663, n27666, n27667, n27668, n27669, n27670, n27673, n27674, n27677, n27678, n27679, n27680, n27683, n27684, n27687, n27688, n27690, n27691, n27692, n27694, n27695, n27696, n27697, n27698, n27700, n27702, n27703, n27705, n27706, n27707, n27709, n27710, n27712, n27714, n27715, n27717, n27718, n27723, n27724, n27725, n27726, n27727, n27730, n27732, n27734, n27736, n27737, n27739, n27740, n27741, n27742, n27743, n27745, n27746, n27747, n27749, n27750, n27753, n27754, n27755, n27758, n27759, n27760, n27761, n27763, n27765, n27766, n27767, n27768, n27771, n27772, n27773, n27774, n27776, n27777, n27779, n27781, n27782, n27784, n27785, n27791, n27793, n27795, n27796, n27797, n27799, n27800, n27801, n27802, n27803, n27806, n27808, n27810, n27812, n27814, n27815, n27816, n27817, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27831, n27832, n27834, n27836, n27838, n27839, n27840, n27843, n27845, n27846, n27847, n27851, n27852, n27853, n27855, n27857, n27858, n27859, n27860, n27862, n27863, n27864, n27865, n27866, n27867, n27869, n27870, n27871, n27872, n27874, n27875, n27876, n27877, n27878, n27880, n27881, n27882, n27884, n27885, n27888, n27889, n27891, n27892, n27893, n27895, n27897, n27898, n27899, n27901, n27902, n27904, n27905, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27916, n27917, n27919, n27920, n27921, n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27933, n27934, n27936, n27937, n27938, n27939, n27940, n27943, n27945, n27946, n27948, n27950, n27951, n27952, n27953, n27956, n27957, n27960, n27961, n27962, n27963, n27964, n27966, n27968, n27969, n27970, n27971, n27972, n27973, n27975, n27978, n27979, n27980, n27981, n27982, n27983, n27985, n27987, n27989, n27991, n27992, n27993, n27995, n27996, n27997, n27998, n27999, n28002, n28004, n28006, n28008, n28009, n28010, n28011, n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28027, n28028, n28029, n28031, n28034, n28036, n28037, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28049, n28050, n28052, n28053, n28055, n28056, n28057, n28058, n28060, n28061, n28063, n28064, n28066, n28069, n28070, n28072, n28076, n28077, n28078, n28079, n28081, n28082, n28083, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28118, n28121, n28122, n28124, n28125, n28126, n28127, n28132, n28133, n28135, n28136, n28137, n28138, n28139, n28141, n28142, n28143, n28144, n28146, n28147, n28148, n28150, n28151, n28154, n28156, n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28169, n28170, n28171, n28172, n28174, n28176, n28177, n28178, n28179, n28182, n28183, n28185, n28186, n28190, n28191, n28192, n28193, n28194, n28195, n28197, n28198, n28199, n28201, n28202, n28203, n28204, n28205, n28206, n28208, n28211, n28214, n28215, n28217, n28218, n28219, n28220, n28222, n28226, n28227, n28229, n28232, n28233, n28234, n28235, n28237, n28238, n28241, n28242, n28244, n28245, n28246, n28248, n28250, n28252, n28253, n28254, n28256, n28257, n28258, n28260, n28264, n28265, n28267, n28269, n28270, n28271, n28272, n28273, n28276, n28277, n28279, n28282, n28284, n28287, n28289, n28290, n28294, n28295, n28297, n28298, n28299, n28301, n28302, n28303, n28304, n28305, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28317, n28318, n28320, n28321, n28324, n28325, n28326, n28328, n28329, n28334, n28335, n28336, n28339, n28342, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28352, n28353, n28354, n28356, n28358, n28359, n28361, n28363, n28364, n28365, n28368, n28371, n28372, n28374, n28375, n28379, n28380, n28381, n28382, n28384, n28385, n28386, n28387, n28389, n28390, n28392, n28393, n28396, n28397, n28399, n28401, n28403, n28404, n28405, n28406, n28408, n28409, n28410, n28411, n28412, n28417, n28418, n28419, n28421, n28422, n28423, n28426, n28427, n28429, n28430, n28431, n28432, n28434, n28435, n28436, n28437, n28439, n28440, n28441, n28443, n28444, n28445, n28446, n28448, n28450, n28451, n28452, n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28463, n28465, n28466, n28467, n28469, n28471, n28472, n28475, n28476, n28477, n28478, n28479, n28481, n28483, n28485, n28486, n28487, n28488, n28490, n28491, n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28503, n28506, n28507, n28508, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28520, n28521, n28522, n28523, n28526, n28528, n28529, n28531, n28532, n28537, n28538, n28540, n28544, n28545, n28546, n28547, n28548, n28551, n28553, n28554, n28555, n28556, n28557, n28559, n28560, n28561, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28574, n28575, n28577, n28578, n28581, n28582, n28585, n28586, n28587, n28588, n28589, n28590, n28594, n28596, n28599, n28600, n28601, n28602, n28603, n28606, n28610, n28611, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28622, n28625, n28627, n28628, n28629, n28630, n28631, n28633, n28634, n28635, n28636, n28637, n28639, n28640, n28642, n28643, n28644, n28645, n28646, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28659, n28660, n28662, n28663, n28664, n28665, n28667, n28668, n28669, n28673, n28674, n28675, n28677, n28678, n28679, n28680, n28681, n28682, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28695, n28697, n28698, n28699, n28701, n28702, n28703, n28704, n28705, n28706, n28708, n28709, n28710, n28711, n28712, n28714, n28716, n28717, n28718, n28719, n28720, n28721, n28724, n28726, n28727, n28729, n28730, n28731, n28732, n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28746, n28747, n28749, n28750, n28753, n28754, n28756, n28757, n28758, n28760, n28761, n28762, n28763, n28764, n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28776, n28777, n28779, n28781, n28782, n28783, n28785, n28786, n28787, n28788, n28789, n28793, n28794, n28795, n28796, n28797, n28798, n28801, n28803, n28804, n28805, n28807, n28808, n28809, n28810, n28813, n28815, n28817, n28819, n28820, n28821, n28822, n28823, n28825, n28828, n28831, n28832, n28833, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28850, n28854, n28855, n28856, n28857, n28859, n28860, n28861, n28864, n28865, n28867, n28868, n28870, n28871, n28873, n28874, n28876, n28877, n28878, n28880, n28882, n28884, n28885, n28886, n28888, n28889, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28901, n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28919, n28920, n28921, n28922, n28923, n28925, n28927, n28930, n28933, n28937, n28938, n28939, n28942, n28943, n28944, n28945, n28946, n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28956, n28957, n28958, n28959, n28960, n28962, n28963, n28964, n28965, n28966, n28968, n28969, n28970, n28973, n28974, n28975, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28986, n28987, n28988, n28989, n28990, n28991, n28993, n28995, n28996, n28997, n28998, n28999, n29000, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29018, n29019, n29021, n29022, n29024, n29025, n29026, n29027, n29028, n29030, n29031, n29032, n29033, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29043, n29044, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29055, n29058, n29061, n29063, n29064, n29065, n29066, n29069, n29071, n29072, n29075, n29078, n29079, n29082, n29083, n29084, n29085, n29087, n29088, n29089, n29090, n29091, n29093, n29094, n29097, n29098, n29099, n29100, n29101, n29102, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29113, n29114, n29116, n29117, n29118, n29119, n29120, n29122, n29125, n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29139, n29144, n29146, n29147, n29148, n29149, n29150, n29151, n29153, n29154, n29156, n29157, n29158, n29159, n29160, n29162, n29163, n29164, n29165, n29167, n29168, n29169, n29170, n29172, n29173, n29174, n29175, n29176, n29179, n29180, n29181, n29182, n29183, n29185, n29186, n29188, n29190, n29191, n29193, n29195, n29196, n29197, n29198, n29201, n29205, n29207, n29208, n29210, n29211, n29212, n29214, n29216, n29217, n29219, n29221, n29222, n29223, n29225, n29226, n29227, n29228, n29230, n29231, n29232, n29233, n29235, n29236, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29253, n29254, n29255, n29257, n29259, n29260, n29262, n29263, n29264, n29265, n29266, n29270, n29271, n29272, n29274, n29275, n29276, n29278, n29279, n29280, n29281, n29282, n29284, n29285, n29286, n29287, n29289, n29292, n29293, n29294, n29295, n29296, n29298, n29299, n29300, n29304, n29305, n29308, n29309, n29310, n29311, n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29329, n29330, n29331, n29332, n29333, n29335, n29337, n29339, n29340, n29343, n29344, n29346, n29347, n29351, n29352, n29353, n29354, n29355, n29358, n29359, n29363, n29364, n29365, n29366, n29367, n29371, n29372, n29374, n29375, n29376, n29377, n29382, n29383, n29384, n29385, n29386, n29388, n29389, n29391, n29392, n29393, n29394, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29405, n29406, n29407, n29408, n29409, n29410, n29412, n29413, n29416, n29418, n29419, n29420, n29422, n29423, n29424, n29425, n29428, n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29449, n29450, n29451, n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29463, n29464, n29465, n29467, n29468, n29470, n29472, n29474, n29475, n29477, n29479, n29480, n29481, n29483, n29484, n29485, n29486, n29487, n29489, n29490, n29491, n29492, n29494, n29495, n29496, n29500, n29502, n29503, n29504, n29505, n29506, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29521, n29522, n29523, n29524, n29525, n29526, n29528, n29531, n29532, n29535, n29536, n29540, n29541, n29542, n29544, n29545, n29546, n29547, n29548, n29551, n29553, n29555, n29556, n29557, n29559, n29560, n29561, n29564, n29565, n29566, n29567, n29569, n29574, n29575, n29577, n29578, n29580, n29582, n29583, n29586, n29587, n29589, n29591, n29592, n29593, n29595, n29596, n29597, n29598, n29599, n29600, n29602, n29603, n29604, n29607, n29608, n29609, n29611, n29612, n29613, n29615, n29616, n29617, n29618, n29619, n29621, n29622, n29623, n29625, n29626, n29629, n29630, n29634, n29635, n29636, n29637, n29638, n29639, n29642, n29644, n29647, n29650, n29653, n29656, n29660, n29661, n29664, n29665, n29667, n29671, n29672, n29673, n29674, n29675, n29677, n29678, n29680, n29681, n29683, n29684, n29685, n29687, n29688, n29689, n29692, n29694, n29695, n29696, n29697, n29698, n29701, n29702, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29725, n29728, n29730, n29732, n29733, n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29743, n29744, n29745, n29749, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29761, n29762, n29763, n29766, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29780, n29781, n29782, n29783, n29784, n29788, n29790, n29791, n29792, n29793, n29797, n29799, n29800, n29801, n29803, n29805, n29806, n29807, n29809, n29810, n29814, n29815, n29818, n29819, n29821, n29823, n29824, n29826, n29827, n29828, n29830, n29831, n29832, n29834, n29835, n29838, n29839, n29841, n29842, n29844, n29847, n29848, n29851, n29854, n29856, n29858, n29859, n29860, n29861, n29862, n29864, n29865, n29867, n29868, n29869, n29870, n29871, n29872, n29877, n29880, n29881, n29882, n29883, n29884, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29895, n29896, n29897, n29898, n29900, n29902, n29903, n29904, n29905, n29906, n29908, n29909, n29910, n29911, n29912, n29914, n29915, n29916, n29917, n29919, n29920, n29921, n29922, n29924, n29929, n29930, n29932, n29933, n29936, n29937, n29938, n29939, n29940, n29941, n29943, n29945, n29949, n29950, n29951, n29954, n29958, n29961, n29962, n29963, n29964, n29967, n29968, n29970, n29971, n29973, n29974, n29977, n29978, n29979, n29982, n29983, n29985, n29986, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30010, n30011, n30013, n30014, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30028, n30029, n30030, n30032, n30033, n30037, n30038, n30039, n30040, n30041, n30043, n30047, n30048, n30049, n30051, n30052, n30053, n30054, n30055, n30056, n30058, n30061, n30062, n30063, n30065, n30067, n30068, n30069, n30071, n30072, n30073, n30074, n30075, n30076, n30078, n30081, n30082, n30083, n30086, n30087, n30088, n30089, n30090, n30092, n30094, n30095, n30099, n30100, n30101, n30103, n30106, n30107, n30112, n30113, n30114, n30115, n30117, n30120, n30121, n30122, n30125, n30126, n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30136, n30145, n30147, n30151, n30152, n30153, n30154, n30156, n30159, n30160, n30166, n30167, n30168, n30172, n30173, n30175, n30182, n30185, n30200, n30202, n30204, n30207, n30209, n30211, n30220, n30229, n30231, n30232, n30234, n30235, n30238, n30240, n30244, n30246, n30250, n30251, n30254, n30257, n30261, n30269, n30271, n30274, n30276, n30277, n30282, n30285, n30287, n30289, n30290, n30291, n30294, n30299, n30300, n30302, n30304, n30306, n30308, n30310, n30311, n30312, n30315, n30318, n30320, n30324, n30327, n30328, n30329, n30332, n30335, n30340, n30342, n30346, n30349, n30351, n30353, n30355, n30356, n30360, n30362, n30368, n30371, n30379, n30380, n30384, n30385, n30387, n30388, n30390, n30392, n30394, n30397, n30399, n30400, n30402, n30403, n30408, n30409, n30410, n30417, n30422, n30423, n30425, n30429, n30430, n30431, n30433, n30436, n30439, n30441, n30445, n30450, n30451, n30464, n30465, n30472, n30473, n30475, n30478, n30482, n30483, n30486, n30489, n30490, n30492, n30494, n30501, n30511, n30512, n30513, n30516, n30518, n30525, n30526, n30535, n30538, n30541, n30542, n30543, n30547, n30548, n30549, n30550, n30552, n30555, n30556, n30558, n30562, n30563, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30573, n30574, n30576, n30581, n30583, n30587, n30594, n30599, n30600, n30604, n30606, n30607, n30610, n30614, n30619, n30624, n30626, n30629, n30630, n30632, n30637, n30640, n30645, n30646, n30647, n30648, n30653, n30657, n30661, n30680, n30684, n30686, n30690, n30695, n30697, n30698, n30700, n30701, n30702, n30707, n30708, n30709, n30711, n30715, n30720, n30722, n30723, n30728, n30729, n30733, n30734, n30736, n30738, n30740, n30745, n30746, n30748, n30752, n30754, n30757, n30760, n30762, n30764, n30765, n30770, n30771, n30775, n30776, n30778, n30783, n30788, n30797, n30798, n30799, n30800, n30802, n30805, n30807, n30811, n30812, n30814, n30820, n30821, n30825, n30830, n30831, n30835, n30841, n30844, n30848, n30854, n30857, n30859, n30860, n30867, n30868, n30870, n30874, n30878, n30884, n30889, n30891, n30892, n30894, n30897, n30899, n30906, n30909, n30910, n30911, n30920, n30924, n30927, n30928, n30929, n30931, n30932, n30938, n30940, n30941, n30943, n30951, n30954, n30955, n30956, n30958, n30961, n30967, n30969, n30973, n30978, n30980, n30984, n30985, n30989, n30990, n30995, n30996, n30997, n31001, n31002, n31008, n31011, n31012, n31013, n31014, n31015, n31024, n31025, n31026, n31027, n31030, n31031, n31034, n31040, n31042, n31044, n31046, n31049, n31055, n31060, n31063, n31066, n31067, n31070, n31073, n31074, n31075, n31076, n31079, n31084, n31086, n31087, n31090, n31091, n31092, n31095, n31099, n31100, n31102, n31104, n31106, n31109, n31114, n31119, n31120, n31121, n31122, n31124, n31126, n31130, n31132, n31135, n31136, n31139, n31140, n31142, n31143, n31144, n31146, n31147, n31150, n31151, n31154, n31156, n31161, n31162, n31168, n31170, n31173, n31175, n31177, n31179, n31181, n31183, n31187, n31190, n31191, n31195, n31198, n31201, n31208, n31209, n31214, n31215, n31216, n31217, n31222, n31226, n31228, n31234, n31237, n31238, n31239, n31242, n31244, n31245, n31247, n31249, n31250, n31254, n31256, n31257, n31261, n31264, n31265, n31267, n31268, n31276, n31278, n31279, n31281, n31288, n31289, n31292, n31296, n31298, n31300, n31302, n31303, n31304, n31305, n31306, n31307, n31311, n31314, n31316, n31318, n31322, n31323, n31327, n31330, n31331, n31334, n31344, n31345, n31347, n31348, n31349, n31351, n31353, n31354, n31358, n31359, n31360, n31363, n31366, n31369, n31373, n31380, n31381, n31384, n31394, n31399, n31400, n31410, n31411, n31413, n31419, n31423, n31426, n31427, n31429, n31435, n31436, n31437, n31440, n31442, n31444, n31445, n31446, n31449, n31454, n31455, n31456, n31457, n31458, n31460, n31461, n31462, n31468, n31470, n31476, n31480, n31486, n31487, n31493, n31494, n31500, n31503, n31504, n31509, n31510, n31515, n31523, n31526, n31530, n31531, n31534, n31539, n31545, n31547, n31549, n31552, n31555, n31558, n31559, n31564, n31569, n31572, n31577, n31578, n31585, n31590, n31592, n31599, n31601, n31602, n31604, n31607, n31609, n31611, n31612, n31613, n31616, n31623, n31625, n31626, n31631, n31633, n31634, n31635, n31636, n31639, n31640, n31641, n31644, n31646, n31650, n31661, n31662, n31663, n31669, n31671, n31675, n31676, n31678, n31680, n31683, n31690, n31702, n31709, n31713, n31716, n31721, n31722, n31723, n31726, n31727, n31729, n31730, n31732, n31733, n31735, n31739, n31741, n31743, n31747, n31748, n31750, n31751, n31755, n31756, n31758, n31769, n31770, n31774, n31779, n31780, n31782, n31784, n31786, n31792, n31795, n31796, n31798, n31799, n31800, n31804, n31809, n31816, n31832, n31835, n31838, n31839, n31844, n31847, n31853, n31856, n31861, n31862, n31863, n31864, n31866, n31869, n31874, n31877, n31878, n31879, n31886, n31889, n31893, n31894, n31897, n31898, n31901, n31902, n31905, n31909, n31914, n31917, n31919, n31921, n31923, n31926, n31927, n31931, n31934, n31935, n31936, n31938, n31943, n31951, n31952, n31955, n31958, n31961, n31968, n31970, n31972, n31975, n31978, n31980, n31986, n31987, n31993, n31995, n31997, n32003, n32005, n32006, n32008, n32009, n32011, n32016, n32022, n32023, n32024, n32025, n32029, n32031, n32033, n32035, n32039, n32043, n32044, n32046, n32049, n32052, n32060, n32061, n32063, n32067, n32071, n32072, n32074, n32085, n32086, n32091, n32094, n32095, n32096, n32100, n32102, n32103, n32107, n32112, n32113, n32115, n32116, n32120, n32122, n32123, n32125, n32126, n32128, n32131, n32132, n32133, n32139, n32140, n32142, n32149, n32156, n32157, n32158, n32159, n32163, n32166, n32168, n32169, n32170, n32172, n32178, n32180, n32181, n32185, n32188, n32191, n32194, n32196, n32197, n32198, n32202, n32204, n32205, n32206, n32207, n32208, n32211, n32213, n32215, n32217, n32220, n32221, n32227, n32231, n32239, n32241, n32242, n32245, n32248, n32254, n32256, n32258, n32261, n32268, n32270, n32271, n32281, n32284, n32285, n32286, n32289, n32297, n32299, n32300, n32306, n32307, n32322, n32323, n32324, n32326, n32331, n32332, n32334, n32335, n32338, n32344, n32358, n32360, n32364, n32366, n32368, n32371, n32375, n32376, n32381, n32390, n32391, n32395, n32398, n32402, n32403, n32413, n32414, n32415, n32417, n32423, n32436, n32443, n32450, n32452, n32453, n32457, n32458, n32462, n32463, n32467, n32468, n32470, n32477, n32478, n32479, n32484, n32485, n32486, n32487, n32488, n32493, n32495, n32497, n32499, n32503, n32504, n32509, n32510, n32512, n32515, n32516, n32518, n32520, n32523, n32524, n32529, n32530, n32533, n32534, n32536, n32537, n32538, n32541, n32545, n32546, n32549, n32551, n32555, n32556, n32561, n32566, n32569, n32571, n32572, n32574, n32578, n32580, n32588, n32591, n32594, n32596, n32601, n32605, n32609, n32611, n32612, n32614, n32620, n32627, n32630, n32632, n32636, n32646, n32647, n32648, n32649, n32651, n32659, n32660, n32664, n32672, n32675, n32680, n32681, n32683, n32684, n32687, n32688, n32692, n32697, n32699, n32701, n32708, n32711, n32715, n32717, n32721, n32724, n32727, n32729, n32734, n32739, n32746, n32751, n32753, n32757, n32761, n32766, n32767, n32768, n32775, n32776, n32780, n32783, n32791, n32803, n32805, n32806, n32808, n32815, n32816, n32826, n32827, n32831, n32835, n32836, n32839, n32840, n32843, n32844, n32845, n32847, n32855, n32856, n32857, n32861, n32864, n32865, n32870, n32889, n32891, n32894, n32895, n32897, n32898, n32902, n32903, n32904, n32910, n32913, n32914, n32915, n32919, n32921, n32922, n32925, n32927, n32928, n32929, n32932, n32933, n32934, n32938, n32941, n32945, n32951, n32954, n32955, n32959, n32961, n32962, n32963, n32964, n32967, n32974, n32975, n32976, n32981, n32984, n32989, n32992, n32996, n32997, n33003, n33004, n33008, n33011, n33014, n33015, n33017, n33019, n33023, n33030, n33033, n33039, n33041, n33042, n33043, n33048, n33050, n33051, n33052, n33053, n33059, n33060, n33062, n33065, n33066, n33067, n33069, n33070, n33071, n33074, n33076, n33080, n33081, n33086, n33089, n33090, n33094, n33095, n33097, n33100, n33102, n33103, n33104, n33106, n33118, n33121, n33123, n33128, n33130, n33134, n33135, n33137, n33139, n33140, n33147, n33148, n33153, n33154, n33155, n33161, n33166, n33169, n33172, n33176, n33184, n33187, n33199, n33200, n33201, n33204, n33205, n33207, n33210, n33212, n33213, n33214, n33218, n33219, n33222, n33225, n33228, n33230, n33235, n33237, n33239, n33243, n33246, n33251, n33252, n33255, n33258, n33260, n33261, n33268, n33270, n33271, n33272, n33273, n33275, n33276, n33278, n33280, n33281, n33283, n33286, n33290, n33296, n33298, n33303, n33308, n33312, n33314, n33322, n33323, n33326, n33328, n33333, n33334, n33350, n33357, n33370, n33371, n33375, n33376, n33381, n33382, n33383, n33389, n33390, n33391, n33393, n33394, n33395, n33397, n33399, n33402, n33403, n33409, n33412, n33417, n33420, n33421, n33425, n33426, n33428, n33429, n33430, n33435, n33438, n33439, n33440, n33444, n33445, n33449, n33454, n33456, n33459, n33460, n33461, n33465, n33470, n33471, n33472, n33473, n33475, n33478, n33480, n33482, n33483, n33484, n33488, n33494, n33495, n33498, n33499, n33505, n33507, n33512, n33520, n33523, n33525, n33533, n33535, n33541, n33542, n33544, n33545, n33549, n33558, n33566, n33567, n33569, n33571, n33572, n33575, n33580, n33581, n33582, n33585, n33589, n33591, n33592, n33595, n33596, n33597, n33598, n33600, n33601, n33602, n33603, n33604, n33605, n33607, n33608, n33612, n33615, n33617, n33624, n33632, n33633, n33634, n33636, n33638, n33644, n33645, n33648, n33649, n33662, n33664, n33665, n33666, n33667, n33668, n33669, n33671, n33676, n33682, n33686, n33688, n33690, n33696, n33698, n33699, n33702, n33704, n33715, n33716, n33717, n33719, n33728, n33732, n33736, n33737, n33739, n33744, n33748, n33756, n33760, n33762, n33768, n33770, n33771, n33781, n33790, n33791, n33806, n33808, n33810, n33816, n33817, n33819, n33823, n33831, n33834, n33838, n33840, n33843, n33845, n33847, n33855, n33857, n33860, n33865, n33868, n33874, n33883, n33885, n33886, n33887, n33893, n33894, n33895, n33902, n33910, n33912, n33913, n33918, n33920, n33923, n33924, n33926, n33931, n33932, n33938, n33939, n33941, n33942, n33954, n33957, n33958, n33959, n33962, n33964, n33981, n33982, n33988, n33989, n33991, n33999, n34007, n34012, n34013, n34014, n34015, n34017, n34018, n34022, n34027, n34029, n34030, n34034, n34038, n34041, n34048, n34051, n34056, n34064, n34069, n34071, n34075, n34078, n34079, n34080, n34083, n34086, n34087, n34089, n34091, n34094, n34099, n34101, n34104, n34111, n34113, n34126, n34134, n34138, n34139, n34140, n34144, n34152, n34154, n34157, n34159, n34162, n34164, n34167, n34168, n34169, n34172, n34173, n34175, n34176, n34182, n34190, n34191, n34192, n34194, n34200, n34203, n34204, n34207, n34208, n34211, n34213, n34215, n34216, n34219, n34220, n34222, n34224, n34226, n34227, n34230, n34234, n34238, n34241, n34249, n34254, n34255, n34256, n34258, n34262, n34264, n34268, n34269, n34272, n34273, n34275, n34280, n34283, n34286, n34288, n34291, n34297, n34304, n34308, n34311, n34315, n34317, n34320, n34326, n34327, n34328, n34329, n34332, n34333, n34335, n34339, n34340, n34342, n34348, n34349, n34353, n34354, n34357, n34360, n34362, n34366, n34367, n34368, n34370, n34377, n34381, n34382, n34383, n34385, n34387, n34391, n34394, n34395, n34398, n34402, n34404, n34407, n34408, n34415, n34423, n34428, n34429, n34431, n34434, n34438, n34441, n34443, n34444, n34452, n34453, n34464, n34465, n34472, n34474, n34475, n34476, n34477, n34479, n34482, n34483, n34485, n34486, n34489, n34491, n34492, n34504, n34506, n34507, n34509, n34510, n34511, n34513, n34515, n34516, n34518, n34520, n34524, n34529, n34530, n34538, n34543, n34550, n34551, n34553, n34559, n34562, n34573, n34575, n34582, n34584, n34588, n34592, n34601, n34603, n34607, n34609, n34610, n34611, n34615, n34617, n34620, n34621, n34632, n34634, n34635, n34639, n34645, n34651, n34652, n34654, n34656, n34658, n34661, n34664, n34666, n34668, n34669, n34676, n34684, n34690, n34691, n34692, n34694, n34695, n34696, n34700, n34702, n34706, n34709, n34710, n34714, n34715, n34716, n34717, n34718, n34721, n34723, n34733, n34734, n34736, n34737, n34739, n34740, n34747, n34755, n34757, n34759, n34760, n34761, n34762, n34765, n34768, n34770, n34776, n34779, n34782, n34783, n34784, n34785, n34786, n34790, n34791, n34792, n34793, n34798, n34801, n34802, n34803, n34805, n34812, n34813, n34816, n34817, n34819, n34820, n34824, n34825, n34828, n34834, n34835, n34838, n34843, n34846, n34849, n34852, n34858, n34859, n34860, n34862, n34864, n34866, n34872, n34873, n34875, n34876, n34880, n34884, n34887, n34888, n34890, n34892, n34894, n34902, n34905, n34916, n34924, n34927, n34930, n34931, n34935, n34936, n34941, n34942, n34943, n34947, n34949, n34950, n34952, n34955, n34964, n34966, n34969, n34971, n34972, n34973, n34974, n34975, n34976, n34980, n34981, n34989, n34991, n34997, n34998, n35003, n35004, n35008, n35010, n35011, n35012, n35014, n35016, n35023, n35031, n35037, n35038, n35040, n35041, n35044, n35047, n35051, n35061, n35068, n35072, n35075, n35076, n35079, n35080, n35081, n35084, n35090, n35094, n35102, n35105, n35106, n35112, n35114, n35116, n35121, n35122, n35124, n35127, n35130, n35137, n35138, n35141, n35142, n35157, n35158, n35162, n35164, n35165, n35170, n35182, n35183, n35184, n35194, n35195, n35201, n35202, n35205, n35213, n35214, n35216, n35219, n35223, n35226, n35229, n35231, n35233, n35235, n35238, n35243, n35245, n35250, n35251, n35255, n35270, n35271, n35272, n35273, n35274, n35276, n35277, n35285, n35287, n35292, n35293, n35294, n35297, n35303, n35306, n35307, n35312, n35316, n35317, n35320, n35325, n35329, n35335, n35336, n35339, n35341, n35347, n35348, n35360, n35361, n35364, n35365, n35367, n35369, n35372, n35382, n35390, n35393, n35397, n35404, n35405, n35410, n35412, n35420, n35421, n35426, n35430, n35432, n35434, n35437, n35447, n35450, n35451, n35452, n35454, n35455, n35461, n35462, n35465, n35466, n35473, n35475, n35478, n35480, n35483, n35484, n35487, n35489, n35491, n35493, n35494, n35505, n35506, n35509, n35510, n35515, n35518, n35520, n35523, n35528, n35535, n35537, n35539, n35540, n35541, n35543, n35546, n35552, n35556, n35559, n35562, n35566, n35568, n35572, n35580, n35581, n35590, n35597, n35599, n35602, n35607, n35610, n35614, n35616, n35617, n35622, n35628, n35634, n35636, n35638, n35639, n35640, n35641, n35644, n35646, n35648, n35651, n35654, n35656, n35657, n35658, n35660, n35662, n35664, n35667, n35671, n35673, n35679, n35683, n35685, n35686, n35688, n35689, n35693, n35696, n35699, n35706, n35708, n35709, n35712, n35713, n35714, n35717, n35719, n35727, n35729, n35730, n35733, n35736, n35738, n35741, n35742, n35744, n35746, n35748, n35750, n35753, n35761, n35763, n35765, n35772, n35773, n35774, n35775, n35778, n35780, n35783, n35784, n35787, n35788, n35789, n35790, n35792, n35794, n35809, n35810, n35812, n35813, n35817, n35819, n35824, n35825, n35826, n35827, n35829, n35830, n35834, n35839, n35850, n35854, n35857, n35859, n35866, n35867, n35871, n35873, n35874, n35877, n35879, n35881, n35882, n35883, n35886, n35887, n35888, n35890, n35902, n35904, n35909, n35912, n35915, n35916, n35920, n35922, n35925, n35928, n35930, n35937, n35939, n35942, n35945, n35946, n35951, n35956, n35960, n35963, n35964, n35967, n35968, n35969, n35970, n35976, n35978, n35985, n35990, n35991, n35993, n35997, n35999, n36007, n36009, n36010, n36012, n36014, n36015, n36018, n36021, n36023, n36028, n36032, n36033, n36034, n36039, n36040, n36045, n36046, n36049, n36054, n36056, n36062, n36064, n36067, n36071, n36075, n36078, n36079, n36082, n36084, n36085, n36088, n36090, n36095, n36096, n36099, n36101, n36104, n36110, n36119, n36120, n36126, n36128, n36129, n36132, n36136, n36137, n36142, n36144, n36147, n36149, n36152, n36156, n36157, n36162, n36165, n36166, n36167, n36168, n36171, n36173, n36179, n36183, n36184, n36185, n36190, n36199, n36200, n36203, n36204, n36207, n36208, n36211, n36213, n36217, n36218, n36220, n36221, n36223, n36237, n36240, n36243, n36244, n36245, n36248, n36253, n36254, n36255, n36258, n36268, n36269, n36270, n36280, n36283, n36287, n36290, n36291, n36292, n36297, n36299, n36302, n36303, n36305, n36306, n36310, n36311, n36312, n36314, n36316, n36320, n36321, n36323, n36324, n36327, n36332, n36334, n36335, n36340, n36343, n36349, n36350, n36352, n36357, n36359, n36360, n36361, n36369, n36370, n36375, n36377, n36379, n36382, n36384, n36386, n36389, n36392, n36397, n36399, n36402, n36405, n36407, n36409, n36411, n36414, n36417, n36418, n36438, n36440, n36441, n36444, n36445, n36446, n36447, n36449, n36450, n36454, n36459, n36460, n36461, n36462, n36476, n36479, n36485, n36486, n36487, n36494, n36495, n36496, n36504, n36508, n36509, n36510, n36511, n36513, n36514, n36517, n36520, n36523, n36530, n36533, n36535, n36538, n36541, n36544, n36547, n36550, n36551, n36555, n36559, n36568, n36572, n36573, n36574, n36579, n36581, n36582, n36586, n36589, n36590, n36591, n36593, n36606, n36612, n36614, n36616, n36620, n36628, n36631, n36632, n36637, n36641, n36643, n36648, n36652, n36658, n36659, n36660, n36670, n36676, n36681, n36685, n36690, n36692, n36693, n36694, n36696, n36698, n36700, n36704, n36708, n36710, n36712, n36714, n36726, n36728, n36731, n36732, n36736, n36739, n36741, n36745, n36750, n36751, n36753, n36757, n36759, n36761, n36762, n36763, n36766, n36772, n36775, n36776, n36781, n36790, n36792, n36794, n36796, n36800, n36801, n36802, n36814, n36815, n36819, n36826, n36827, n36830, n36832, n36833, n36836, n36837, n36838, n36841, n36843, n36844, n36847, n36849, n36856, n36857, n36860, n36868, n36875, n36876, n36877, n36878, n36883, n36884, n36885, n36894, n36895, n36899, n36901, n36903, n36904, n36905, n36913, n36914, n36919, n36924, n36927, n36935, n36940, n36941, n36942, n36943, n36944, n36945, n36947, n36953, n36957, n36963, n36965, n36966, n36968, n36969, n36971, n36973, n36974, n36975, n36976, n36979, n36983, n36984, n36986, n36987, n36988, n36989, n36993, n36994, n36996, n36997, n37005, n37007, n37008, n37009, n37010, n37012, n37015, n37022, n37027, n37030, n37033, n37034, n37036, n37040, n37041, n37045, n37047, n37049, n37050, n37051, n37056, n37057, n37058, n37060, n37062, n37064, n37069, n37072, n37073, n37074, n37076, n37077, n37078, n37080, n37081, n37082, n37086, n37095, n37096, n37098, n37101, n37102, n37104, n37105, n37106, n37107, n37110, n37112, n37114, n37116, n37118, n37119, n37122, n37126, n37127, n37129, n37130, n37132, n37133, n37134, n37135, n37136, n37138, n37143, n37146, n37147, n37151, n37160, n37168, n37172, n37174, n37175, n37178, n37183, n37184, n37188, n37189, n37190, n37191, n37203, n37207, n37208, n37209, n37210, n37217, n37219, n37221, n37223, n37224, n37225, n37227, n37229, n37233, n37236, n37240, n37241, n37246, n37250, n37255, n37257, n37258, n37259, n37261, n37262, n37263, n37268, n37270, n37281, n37283, n37287, n37291, n37292, n37293, n37295, n37296, n37298, n37301, n37303, n37314, n37315, n37317, n37318, n37323, n37329, n37330, n37332, n37333, n37337, n37340, n37344, n37356, n37357, n37361, n37362, n37364, n37367, n37369, n37370, n37372, n37384, n37385, n37395, n37396, n37397, n37398, n37400, n37406, n37412, n37413, n37416, n37422, n37423, n37429, n37431, n37436, n37441, n37447, n37449, n37451, n37452, n37456, n37458, n37459, n37461, n37462, n37465, n37468, n37471, n37472, n37473, n37474, n37476, n37478, n37484, n37487, n37489, n37491, n37493, n37494, n37495, n37499, n37507, n37510, n37511, n37516, n37522, n37525, n37530, n37539, n37541, n37544, n37555, n37560, n37561, n37562, n37567, n37568, n37569, n37570, n37577, n37587, n37589, n37594, n37597, n37599, n37606, n37615, n37619, n37626, n37627, n37634, n37637, n37640, n37641, n37642, n37652, n37653, n37657, n37662, n37665, n37667, n37669, n37675, n37676, n37679, n37681, n37682, n37683, n37685, n37686, n37689, n37694, n37698, n37699, n37700, n37702, n37703, n37704, n37706, n37718, n37719, n37721, n37722, n37725, n37732, n37733, n37735, n37741, n37744, n37755, n37758, n37760, n37762, n37765, n37767, n37771, n37784, n37785, n37787, n37794, n37799, n37800, n37801, n37802, n37805, n37810, n37812, n37815, n37817, n37818, n37821, n37822, n37823, n37824, n37825, n37829, n37834, n37835, n37836, n37839, n37842, n37843, n37845, n37848, n37849, n37850, n37856, n37870, n37873, n37880, n37881, n37883, n37886, n37897, n37899, n37901, n37902, n37906, n37910, n37916, n37925, n37926, n37931, n37936, n37942, n37947, n37951, n37954, n37955, n37956, n37958, n37962, n37963, n37974, n37975, n37976, n37978, n37984, n37985, n37991, n37992, n37993, n37995, n37996, n37997, n38001, n38002, n38004, n38007, n38008, n38013, n38014, n38018, n38020, n38021, n38028, n38036, n38037, n38038, n38039, n38042, n38044, n38058, n38060, n38061, n38068, n38070, n38072, n38073, n38076, n38079, n38081, n38085, n38086, n38087, n38089, n38101, n38102, n38106, n38107, n38110, n38112, n38115, n38120, n38123, n38130, n38131, n38138, n38140, n38156, n38158, n38162, n38165, n38167, n38169, n38170, n38172, n38173, n38174, n38176, n38180, n38181, n38184, n38185, n38195, n38198, n38200, n38201, n38203, n38208, n38211, n38214, n38215, n38216, n38219, n38223, n38229, n38231, n38236, n38239, n38241, n38242, n38244, n38251, n38252, n38253, n38254, n38256, n38257, n38258, n38265, n38266, n38269, n38272, n38273, n38274, n38280, n38282, n38286, n38291, n38292, n38295, n38298, n38300, n38301, n38303, n38306, n38310, n38311, n38317, n38320, n38323, n38327, n38330, n38333, n38334, n38343, n38344, n38347, n38348, n38352, n38355, n38356, n38357, n38358, n38361, n38363, n38364, n38366, n38367, n38370, n38373, n38377, n38382, n38383, n38390, n38395, n38401, n38406, n38414, n38417, n38420, n38425, n38432, n38441, n38442, n38450, n38451, n38456, n38457, n38463, n38466, n38475, n38477, n38481, n38484, n38485, n38490, n38491, n38492, n38499, n38500, n38502, n38503, n38513, n38514, n38516, n38519, n38523, n38526, n38529, n38532, n38534, n38537, n38543, n38554, n38560, n38564, n38565, n38566, n38568, n38578, n38581, n38584, n38590, n38592, n38593, n38594, n38595, n38600, n38601, n38603, n38605, n38606, n38607, n38610, n38611, n38612, n38613, n38617, n38621, n38624, n38625, n38626, n38635, n38640, n38641, n38642, n38644, n38645, n38647, n38649, n38651, n38661, n38666, n38673, n38677, n38678, n38681, n38683, n38685, n38690, n38691, n38692, n38693, n38694, n38698, n38701, n38702, n38703, n38706, n38709, n38711, n38716, n38724, n38727, n38729, n38732, n38735, n38738, n38742, n38743, n38745, n38748, n38752, n38754, n38760, n38763, n38773, n38774, n38777, n38783, n38787, n38789, n38790, n38797, n38799, n38800, n38804, n38807, n38809, n38810, n38811, n38814, n38816, n38818, n38820, n38822, n38824, n38825, n38828, n38831, n38833, n38837, n38839, n38843, n38846, n38847, n38848, n38852, n38854, n38855, n38860, n38861, n38863, n38864, n38866, n38871, n38872, n38873, n38875, n38878, n38879, n38881, n38894, n38896, n38899, n38900, n38902, n38908, n38909, n38912, n38927, n38929, n38930, n38935, n38936, n38942, n38943, n38945, n38948, n38955, n38958, n38959, n38963, n38965, n38969, n38973, n38975, n38978, n38979, n38981, n38982, n38983, n38985, n38988, n38989, n38991, n38992, n38995, n38996, n38997, n38998, n39004, n39006, n39009, n39012, n39013, n39015, n39018, n39022, n39027, n39032, n39039, n39040, n39052, n39056, n39058, n39067, n39072, n39075, n39080, n39083, n39085, n39087, n39088, n39094, n39095, n39096, n39099, n39100, n39113, n39114, n39115, n39116, n39118, n39120, n39121, n39127, n39130, n39138, n39140, n39141, n39145, n39146, n39147, n39150, n39152, n39158, n39159, n39162, n39167, n39174, n39179, n39180, n39183, n39189, n39191, n39192, n39193, n39198, n39199, n39202, n39205, n39207, n39210, n39212, n39215, n39221, n39226, n39231, n39232, n39235, n39237, n39239, n39240, n39245, n39246, n39254, n39256, n39259, n39263, n39264, n39265, n39266, n39269, n39275, n39276, n39279, n39280, n39282, n39288, n39292, n39296, n39300, n39302, n39307, n39309, n39312, n39313, n39314, n39315, n39317, n39319, n39323, n39326, n39333, n39341, n39343, n39344, n39346, n39349, n39350, n39355, n39356, n39362, n39363, n39364, n39365, n39367, n39370, n39371, n39374, n39377, n39381, n39382, n39385, n39386, n39387, n39392, n39397, n39399, n39400, n39402, n39405, n39408, n39412, n39415, n39416, n39424, n39426, n39427, n39428, n39430, n39434, n39435, n39446, n39447, n39448, n39449, n39454, n39455, n39457, n39458, n39460, n39462, n39464, n39466, n39469, n39470, n39471, n39474, n39476, n39478, n39479, n39481, n39483, n39492, n39493, n39495, n39498, n39504, n39505, n39510, n39513, n39514, n39515, n39518, n39520, n39523, n39525, n39529, n39532, n39538, n39541, n39542, n39546, n39549, n39550, n39559, n39562, n39577, n39580, n39583, n39585, n39590, n39594, n39597, n39599, n39600, n39601, n39604, n39605, n39607, n39612, n39614, n39619, n39620, n39630, n39632, n39639, n39640, n39641, n39644, n39648, n39650, n39651, n39652, n39655, n39657, n39659, n39660, n39665, n39667, n39668, n39670, n39671, n39673, n39675, n39676, n39677, n39678, n39683, n39684, n39688, n39689, n39690, n39691, n39693, n39694, n39696, n39705, n39710, n39712, n39716, n39719, n39723, n39728, n39732, n39735, n39738, n39739, n39742, n39744, n39746, n39747, n39749, n39750, n39752, n39753, n39762, n39764, n39767, n39769, n39772, n39774, n39775, n39777, n39780, n39784, n39785, n39796, n39799, n39802, n39807, n39812, n39819, n39824, n39826, n39829, n39832, n39835, n39836, n39840, n39844, n39845, n39857, n39858, n39859, n39861, n39869, n39873, n39874, n39878, n39881, n39887, n39888, n39891, n39893, n39898, n39900, n39903, n39908, n39909, n39911, n39916, n39919, n39932, n39934, n39937, n39938, n39941, n39943, n39945, n39947, n39949, n39953, n39958, n39964, n39967, n39970, n39971, n39979, n39981, n39983, n39986, n39989, n39997, n39998, n40000, n40002, n40004, n40010, n40012, n40015, n40018, n40020, n40021, n40022, n40025, n40026, n40029, n40030, n40033, n40034, n40035, n40040, n40041, n40042, n40043, n40045, n40049, n40050, n40059, n40060, n40065, n40067, n40072, n40075, n40079, n40086, n40087, n40093, n40095, n40097, n40098, n40100, n40105, n40110, n40113, n40117, n40122, n40123, n40130, n40131, n40132, n40135, n40140, n40141, n40146, n40149, n40150, n40151, n40162, n40163, n40165, n40167, n40175, n40182, n40183, n40184, n40185, n40186, n40187, n40189, n40190, n40193, n40194, n40195, n40197, n40198, n40203, n40215, n40219, n40224, n40226, n40228, n40235, n40241, n40243, n40246, n40251, n40255, n40256, n40257, n40262, n40264, n40265, n40266, n40269, n40271, n40273, n40277, n40283, n40285, n40286, n40290, n40292, n40293, n40295, n40297, n40298, n40304, n40305, n40310, n40312, n40317, n40323, n40327, n40328, n40337, n40340, n40343, n40356, n40359, n40366, n40368, n40374, n40378, n40380, n40383, n40387, n40388, n40391, n40395, n40401, n40402, n40403, n40407, n40411, n40414, n40419, n40426, n40429, n40430, n40431, n40432, n40440, n40442, n40448, n40449, n40451, n40453, n40460, n40463, n40471, n40473, n40475, n40476, n40480, n40482, n40485, n40487, n40496, n40501, n40503, n40504, n40508, n40512, n40515, n40519, n40520, n40521, n40524, n40529, n40532, n40534, n40536, n40538, n40539, n40540, n40541, n40543, n40548, n40555, n40556, n40559, n40569, n40570, n40572, n40576, n40580, n40581, n40582, n40584, n40586, n40588, n40593, n40597, n40600, n40603, n40606, n40609, n40611, n40622, n40623, n40624, n40625, n40628, n40629, n40635, n40638, n40639, n40641, n40643, n40644, n40646, n40651, n40652, n40653, n40656, n40660, n40663, n40666, n40667, n40669, n40672, n40674, n40679, n40689, n40690, n40692, n40703, n40704, n40705, n40706, n40707, n40717, n40718, n40725, n40726, n40727, n40730, n40734, n40737, n40741, n40743, n40745, n40751, n40752, n40753, n40754, n40755, n40759, n40764, n40765, n40774, n40777, n40781, n40782, n40783, n40784, n40785, n40792, n40796, n40799, n40800, n40802, n40803, n40806, n40807, n40808, n40812, n40814, n40815, n40817, n40818, n40819, n40820, n40821, n40824, n40825, n40835, n40842, n40847, n40848, n40851, n40853, n40864, n40867, n40873, n40874, n40877, n40881, n40882, n40883, n40884, n40885, n40887, n40889, n40890, n40891, n40894, n40895, n40897, n40898, n40900, n40901, n40912, n40914, n40916, n40918, n40921, n40925, n40927, n40928, n40932, n40938, n40941, n40943, n40948, n40951, n40952, n40953, n40958, n40964, n40966, n40967, n40968, n40970, n40972, n40975, n40976, n40977, n40980, n40982, n40985, n40988, n40992, n40996, n41001, n41002, n41004, n41005, n41007, n41009, n41011, n41014, n41015, n41016, n41019, n41025, n41030, n41040, n41042, n41044, n41051, n41056, n41058, n41061, n41077, n41082, n41086, n41087, n41089, n41090, n41091, n41092, n41099, n41102, n41109, n41112, n41113, n41116, n41118, n41125, n41126, n41133, n41137, n41140, n41141, n41142, n41143, n41155, n41156, n41157, n41158, n41163, n41164, n41169, n41175, n41177, n41180, n41188, n41191, n41192, n41197, n41198, n41203, n41205, n41206, n41207, n41217, n41218, n41221, n41222, n41230, n41231, n41233, n41238, n41241, n41243, n41245, n41251, n41254, n41258, n41261, n41264, n41268, n41269, n41270, n41272, n41274, n41275, n41277, n41281, n41288, n41291, n41292, n41298, n41301, n41307, n41308, n41314, n41317, n41320, n41326, n41327, n41328, n41332, n41335, n41338, n41340, n41345, n41346, n41347, n41351, n41358, n41361, n41365, n41366, n41370, n41383, n41385, n41396, n41398, n41402, n41408, n41411, n41413, n41416, n41420, n41422, n41423, n41427, n41429, n41436, n41442, n41444, n41447, n41448, n41449, n41451, n41454, n41455, n41463, n41465, n41468, n41469, n41472, n41475, n41477, n41478, n41480, n41482, n41485, n41487, n41488, n41492, n41498, n41501, n41502, n41503, n41507, n41508, n41509, n41510, n41516, n41517, n41523, n41524, n41533, n41534, n41535, n41538, n41539, n41546, n41548, n41557, n41563, n41581, n41585, n41592, n41594, n41599, n41602, n41605, n41610, n41611, n41614, n41615, n41617, n41618, n41620, n41624, n41625, n41626, n41627, n41629, n41630, n41631, n41634, n41635, n41637, n41641, n41644, n41647, n41648, n41653, n41656, n41663, n41672, n41676, n41677, n41678, n41682, n41683, n41684, n41686, n41688, n41689, n41690, n41691, n41693, n41694, n41696, n41702, n41703, n41704, n41705, n41706, n41711, n41713, n41718, n41719, n41721, n41722, n41723, n41729, n41730, n41734, n41735, n41738, n41739, n41740, n41742, n41744, n41746, n41747, n41748, n41755, n41756, n41757, n41762, n41771, n41772, n41773, n41774, n41779, n41780, n41782, n41784, n41785, n41789, n41790, n41791, n41794, n41799, n41801, n41808, n41809, n41816, n41817, n41819, n41821, n41824, n41825, n41826, n41828, n41834, n41841, n41847, n41850, n41852, n41853, n41854, n41855, n41857, n41858, n41863, n41864, n41868, n41870, n41872, n41879, n41884, n41886, n41905, n41909, n41913, n41914, n41922, n41925, n41926, n41928, n41930, n41934, n41939, n41940, n41946, n41949, n41954, n41955, n41961, n41963, n41967, n41971, n41974, n41976, n41978, n41981, n41987, n41989, n41997, n41999, n42007, n42009, n42010, n42017, n42021, n42023, n42027, n42032, n42034, n42036, n42037, n42038, n42042, n42043, n42044, n42046, n42048, n42049, n42050, n42052, n42053, n42057, n42058, n42060, n42063, n42065, n42067, n42073, n42075, n42077, n42079, n42081, n42083, n42090, n42093, n42098, n42099, n42102, n42111, n42112, n42117, n42119, n42120, n42121, n42122, n42123, n42124, n42126, n42130, n42134, n42135, n42137, n42139, n42143, n42147, n42148, n42155, n42157, n42159, n42161, n42163, n42165, n42166, n42167, n42171, n42172, n42173, n42179, n42183, n42184, n42190, n42193, n42196, n42202, n42205, n42215, n42216, n42223, n42226, n42228, n42231, n42236, n42239, n42244, n42251, n42253, n42261, n42266, n42268, n42274, n42275, n42277, n42278, n42282, n42285, n42289, n42291, n42293, n42298, n42307, n42309, n42312, n42314, n42316, n42319, n42321, n42324, n42325, n42329, n42333, n42334, n42335, n42338, n42339, n42340, n42341, n42346, n42347, n42348, n42349, n42358, n42359, n42361, n42366, n42371, n42372, n42373, n42374, n42375, n42377, n42379, n42380, n42383, n42387, n42391, n42394, n42396, n42401, n42402, n42403, n42405, n42408, n42409, n42416, n42419, n42424, n42425, n42429, n42435, n42437, n42442, n42443, n42444, n42445, n42447, n42452, n42454, n42455, n42456, n42467, n42474, n42478, n42479, n42481, n42485, n42486, n42489, n42490, n42495, n42497, n42501, n42504, n42506, n42507, n42509, n42510, n42511, n42514, n42518, n42520, n42521, n42525, n42526, n42530, n42533, n42536, n42537, n42538, n42539, n42540, n42543, n42544, n42546, n42550, n42555, n42557, n42558, n42560, n42566, n42567, n42568, n42570, n42574, n42576, n42580, n42583, n42593, n42594, n42595, n42597, n42598, n42600, n42604, n42608, n42613, n42617, n42618, n42621, n42623, n42625, n42626, n42627, n42633, n42634, n42637, n42640, n42641, n42643, n42644, n42647, n42648, n42652, n42654, n42656, n42658, n42660, n42661, n42663, n42666, n42668, n42669, n42670, n42674, n42675, n42676, n42677, n42678, n42680, n42689, n42690, n42692, n42694, n42695, n42696, n42697, n42705, n42706, n42707, n42709, n42712, n42715, n42716, n42720, n42722, n42728, n42735, n42736, n42738, n42743, n42744, n42749, n42750, n42751, n42752, n42759, n42761, n42762, n42767, n42770, n42772, n42783, n42788, n42790, n42792, n42793, n42798, n42800, n42806, n42807, n42812, n42819, n42827, n42828, n42829, n42832, n42834, n42835, n42836, n42839, n42840, n42841, n42844, n42851, n42856, n42858, n42861, n42862, n42865, n42867, n42870, n42873, n42877, n42878, n42879, n42881, n42883, n42886, n42890, n42891, n42895, n42899, n42901, n42907, n42916, n42930, n42931, n42933, n42934, n42935, n42937, n42943, n42945, n42948, n42954, n42955, n42960, n42961, n42962, n42967, n42968, n42970, n42975, n42976, n42978, n42980, n42981, n42982, n42992, n42998, n43000, n43007, n43015, n43017, n43023, n43025, n43032, n43045, n43046, n43053, n43055, n43056, n43067, n43073, n43074, n43076, n43077, n43078, n43085, n43086, n43087, n43090, n43092, n43096, n43097, n43099, n43100, n43101, n43102, n43103, n43104, n43109, n43120, n43128, n43129, n43133, n43136, n43138, n43149, n43155, n43160, n43167, n43171, n43172, n43176, n43177, n43178, n43182, n43184, n43185, n43186, n43195, n43198, n43199, n43201, n43202, n43205, n43208, n43209, n43213, n43217, n43218, n43220, n43221, n43224, n43227, n43228, n43229, n43231, n43235, n43239, n43249, n43251, n43254, n43257, n43261, n43264, n43265, n43268, n43269, n43271, n43272, n43273, n43276, n43278, n43282, n43286, n43291, n43292, n43293, n43296, n43303, n43304, n43309, n43311, n43312, n43314, n43315, n43324, n43325, n43326, n43327, n43329, n43330, n43331, n43333, n43344, n43346, n43347, n43358, n43359, n43360, n43363, n43366, n43367, n43370, n43371, n43375, n43385, n43389, n43395, n43396, n43398, n43405, n43406, n43408, n43410, n43415, n43419, n43427, n43429, n43435, n43436, n43441, n43445, n43451, n43453, n43454, n43464, n43471, n43475, n43523, n43534, n43539, n43543, n43554, n43557, n43559, n43561, n43564, n43575, n43582, n43585, n43593, n43620, n43627, n43631, n43633, n43643, n43675, n43690, n43703, n43729, n43747, n43760, n43762, n43764, n43770, n43771, n43776, n43796, n43803, n43844, n43858, n43878, n43890, n43899, n43920, n43933, n43940, n43941, n43954, n43963, n43993, n43998, n44006, n44054, n44068, n44096, n44104, n44120, n44134, n44138, n44140, n44157, n44170, n44173, n44176, n44179, n44180, n44211, n44214, n44223, n44228, n44231, n44245, n44247, n44253, n44260, n44270, n44280, n44287, n44315, n44336, n44337, n44340, n44344, n44351, n44358, n44361, n44362, n44374, n44382, n44383, n44398, n44439, n44449, n44454, n44455, n44460, n44468, n44477, n44485, n44487, n44490, n44501, n44524, n44535, n44542, n44546, n44565, n44571, n44584, n44591, n44603, n44623, n44624, n44640, n44642, n44663, n44665, n44697, n44703, n44708, n44710, n44720, n44721, n44727, n44731, n44747, n44765, n44766, n44767, n44790, n44794, n44796, n44800, n44822, n44834, n44849, n44887, n44892, n44895, n44937, n44944, n44951, n44967, n44970, n44975, n44987, n44988, n45019, n45035, n45049, n45062, n45077, n45083, n45104, n45112, n45126, n45134, n45137, n45140, n45141, n45152, n45156, n45177, n45184, n45204, n45207, n45211, n45218, n45226, n45239, n45240, n45241, n45264, n45265, n45266, n45268, n45302, n45306, n45315, n45334, n45350, n45351, n45368, n45371, n45392, n45400, n45401, n45404, n45428, n45432, n45437, n45446, n45453, n45454, n45455, n45456, n45457, n45463, n45470, n45482, n45510, n45512, n45528, n45529, n45534, n45546, n45560, n45565, n45582, n45583, n45591, n45594, n45596, n45598, n45604, n45624, n45626, n45632, n45644, n45645, n45651, n45668, n45670, n45672, n45675, n45684, n45700, n45704, n45715, n45731, n45734, n45738, n45755, n45767, n45777, n45781, n45785, n45788, n45794, n45832, n45864, n45900, n45937, n45943, n45959, n45970, n45977, n45978, n45982, n45998, n46001, n46009, n46010, n46033, n46046, n46050, n46055, n46062, n46076, n46083, n46084, n46088, n46119, n46120, n46130, n46138, n46165, n46189, n46199, n46224, n46225, n46240, n46250, n46259, n46266, n46279, n46287, n46294, n46300, n46301, n46308, n46313, n46334, n46335, n46363, n46364, n46383, n46386, n46390, n46392, n46418, n46427, n46458, n46482, n46488, n46502, n46504, n46516, n46522, n46535, n46595, n46600, n46607, n46630, n46652, n46663, n46670, n46698, n46706, n46711, n46724, n46739, n46755, n46770, n46771, n46789, n46811, n46831, n46842, n46849, n46858, n46861, n46901, n46927, n46930, n46938, n46943, n46944, n46974, n46986, n46996, n47000, n47022, n47033, n47057, n47085, n47114, n47117, n47126, n47132, n47140, n47144, n47154, n47169, n47183, n47194, n47195, n47218, n47233, n47245, n47265, n47333, n47334, n47375, n47377, n47419, n47431, n47451, n47454, n47471, n47475, n47495, n47499, n47509, n47514, n47516, n47535, n47546, n47611, n47621, n47629, n47635, n47637, n47638, n47640, n47645, n47661, n47663, n47669, n47673, n47715, n47717, n47727, n47740, n47752, n47758, n47771, n47809, n47838, n47844, n47873, n47879, n47902, n47921, n47924, n47947, n47956, n48028, n48039, n48048, n48057, n48060, n48086, n48101, n48112, n48114, n48128, n48134, n48136, n48144, n48146, n48151, n48163, n48166, n48186, n48209, n48215, n48218, n48232, n48239, n48247, n48261, n48266, n48276, n48285, n48301, n48304, n48305, n48310, n48322, n48324, n48330, n48348, n48355, n48361, n48373, n48376, n48378, n48381, n48402, n48403, n48434, n48453, n48458, n48460, n48467, n48487, n48509, n48510, n48514, n48520, n48522, n48544, n48548, n48554, n48556, n48577, n48580, n48599, n48608, n48640, n48648, n48678, n48703, n48717, n48719, n48733, n48743, n48761, n48816, n48827, n48831, n48834, n48891, n48893, n48896, n48908, n48931, n48942, n48953, n48968, n48970, n48976, n48987, n48993, n49010, n49027, n49029, n49031, n49032, n49047, n49067, n49089, n49096, n49106, n49116, n49117, n49122, n49129, n49134, n49152, n49179, n49184, n49194, n49203, n49219, n49221, n49238, n49264, n49273, n49278, n49283, n49299, n49307, n49316, n49329, n49332, n49337, n49361, n49362, n49365, n49376, n49379, n49421, n49427, n49440, n49455, n49458, n49466, n49472, n49482, n49505, n49553, n49554, n49561, n49588, n49615, n49621, n49623, n49627, n49642, n49654, n49659, n49671, n49686, n49704, n49738, n49762, n49764, n49766, n49775, n49786, n49793, n49833, n49834, n49859, n49893, n49897, n49900, n49902, n49916, n49922, n49968, n49971, n49978, n49984, n49990, n50002, n50029, n50052, n50083, n50088, n50097, n50107, n50112, n50114, n50118, n50127, n50128, n50141, n50155, n50156, n50176, n50178, n50184, n50198, n50199, n50202, n50207, n50219, n50228, n50233, n50245, n50257, n50261, n50269, n50271, n50275, n50311, n50314, n50322, n50348, n50365, n50394, n50395, n50423, n50431, n50455, n50460, n50505, n50511, n50534, n50568, n50587, n50591, n50594, n50595, n50597, n50602, n50626, n50634, n50647, n50666, n50686, n50692, n50704, n50727, n50740, n50823, n50854, n50861, n50863, n50877, n50889, n50890, n50897, n50907, n50909, n50917, n50931, n50935, n50938, n50940, n50943, n50947, n50948, n50951, n50967, n50974, n50977, n50987, n51024, n51025, n51035, n51038, n51042, n51046, n51051, n51063, n51088, n51092, n51099, n51100, n51104, n51109, n51138, n51149, n51158, n51192, n51196, n51199, n51218, n51227, n51241, n51243, n51247, n51264, n51275, n51293, n51307, n51323, n51330, n51337, n51339, n51354, n51356, n51370, n51373, n51380, n51391, n51393, n51404, n51429, n51451, n51462, n51472, n51498, n51501, n51503, n51516, n51521, n51532, n51535, n51536, n51540, n51549, n51571, n51585, n51611, n51734, n51744, n51753, n51843, n51866, n51895, n51925, n51936, n51972, n52010, n52024, n52068, n52084, n52088, n52093, n52104, n52181, n52206, n52238, n52326, n52328, n52430, n52454, n52518, n52545, n52577, n52605, n52607, n52612, n52635, n52660, n52799, n52813, n52837, n52881, n52939, n52966, n53023, n53027, n53065, n53076, n53203, n53232, n53324, n53352, n53362, n53365, n53392, n53453, n53600, n53631, n53799, n53862, n53995, n54070;

    NANDX1 U1 (.A1(N1), .A2(N2), .ZN(n12873));
    NANDX1 U2 (.A1(N3), .A2(N4), .ZN(N12874));
    NANDX1 U3 (.A1(N5), .A2(N6), .ZN(n12875));
    NANDX1 U4 (.A1(N7), .A2(N8), .ZN(n12876));
    NOR2X1 U5 (.A1(N9), .A2(N10), .ZN(N12877));
    NOR2X1 U6 (.A1(N11), .A2(N12), .ZN(n12878));
    NANDX1 U7 (.A1(N13), .A2(N14), .ZN(n12879));
    NANDX1 U8 (.A1(N15), .A2(N16), .ZN(n12880));
    NOR2X1 U9 (.A1(N17), .A2(N18), .ZN(N12881));
    NANDX1 U10 (.A1(N19), .A2(N20), .ZN(n12882));
    NOR2X1 U11 (.A1(N21), .A2(N22), .ZN(n12883));
    NANDX1 U12 (.A1(N23), .A2(N24), .ZN(n12884));
    NANDX1 U13 (.A1(N25), .A2(N26), .ZN(n12885));
    NOR2X1 U14 (.A1(N27), .A2(N28), .ZN(n12886));
    NOR2X1 U15 (.A1(N29), .A2(N30), .ZN(n12887));
    NOR2X1 U16 (.A1(N31), .A2(N32), .ZN(n12888));
    NOR2X1 U17 (.A1(N33), .A2(N34), .ZN(n12889));
    NOR2X1 U18 (.A1(N35), .A2(N36), .ZN(n12890));
    NANDX1 U19 (.A1(N37), .A2(N38), .ZN(N12891));
    NOR2X1 U20 (.A1(N39), .A2(N40), .ZN(N12892));
    NANDX1 U21 (.A1(N41), .A2(N42), .ZN(n12893));
    NANDX1 U22 (.A1(N43), .A2(N44), .ZN(n12894));
    NOR2X1 U23 (.A1(N45), .A2(N46), .ZN(n12895));
    NOR2X1 U24 (.A1(N47), .A2(N48), .ZN(n12896));
    NOR2X1 U25 (.A1(N49), .A2(N50), .ZN(N12897));
    NANDX1 U26 (.A1(N51), .A2(N52), .ZN(n12898));
    NANDX1 U27 (.A1(N53), .A2(N54), .ZN(N12899));
    NANDX1 U28 (.A1(N55), .A2(N56), .ZN(n12900));
    NANDX1 U29 (.A1(N57), .A2(N58), .ZN(n12901));
    NOR2X1 U30 (.A1(N59), .A2(N60), .ZN(n12902));
    NOR2X1 U31 (.A1(N61), .A2(N62), .ZN(n12903));
    NOR2X1 U32 (.A1(N63), .A2(N64), .ZN(n12904));
    NANDX1 U33 (.A1(N65), .A2(N66), .ZN(N12905));
    NANDX1 U34 (.A1(N67), .A2(N68), .ZN(n12906));
    NANDX1 U35 (.A1(N69), .A2(N70), .ZN(n12907));
    NOR2X1 U36 (.A1(N71), .A2(N72), .ZN(N12908));
    NANDX1 U37 (.A1(N73), .A2(N74), .ZN(n12909));
    NOR2X1 U38 (.A1(N75), .A2(N76), .ZN(n12910));
    NANDX1 U39 (.A1(N77), .A2(N78), .ZN(N12911));
    NANDX1 U40 (.A1(N79), .A2(N80), .ZN(n12912));
    NANDX1 U41 (.A1(N81), .A2(N82), .ZN(n12913));
    NANDX1 U42 (.A1(N83), .A2(N84), .ZN(n12914));
    NOR2X1 U43 (.A1(N85), .A2(N86), .ZN(n12915));
    NANDX1 U44 (.A1(N87), .A2(N88), .ZN(N12916));
    NOR2X1 U45 (.A1(N89), .A2(N90), .ZN(n12917));
    NOR2X1 U46 (.A1(N91), .A2(N92), .ZN(N12918));
    NANDX1 U47 (.A1(N93), .A2(N94), .ZN(n12919));
    NOR2X1 U48 (.A1(N95), .A2(N96), .ZN(N12920));
    NANDX1 U49 (.A1(N97), .A2(N98), .ZN(n12921));
    NOR2X1 U50 (.A1(N99), .A2(N100), .ZN(n12922));
    NANDX1 U51 (.A1(N101), .A2(N102), .ZN(n12923));
    NOR2X1 U52 (.A1(N103), .A2(N104), .ZN(N12924));
    NOR2X1 U53 (.A1(N105), .A2(N106), .ZN(N12925));
    NANDX1 U54 (.A1(N107), .A2(N108), .ZN(n12926));
    NOR2X1 U55 (.A1(N109), .A2(N110), .ZN(n12927));
    NOR2X1 U56 (.A1(N111), .A2(N112), .ZN(n12928));
    NOR2X1 U57 (.A1(N113), .A2(N114), .ZN(n12929));
    NANDX1 U58 (.A1(N115), .A2(N116), .ZN(n12930));
    NANDX1 U59 (.A1(N117), .A2(N118), .ZN(N12931));
    NANDX1 U60 (.A1(N119), .A2(N120), .ZN(n12932));
    NOR2X1 U61 (.A1(N121), .A2(N122), .ZN(N12933));
    NANDX1 U62 (.A1(N123), .A2(N124), .ZN(n12934));
    NOR2X1 U63 (.A1(N125), .A2(N126), .ZN(n12935));
    NANDX1 U64 (.A1(N127), .A2(N128), .ZN(n12936));
    NOR2X1 U65 (.A1(N129), .A2(N130), .ZN(n12937));
    NANDX1 U66 (.A1(N131), .A2(N132), .ZN(n12938));
    NANDX1 U67 (.A1(N133), .A2(N134), .ZN(n12939));
    NANDX1 U68 (.A1(N135), .A2(N136), .ZN(n12940));
    NOR2X1 U69 (.A1(N137), .A2(N138), .ZN(n12941));
    NANDX1 U70 (.A1(N139), .A2(N140), .ZN(n12942));
    NOR2X1 U71 (.A1(N141), .A2(N142), .ZN(N12943));
    NANDX1 U72 (.A1(N143), .A2(N144), .ZN(n12944));
    NOR2X1 U73 (.A1(N145), .A2(N146), .ZN(n12945));
    NANDX1 U74 (.A1(N147), .A2(N148), .ZN(n12946));
    NOR2X1 U75 (.A1(N149), .A2(N150), .ZN(n12947));
    NOR2X1 U76 (.A1(N151), .A2(N152), .ZN(n12948));
    NANDX1 U77 (.A1(N153), .A2(N154), .ZN(N12949));
    NOR2X1 U78 (.A1(N155), .A2(N156), .ZN(n12950));
    NANDX1 U79 (.A1(N157), .A2(N158), .ZN(n12951));
    NOR2X1 U80 (.A1(N159), .A2(N160), .ZN(N12952));
    NOR2X1 U81 (.A1(N161), .A2(N162), .ZN(n12953));
    NOR2X1 U82 (.A1(N163), .A2(N164), .ZN(n12954));
    NOR2X1 U83 (.A1(N165), .A2(N166), .ZN(n12955));
    NOR2X1 U84 (.A1(N167), .A2(N168), .ZN(n12956));
    NANDX1 U85 (.A1(N169), .A2(N170), .ZN(n12957));
    NANDX1 U86 (.A1(N171), .A2(N172), .ZN(N12958));
    NOR2X1 U87 (.A1(N173), .A2(N174), .ZN(n12959));
    NANDX1 U88 (.A1(N175), .A2(N176), .ZN(n12960));
    NOR2X1 U89 (.A1(N177), .A2(N178), .ZN(n12961));
    NOR2X1 U90 (.A1(N179), .A2(N180), .ZN(n12962));
    NOR2X1 U91 (.A1(N181), .A2(N182), .ZN(n12963));
    NOR2X1 U92 (.A1(N183), .A2(N184), .ZN(n12964));
    NANDX1 U93 (.A1(N185), .A2(N186), .ZN(N12965));
    NOR2X1 U94 (.A1(N187), .A2(N188), .ZN(n12966));
    NOR2X1 U95 (.A1(N189), .A2(N190), .ZN(n12967));
    NOR2X1 U96 (.A1(N191), .A2(N192), .ZN(n12968));
    NOR2X1 U97 (.A1(N193), .A2(N194), .ZN(N12969));
    NANDX1 U98 (.A1(N195), .A2(N196), .ZN(n12970));
    NANDX1 U99 (.A1(N197), .A2(N198), .ZN(n12971));
    NOR2X1 U100 (.A1(N199), .A2(N200), .ZN(n12972));
    NOR2X1 U101 (.A1(N201), .A2(N202), .ZN(N12973));
    NOR2X1 U102 (.A1(N203), .A2(N204), .ZN(n12974));
    NANDX1 U103 (.A1(N205), .A2(N206), .ZN(n12975));
    NANDX1 U104 (.A1(N207), .A2(N208), .ZN(n12976));
    NANDX1 U105 (.A1(N209), .A2(N210), .ZN(n12977));
    NOR2X1 U106 (.A1(N211), .A2(N212), .ZN(n12978));
    NANDX1 U107 (.A1(N213), .A2(N214), .ZN(n12979));
    NOR2X1 U108 (.A1(N215), .A2(N216), .ZN(N12980));
    NOR2X1 U109 (.A1(N217), .A2(N218), .ZN(N12981));
    NOR2X1 U110 (.A1(N219), .A2(N220), .ZN(n12982));
    NANDX1 U111 (.A1(N221), .A2(N222), .ZN(n12983));
    NOR2X1 U112 (.A1(N223), .A2(N224), .ZN(n12984));
    NOR2X1 U113 (.A1(N225), .A2(N226), .ZN(n12985));
    NANDX1 U114 (.A1(N227), .A2(N228), .ZN(n12986));
    NANDX1 U115 (.A1(N229), .A2(N230), .ZN(n12987));
    NANDX1 U116 (.A1(N231), .A2(N232), .ZN(n12988));
    NOR2X1 U117 (.A1(N233), .A2(N234), .ZN(n12989));
    NANDX1 U118 (.A1(N235), .A2(N236), .ZN(n12990));
    NOR2X1 U119 (.A1(N237), .A2(N238), .ZN(N12991));
    NANDX1 U120 (.A1(N239), .A2(N240), .ZN(n12992));
    NANDX1 U121 (.A1(N241), .A2(N242), .ZN(n12993));
    NANDX1 U122 (.A1(N243), .A2(N244), .ZN(n12994));
    NANDX1 U123 (.A1(N245), .A2(N246), .ZN(N12995));
    NANDX1 U124 (.A1(N247), .A2(N248), .ZN(N12996));
    NANDX1 U125 (.A1(N249), .A2(N250), .ZN(n12997));
    NANDX1 U126 (.A1(N251), .A2(N252), .ZN(n12998));
    NANDX1 U127 (.A1(N253), .A2(N254), .ZN(n12999));
    NANDX1 U128 (.A1(N255), .A2(N256), .ZN(n13000));
    NANDX1 U129 (.A1(N257), .A2(N258), .ZN(n13001));
    NOR2X1 U130 (.A1(N259), .A2(N260), .ZN(n13002));
    NANDX1 U131 (.A1(N261), .A2(N262), .ZN(n13003));
    NANDX1 U132 (.A1(N263), .A2(N264), .ZN(n13004));
    NOR2X1 U133 (.A1(N265), .A2(N266), .ZN(n13005));
    NANDX1 U134 (.A1(N267), .A2(N268), .ZN(n13006));
    NOR2X1 U135 (.A1(N269), .A2(N270), .ZN(n13007));
    NANDX1 U136 (.A1(N271), .A2(N272), .ZN(N13008));
    NANDX1 U137 (.A1(N273), .A2(N274), .ZN(n13009));
    NOR2X1 U138 (.A1(N275), .A2(N276), .ZN(n13010));
    NOR2X1 U139 (.A1(N277), .A2(N278), .ZN(n13011));
    NANDX1 U140 (.A1(N279), .A2(N280), .ZN(n13012));
    NOR2X1 U141 (.A1(N281), .A2(N282), .ZN(n13013));
    NANDX1 U142 (.A1(N283), .A2(N284), .ZN(n13014));
    NANDX1 U143 (.A1(N285), .A2(N286), .ZN(N13015));
    NANDX1 U144 (.A1(N287), .A2(N288), .ZN(n13016));
    NOR2X1 U145 (.A1(N289), .A2(N290), .ZN(n13017));
    NOR2X1 U146 (.A1(N291), .A2(N292), .ZN(n13018));
    NOR2X1 U147 (.A1(N293), .A2(N294), .ZN(n13019));
    NANDX1 U148 (.A1(N295), .A2(N296), .ZN(n13020));
    NOR2X1 U149 (.A1(N297), .A2(N298), .ZN(N13021));
    NANDX1 U150 (.A1(N299), .A2(N300), .ZN(n13022));
    NOR2X1 U151 (.A1(N301), .A2(N302), .ZN(N13023));
    NANDX1 U152 (.A1(N303), .A2(N304), .ZN(N13024));
    NOR2X1 U153 (.A1(N305), .A2(N306), .ZN(n13025));
    NANDX1 U154 (.A1(N307), .A2(N308), .ZN(n13026));
    NOR2X1 U155 (.A1(N309), .A2(N310), .ZN(n13027));
    NANDX1 U156 (.A1(N311), .A2(N312), .ZN(N13028));
    NANDX1 U157 (.A1(N313), .A2(N314), .ZN(n13029));
    NANDX1 U158 (.A1(N315), .A2(N316), .ZN(n13030));
    NANDX1 U159 (.A1(N317), .A2(N318), .ZN(n13031));
    NOR2X1 U160 (.A1(N319), .A2(N320), .ZN(n13032));
    NOR2X1 U161 (.A1(N321), .A2(N322), .ZN(N13033));
    NOR2X1 U162 (.A1(N323), .A2(N324), .ZN(n13034));
    NANDX1 U163 (.A1(N325), .A2(N326), .ZN(N13035));
    NOR2X1 U164 (.A1(N327), .A2(N328), .ZN(n13036));
    NANDX1 U165 (.A1(N329), .A2(N330), .ZN(n13037));
    NOR2X1 U166 (.A1(N331), .A2(N332), .ZN(n13038));
    NOR2X1 U167 (.A1(N333), .A2(N334), .ZN(n13039));
    NOR2X1 U168 (.A1(N335), .A2(N336), .ZN(N13040));
    NOR2X1 U169 (.A1(N337), .A2(N338), .ZN(n13041));
    NOR2X1 U170 (.A1(N339), .A2(N340), .ZN(n13042));
    NANDX1 U171 (.A1(N341), .A2(N342), .ZN(N13043));
    NOR2X1 U172 (.A1(N343), .A2(N344), .ZN(n13044));
    NANDX1 U173 (.A1(N345), .A2(N346), .ZN(n13045));
    NANDX1 U174 (.A1(N347), .A2(N348), .ZN(n13046));
    NANDX1 U175 (.A1(N349), .A2(N350), .ZN(n13047));
    NANDX1 U176 (.A1(N351), .A2(N352), .ZN(n13048));
    NANDX1 U177 (.A1(N353), .A2(N354), .ZN(n13049));
    NOR2X1 U178 (.A1(N355), .A2(N356), .ZN(n13050));
    NOR2X1 U179 (.A1(N357), .A2(N358), .ZN(n13051));
    NANDX1 U180 (.A1(N359), .A2(N360), .ZN(n13052));
    NANDX1 U181 (.A1(N361), .A2(N362), .ZN(n13053));
    NOR2X1 U182 (.A1(N363), .A2(N364), .ZN(n13054));
    NANDX1 U183 (.A1(N365), .A2(N366), .ZN(n13055));
    NANDX1 U184 (.A1(N367), .A2(N368), .ZN(n13056));
    NOR2X1 U185 (.A1(N369), .A2(N370), .ZN(n13057));
    NANDX1 U186 (.A1(N371), .A2(N372), .ZN(n13058));
    NOR2X1 U187 (.A1(N373), .A2(N374), .ZN(n13059));
    NANDX1 U188 (.A1(N375), .A2(N376), .ZN(n13060));
    NANDX1 U189 (.A1(N377), .A2(N378), .ZN(n13061));
    NANDX1 U190 (.A1(N379), .A2(N380), .ZN(n13062));
    NANDX1 U191 (.A1(N381), .A2(N382), .ZN(n13063));
    NANDX1 U192 (.A1(N383), .A2(N384), .ZN(n13064));
    NOR2X1 U193 (.A1(N385), .A2(N386), .ZN(N13065));
    NOR2X1 U194 (.A1(N387), .A2(N388), .ZN(n13066));
    NANDX1 U195 (.A1(N389), .A2(N390), .ZN(n13067));
    NANDX1 U196 (.A1(N391), .A2(N392), .ZN(n13068));
    NOR2X1 U197 (.A1(N393), .A2(N394), .ZN(n13069));
    NANDX1 U198 (.A1(N395), .A2(N396), .ZN(n13070));
    NOR2X1 U199 (.A1(N397), .A2(N398), .ZN(N13071));
    NOR2X1 U200 (.A1(N399), .A2(N400), .ZN(n13072));
    NANDX1 U201 (.A1(N401), .A2(N402), .ZN(n13073));
    NANDX1 U202 (.A1(N403), .A2(N404), .ZN(n13074));
    NANDX1 U203 (.A1(N405), .A2(N406), .ZN(n13075));
    NOR2X1 U204 (.A1(N407), .A2(N408), .ZN(n13076));
    NOR2X1 U205 (.A1(N409), .A2(N410), .ZN(n13077));
    NOR2X1 U206 (.A1(N411), .A2(N412), .ZN(n13078));
    NOR2X1 U207 (.A1(N413), .A2(N414), .ZN(n13079));
    NOR2X1 U208 (.A1(N415), .A2(N416), .ZN(n13080));
    NOR2X1 U209 (.A1(N417), .A2(N418), .ZN(n13081));
    NOR2X1 U210 (.A1(N419), .A2(N420), .ZN(n13082));
    NANDX1 U211 (.A1(N421), .A2(N422), .ZN(n13083));
    NANDX1 U212 (.A1(N423), .A2(N424), .ZN(N13084));
    NANDX1 U213 (.A1(N425), .A2(N426), .ZN(n13085));
    NOR2X1 U214 (.A1(N427), .A2(N428), .ZN(n13086));
    NOR2X1 U215 (.A1(N429), .A2(N430), .ZN(n13087));
    NANDX1 U216 (.A1(N431), .A2(N432), .ZN(n13088));
    NOR2X1 U217 (.A1(N433), .A2(N434), .ZN(n13089));
    NANDX1 U218 (.A1(N435), .A2(N436), .ZN(n13090));
    NOR2X1 U219 (.A1(N437), .A2(N438), .ZN(n13091));
    NANDX1 U220 (.A1(N439), .A2(N440), .ZN(n13092));
    NOR2X1 U221 (.A1(N441), .A2(N442), .ZN(n13093));
    NANDX1 U222 (.A1(N443), .A2(N444), .ZN(n13094));
    NOR2X1 U223 (.A1(N445), .A2(N446), .ZN(n13095));
    NOR2X1 U224 (.A1(N447), .A2(N448), .ZN(N13096));
    NANDX1 U225 (.A1(N449), .A2(N450), .ZN(n13097));
    NANDX1 U226 (.A1(N451), .A2(N452), .ZN(n13098));
    NOR2X1 U227 (.A1(N453), .A2(N454), .ZN(n13099));
    NOR2X1 U228 (.A1(N455), .A2(N456), .ZN(n13100));
    NANDX1 U229 (.A1(N457), .A2(N458), .ZN(n13101));
    NOR2X1 U230 (.A1(N459), .A2(N460), .ZN(n13102));
    NOR2X1 U231 (.A1(N461), .A2(N462), .ZN(n13103));
    NOR2X1 U232 (.A1(N463), .A2(N464), .ZN(n13104));
    NANDX1 U233 (.A1(N465), .A2(N466), .ZN(n13105));
    NANDX1 U234 (.A1(N467), .A2(N468), .ZN(n13106));
    NANDX1 U235 (.A1(N469), .A2(N470), .ZN(n13107));
    NOR2X1 U236 (.A1(N471), .A2(N472), .ZN(n13108));
    NOR2X1 U237 (.A1(N473), .A2(N474), .ZN(n13109));
    NANDX1 U238 (.A1(N475), .A2(N476), .ZN(N13110));
    NOR2X1 U239 (.A1(N477), .A2(N478), .ZN(n13111));
    NOR2X1 U240 (.A1(N479), .A2(N480), .ZN(n13112));
    NANDX1 U241 (.A1(N481), .A2(N482), .ZN(n13113));
    NANDX1 U242 (.A1(N483), .A2(N484), .ZN(n13114));
    NOR2X1 U243 (.A1(N485), .A2(N486), .ZN(n13115));
    NOR2X1 U244 (.A1(N487), .A2(N488), .ZN(n13116));
    NOR2X1 U245 (.A1(N489), .A2(N490), .ZN(n13117));
    NOR2X1 U246 (.A1(N491), .A2(N492), .ZN(N13118));
    NANDX1 U247 (.A1(N493), .A2(N494), .ZN(n13119));
    NOR2X1 U248 (.A1(N495), .A2(N496), .ZN(N13120));
    NANDX1 U249 (.A1(N497), .A2(N498), .ZN(n13121));
    NANDX1 U250 (.A1(N499), .A2(N500), .ZN(n13122));
    NANDX1 U251 (.A1(N501), .A2(N502), .ZN(N13123));
    NOR2X1 U252 (.A1(N503), .A2(N504), .ZN(N13124));
    NOR2X1 U253 (.A1(N505), .A2(N506), .ZN(n13125));
    NANDX1 U254 (.A1(N507), .A2(N508), .ZN(n13126));
    NOR2X1 U255 (.A1(N509), .A2(N510), .ZN(n13127));
    NOR2X1 U256 (.A1(N511), .A2(N512), .ZN(n13128));
    NOR2X1 U257 (.A1(N513), .A2(N514), .ZN(n13129));
    NOR2X1 U258 (.A1(N515), .A2(N516), .ZN(n13130));
    NOR2X1 U259 (.A1(N517), .A2(N518), .ZN(n13131));
    NANDX1 U260 (.A1(N519), .A2(N520), .ZN(N13132));
    NOR2X1 U261 (.A1(N521), .A2(N522), .ZN(n13133));
    NOR2X1 U262 (.A1(N523), .A2(N524), .ZN(n13134));
    NOR2X1 U263 (.A1(N525), .A2(N526), .ZN(n13135));
    NOR2X1 U264 (.A1(N527), .A2(N528), .ZN(n13136));
    NOR2X1 U265 (.A1(N529), .A2(N530), .ZN(n13137));
    NANDX1 U266 (.A1(N531), .A2(N532), .ZN(n13138));
    NOR2X1 U267 (.A1(N533), .A2(N534), .ZN(n13139));
    NOR2X1 U268 (.A1(N535), .A2(N536), .ZN(n13140));
    NOR2X1 U269 (.A1(N537), .A2(N538), .ZN(n13141));
    NOR2X1 U270 (.A1(N539), .A2(N540), .ZN(n13142));
    NOR2X1 U271 (.A1(N541), .A2(N542), .ZN(n13143));
    NANDX1 U272 (.A1(N543), .A2(N544), .ZN(N13144));
    NANDX1 U273 (.A1(N545), .A2(N546), .ZN(n13145));
    NOR2X1 U274 (.A1(N547), .A2(N548), .ZN(n13146));
    NOR2X1 U275 (.A1(N549), .A2(N550), .ZN(n13147));
    NANDX1 U276 (.A1(N551), .A2(N552), .ZN(n13148));
    NANDX1 U277 (.A1(N553), .A2(N554), .ZN(n13149));
    NANDX1 U278 (.A1(N555), .A2(N556), .ZN(n13150));
    NANDX1 U279 (.A1(N557), .A2(N558), .ZN(n13151));
    NOR2X1 U280 (.A1(N559), .A2(N560), .ZN(n13152));
    NANDX1 U281 (.A1(N561), .A2(N562), .ZN(n13153));
    NOR2X1 U282 (.A1(N563), .A2(N564), .ZN(N13154));
    NOR2X1 U283 (.A1(N565), .A2(N566), .ZN(n13155));
    NANDX1 U284 (.A1(N567), .A2(N568), .ZN(n13156));
    NANDX1 U285 (.A1(N569), .A2(N570), .ZN(N13157));
    NANDX1 U286 (.A1(N571), .A2(N572), .ZN(n13158));
    NANDX1 U287 (.A1(N573), .A2(N574), .ZN(n13159));
    NOR2X1 U288 (.A1(N575), .A2(N576), .ZN(n13160));
    NANDX1 U289 (.A1(N577), .A2(N578), .ZN(n13161));
    NANDX1 U290 (.A1(N579), .A2(N580), .ZN(n13162));
    NANDX1 U291 (.A1(N581), .A2(N582), .ZN(n13163));
    NOR2X1 U292 (.A1(N583), .A2(N584), .ZN(n13164));
    NOR2X1 U293 (.A1(N585), .A2(N586), .ZN(N13165));
    NANDX1 U294 (.A1(N587), .A2(N588), .ZN(n13166));
    NOR2X1 U295 (.A1(N589), .A2(N590), .ZN(n13167));
    NOR2X1 U296 (.A1(N591), .A2(N592), .ZN(N13168));
    NOR2X1 U297 (.A1(N593), .A2(N594), .ZN(n13169));
    NOR2X1 U298 (.A1(N595), .A2(N596), .ZN(N13170));
    NOR2X1 U299 (.A1(N597), .A2(N598), .ZN(n13171));
    NOR2X1 U300 (.A1(N599), .A2(N600), .ZN(n13172));
    NOR2X1 U301 (.A1(N601), .A2(N602), .ZN(n13173));
    NOR2X1 U302 (.A1(N603), .A2(N604), .ZN(n13174));
    NOR2X1 U303 (.A1(N605), .A2(N606), .ZN(n13175));
    NANDX1 U304 (.A1(N607), .A2(N608), .ZN(n13176));
    NANDX1 U305 (.A1(N609), .A2(N610), .ZN(n13177));
    NOR2X1 U306 (.A1(N611), .A2(N612), .ZN(n13178));
    NANDX1 U307 (.A1(N613), .A2(N614), .ZN(n13179));
    NOR2X1 U308 (.A1(N615), .A2(N616), .ZN(n13180));
    NANDX1 U309 (.A1(N617), .A2(N618), .ZN(n13181));
    NOR2X1 U310 (.A1(N619), .A2(N620), .ZN(N13182));
    NOR2X1 U311 (.A1(N621), .A2(N622), .ZN(n13183));
    NOR2X1 U312 (.A1(N623), .A2(N624), .ZN(n13184));
    NANDX1 U313 (.A1(N625), .A2(N626), .ZN(n13185));
    NANDX1 U314 (.A1(N627), .A2(N628), .ZN(n13186));
    NOR2X1 U315 (.A1(N629), .A2(N630), .ZN(n13187));
    NOR2X1 U316 (.A1(N631), .A2(N632), .ZN(n13188));
    NOR2X1 U317 (.A1(N633), .A2(N634), .ZN(N13189));
    NANDX1 U318 (.A1(N635), .A2(N636), .ZN(n13190));
    NOR2X1 U319 (.A1(N637), .A2(N638), .ZN(n13191));
    NANDX1 U320 (.A1(N639), .A2(N640), .ZN(n13192));
    NANDX1 U321 (.A1(N641), .A2(N642), .ZN(n13193));
    NOR2X1 U322 (.A1(N643), .A2(N644), .ZN(n13194));
    NANDX1 U323 (.A1(N645), .A2(N646), .ZN(n13195));
    NANDX1 U324 (.A1(N647), .A2(N648), .ZN(n13196));
    NANDX1 U325 (.A1(N649), .A2(N650), .ZN(n13197));
    NANDX1 U326 (.A1(N651), .A2(N652), .ZN(n13198));
    NANDX1 U327 (.A1(N653), .A2(N654), .ZN(n13199));
    NOR2X1 U328 (.A1(N655), .A2(N656), .ZN(N13200));
    NANDX1 U329 (.A1(N657), .A2(N658), .ZN(n13201));
    NANDX1 U330 (.A1(N659), .A2(N660), .ZN(n13202));
    NOR2X1 U331 (.A1(N661), .A2(N662), .ZN(n13203));
    NANDX1 U332 (.A1(N663), .A2(N664), .ZN(n13204));
    NANDX1 U333 (.A1(N665), .A2(N666), .ZN(n13205));
    NOR2X1 U334 (.A1(N667), .A2(N668), .ZN(N13206));
    NANDX1 U335 (.A1(N669), .A2(N670), .ZN(n13207));
    NOR2X1 U336 (.A1(N671), .A2(N672), .ZN(n13208));
    NOR2X1 U337 (.A1(N673), .A2(N674), .ZN(n13209));
    NOR2X1 U338 (.A1(N675), .A2(N676), .ZN(n13210));
    NOR2X1 U339 (.A1(N677), .A2(N678), .ZN(N13211));
    NOR2X1 U340 (.A1(N679), .A2(N680), .ZN(n13212));
    NOR2X1 U341 (.A1(N681), .A2(N682), .ZN(n13213));
    NANDX1 U342 (.A1(N683), .A2(N684), .ZN(n13214));
    NOR2X1 U343 (.A1(N685), .A2(N686), .ZN(n13215));
    NANDX1 U344 (.A1(N687), .A2(N688), .ZN(n13216));
    NOR2X1 U345 (.A1(N689), .A2(N690), .ZN(N13217));
    NOR2X1 U346 (.A1(N691), .A2(N692), .ZN(n13218));
    NOR2X1 U347 (.A1(N693), .A2(N694), .ZN(n13219));
    NOR2X1 U348 (.A1(N695), .A2(N696), .ZN(n13220));
    NOR2X1 U349 (.A1(N697), .A2(N698), .ZN(n13221));
    NOR2X1 U350 (.A1(N699), .A2(N700), .ZN(n13222));
    NANDX1 U351 (.A1(N701), .A2(N702), .ZN(n13223));
    NANDX1 U352 (.A1(N703), .A2(N704), .ZN(n13224));
    NOR2X1 U353 (.A1(N705), .A2(N706), .ZN(N13225));
    NANDX1 U354 (.A1(N707), .A2(N708), .ZN(n13226));
    NOR2X1 U355 (.A1(N709), .A2(N710), .ZN(n13227));
    NOR2X1 U356 (.A1(N711), .A2(N712), .ZN(N13228));
    NOR2X1 U357 (.A1(N713), .A2(N714), .ZN(n13229));
    NANDX1 U358 (.A1(N715), .A2(N716), .ZN(n13230));
    NOR2X1 U359 (.A1(N717), .A2(N718), .ZN(n13231));
    NOR2X1 U360 (.A1(N719), .A2(N720), .ZN(n13232));
    NOR2X1 U361 (.A1(N721), .A2(N722), .ZN(N13233));
    NOR2X1 U362 (.A1(N723), .A2(N724), .ZN(n13234));
    NANDX1 U363 (.A1(N725), .A2(N726), .ZN(n13235));
    NANDX1 U364 (.A1(N727), .A2(N728), .ZN(n13236));
    NANDX1 U365 (.A1(N729), .A2(N730), .ZN(n13237));
    NOR2X1 U366 (.A1(N731), .A2(N732), .ZN(n13238));
    NOR2X1 U367 (.A1(N733), .A2(N734), .ZN(n13239));
    NANDX1 U368 (.A1(N735), .A2(N736), .ZN(n13240));
    NOR2X1 U369 (.A1(N737), .A2(N738), .ZN(N13241));
    NOR2X1 U370 (.A1(N739), .A2(N740), .ZN(N13242));
    NANDX1 U371 (.A1(N741), .A2(N742), .ZN(n13243));
    NANDX1 U372 (.A1(N743), .A2(N744), .ZN(n13244));
    NANDX1 U373 (.A1(N745), .A2(N746), .ZN(n13245));
    NOR2X1 U374 (.A1(N747), .A2(N748), .ZN(n13246));
    NOR2X1 U375 (.A1(N749), .A2(N750), .ZN(n13247));
    NANDX1 U376 (.A1(N751), .A2(N752), .ZN(n13248));
    NOR2X1 U377 (.A1(N753), .A2(N754), .ZN(n13249));
    NOR2X1 U378 (.A1(N755), .A2(N756), .ZN(N13250));
    NANDX1 U379 (.A1(N757), .A2(N758), .ZN(n13251));
    NOR2X1 U380 (.A1(N759), .A2(N760), .ZN(n13252));
    NANDX1 U381 (.A1(N761), .A2(N762), .ZN(n13253));
    NANDX1 U382 (.A1(N763), .A2(N764), .ZN(n13254));
    NANDX1 U383 (.A1(N765), .A2(N766), .ZN(n13255));
    NANDX1 U384 (.A1(N767), .A2(N768), .ZN(n13256));
    NOR2X1 U385 (.A1(N769), .A2(N770), .ZN(N13257));
    NANDX1 U386 (.A1(N771), .A2(N772), .ZN(n13258));
    NANDX1 U387 (.A1(N773), .A2(N774), .ZN(n13259));
    NOR2X1 U388 (.A1(N775), .A2(N776), .ZN(n13260));
    NOR2X1 U389 (.A1(N777), .A2(N778), .ZN(n13261));
    NANDX1 U390 (.A1(N779), .A2(N780), .ZN(n13262));
    NOR2X1 U391 (.A1(N781), .A2(N782), .ZN(n13263));
    NOR2X1 U392 (.A1(N783), .A2(N784), .ZN(n13264));
    NOR2X1 U393 (.A1(N785), .A2(N786), .ZN(n13265));
    NOR2X1 U394 (.A1(N787), .A2(N788), .ZN(n13266));
    NOR2X1 U395 (.A1(N789), .A2(N790), .ZN(n13267));
    NANDX1 U396 (.A1(N791), .A2(N792), .ZN(n13268));
    NOR2X1 U397 (.A1(N793), .A2(N794), .ZN(n13269));
    NOR2X1 U398 (.A1(N795), .A2(N796), .ZN(n13270));
    NOR2X1 U399 (.A1(N797), .A2(N798), .ZN(n13271));
    NANDX1 U400 (.A1(N799), .A2(N800), .ZN(n13272));
    NOR2X1 U401 (.A1(N801), .A2(N802), .ZN(n13273));
    NOR2X1 U402 (.A1(N803), .A2(N804), .ZN(n13274));
    NOR2X1 U403 (.A1(N805), .A2(N806), .ZN(n13275));
    NOR2X1 U404 (.A1(N807), .A2(N808), .ZN(N13276));
    NOR2X1 U405 (.A1(N809), .A2(N810), .ZN(N13277));
    NOR2X1 U406 (.A1(N811), .A2(N812), .ZN(n13278));
    NANDX1 U407 (.A1(N813), .A2(N814), .ZN(n13279));
    NOR2X1 U408 (.A1(N815), .A2(N816), .ZN(n13280));
    NANDX1 U409 (.A1(N817), .A2(N818), .ZN(n13281));
    NANDX1 U410 (.A1(N819), .A2(N820), .ZN(n13282));
    NANDX1 U411 (.A1(N821), .A2(N822), .ZN(N13283));
    NOR2X1 U412 (.A1(N823), .A2(N824), .ZN(n13284));
    NOR2X1 U413 (.A1(N825), .A2(N826), .ZN(n13285));
    NOR2X1 U414 (.A1(N827), .A2(N828), .ZN(n13286));
    NANDX1 U415 (.A1(N829), .A2(N830), .ZN(n13287));
    NOR2X1 U416 (.A1(N831), .A2(N832), .ZN(n13288));
    NOR2X1 U417 (.A1(N833), .A2(N834), .ZN(n13289));
    NANDX1 U418 (.A1(N835), .A2(N836), .ZN(n13290));
    NOR2X1 U419 (.A1(N837), .A2(N838), .ZN(n13291));
    NOR2X1 U420 (.A1(N839), .A2(N840), .ZN(n13292));
    NOR2X1 U421 (.A1(N841), .A2(N842), .ZN(n13293));
    NANDX1 U422 (.A1(N843), .A2(N844), .ZN(n13294));
    NANDX1 U423 (.A1(N845), .A2(N846), .ZN(n13295));
    NOR2X1 U424 (.A1(N847), .A2(N848), .ZN(n13296));
    NANDX1 U425 (.A1(N849), .A2(N850), .ZN(n13297));
    NANDX1 U426 (.A1(N851), .A2(N852), .ZN(n13298));
    NANDX1 U427 (.A1(N853), .A2(N854), .ZN(n13299));
    NANDX1 U428 (.A1(N855), .A2(N856), .ZN(n13300));
    NANDX1 U429 (.A1(N857), .A2(N858), .ZN(n13301));
    NOR2X1 U430 (.A1(N859), .A2(N860), .ZN(n13302));
    NOR2X1 U431 (.A1(N861), .A2(N862), .ZN(n13303));
    NANDX1 U432 (.A1(N863), .A2(N864), .ZN(n13304));
    NOR2X1 U433 (.A1(N865), .A2(N866), .ZN(n13305));
    NOR2X1 U434 (.A1(N867), .A2(N868), .ZN(n13306));
    NANDX1 U435 (.A1(N869), .A2(N870), .ZN(N13307));
    NOR2X1 U436 (.A1(N871), .A2(N872), .ZN(n13308));
    NANDX1 U437 (.A1(N873), .A2(N874), .ZN(N13309));
    NANDX1 U438 (.A1(N875), .A2(N876), .ZN(N13310));
    NOR2X1 U439 (.A1(N877), .A2(N878), .ZN(n13311));
    NOR2X1 U440 (.A1(N879), .A2(N880), .ZN(n13312));
    NOR2X1 U441 (.A1(N881), .A2(N882), .ZN(n13313));
    NANDX1 U442 (.A1(N883), .A2(N884), .ZN(n13314));
    NOR2X1 U443 (.A1(N885), .A2(N886), .ZN(n13315));
    NOR2X1 U444 (.A1(N887), .A2(N888), .ZN(n13316));
    NOR2X1 U445 (.A1(N889), .A2(N890), .ZN(n13317));
    NANDX1 U446 (.A1(N891), .A2(N892), .ZN(n13318));
    NOR2X1 U447 (.A1(N893), .A2(N894), .ZN(n13319));
    NOR2X1 U448 (.A1(N895), .A2(N896), .ZN(n13320));
    NOR2X1 U449 (.A1(N897), .A2(N898), .ZN(n13321));
    NOR2X1 U450 (.A1(N899), .A2(N900), .ZN(n13322));
    NOR2X1 U451 (.A1(N901), .A2(N902), .ZN(n13323));
    NANDX1 U452 (.A1(N903), .A2(N904), .ZN(n13324));
    NANDX1 U453 (.A1(N905), .A2(N906), .ZN(n13325));
    NANDX1 U454 (.A1(N907), .A2(N908), .ZN(N13326));
    NANDX1 U455 (.A1(N909), .A2(N910), .ZN(N13327));
    NOR2X1 U456 (.A1(N911), .A2(N912), .ZN(n13328));
    NOR2X1 U457 (.A1(N913), .A2(N914), .ZN(n13329));
    NANDX1 U458 (.A1(N915), .A2(N916), .ZN(N13330));
    NOR2X1 U459 (.A1(N917), .A2(N918), .ZN(n13331));
    NANDX1 U460 (.A1(N919), .A2(N920), .ZN(n13332));
    NANDX1 U461 (.A1(N921), .A2(N922), .ZN(n13333));
    NOR2X1 U462 (.A1(N923), .A2(N924), .ZN(n13334));
    NANDX1 U463 (.A1(N925), .A2(N926), .ZN(n13335));
    NANDX1 U464 (.A1(N927), .A2(N928), .ZN(n13336));
    NANDX1 U465 (.A1(N929), .A2(N930), .ZN(n13337));
    NOR2X1 U466 (.A1(N931), .A2(N932), .ZN(n13338));
    NANDX1 U467 (.A1(N933), .A2(N934), .ZN(N13339));
    NOR2X1 U468 (.A1(N935), .A2(N936), .ZN(n13340));
    NANDX1 U469 (.A1(N937), .A2(N938), .ZN(n13341));
    NANDX1 U470 (.A1(N939), .A2(N940), .ZN(N13342));
    NOR2X1 U471 (.A1(N941), .A2(N942), .ZN(n13343));
    NANDX1 U472 (.A1(N943), .A2(N944), .ZN(n13344));
    NANDX1 U473 (.A1(N945), .A2(N946), .ZN(n13345));
    NOR2X1 U474 (.A1(N947), .A2(N948), .ZN(n13346));
    NANDX1 U475 (.A1(N949), .A2(N950), .ZN(n13347));
    NANDX1 U476 (.A1(N951), .A2(N952), .ZN(N13348));
    NANDX1 U477 (.A1(N953), .A2(N954), .ZN(n13349));
    NANDX1 U478 (.A1(N955), .A2(N956), .ZN(n13350));
    NANDX1 U479 (.A1(N957), .A2(N958), .ZN(n13351));
    NOR2X1 U480 (.A1(N959), .A2(N960), .ZN(n13352));
    NOR2X1 U481 (.A1(N961), .A2(N962), .ZN(N13353));
    NANDX1 U482 (.A1(N963), .A2(N964), .ZN(n13354));
    NANDX1 U483 (.A1(N965), .A2(N966), .ZN(n13355));
    NANDX1 U484 (.A1(N967), .A2(N968), .ZN(n13356));
    NANDX1 U485 (.A1(N969), .A2(N970), .ZN(n13357));
    NOR2X1 U486 (.A1(N971), .A2(N972), .ZN(n13358));
    NOR2X1 U487 (.A1(N973), .A2(N974), .ZN(n13359));
    NANDX1 U488 (.A1(N975), .A2(N976), .ZN(N13360));
    NANDX1 U489 (.A1(N977), .A2(N978), .ZN(N13361));
    NOR2X1 U490 (.A1(N979), .A2(N980), .ZN(N13362));
    NANDX1 U491 (.A1(N981), .A2(N982), .ZN(n13363));
    NOR2X1 U492 (.A1(N983), .A2(N984), .ZN(n13364));
    NOR2X1 U493 (.A1(N985), .A2(N986), .ZN(n13365));
    NOR2X1 U494 (.A1(N987), .A2(N988), .ZN(n13366));
    NANDX1 U495 (.A1(N989), .A2(N990), .ZN(n13367));
    NANDX1 U496 (.A1(N991), .A2(N992), .ZN(n13368));
    NOR2X1 U497 (.A1(N993), .A2(N994), .ZN(N13369));
    NOR2X1 U498 (.A1(N995), .A2(N996), .ZN(n13370));
    NANDX1 U499 (.A1(N997), .A2(N998), .ZN(n13371));
    NOR2X1 U500 (.A1(N999), .A2(N1000), .ZN(n13372));
    NOR2X1 U501 (.A1(N1001), .A2(N1002), .ZN(N13373));
    NANDX1 U502 (.A1(N1003), .A2(N1004), .ZN(n13374));
    NANDX1 U503 (.A1(N1005), .A2(N1006), .ZN(n13375));
    NANDX1 U504 (.A1(N1007), .A2(N1008), .ZN(N13376));
    NANDX1 U505 (.A1(N1009), .A2(N1010), .ZN(N13377));
    NANDX1 U506 (.A1(N1011), .A2(N1012), .ZN(n13378));
    NOR2X1 U507 (.A1(N1013), .A2(N1014), .ZN(n13379));
    NANDX1 U508 (.A1(N1015), .A2(N1016), .ZN(n13380));
    NOR2X1 U509 (.A1(N1017), .A2(N1018), .ZN(N13381));
    NANDX1 U510 (.A1(N1019), .A2(N1020), .ZN(n13382));
    NANDX1 U511 (.A1(N1021), .A2(N1022), .ZN(n13383));
    NOR2X1 U512 (.A1(N1023), .A2(N1024), .ZN(n13384));
    NOR2X1 U513 (.A1(N1025), .A2(N1026), .ZN(n13385));
    NOR2X1 U514 (.A1(N1027), .A2(N1028), .ZN(n13386));
    NOR2X1 U515 (.A1(N1029), .A2(N1030), .ZN(n13387));
    NANDX1 U516 (.A1(N1031), .A2(N1032), .ZN(n13388));
    NOR2X1 U517 (.A1(N1033), .A2(N1034), .ZN(n13389));
    NOR2X1 U518 (.A1(N1035), .A2(N1036), .ZN(n13390));
    NANDX1 U519 (.A1(N1037), .A2(N1038), .ZN(n13391));
    NOR2X1 U520 (.A1(N1039), .A2(N1040), .ZN(n13392));
    NOR2X1 U521 (.A1(N1041), .A2(N1042), .ZN(n13393));
    NOR2X1 U522 (.A1(N1043), .A2(N1044), .ZN(n13394));
    NOR2X1 U523 (.A1(N1045), .A2(N1046), .ZN(n13395));
    NOR2X1 U524 (.A1(N1047), .A2(N1048), .ZN(N13396));
    NOR2X1 U525 (.A1(N1049), .A2(N1050), .ZN(n13397));
    NOR2X1 U526 (.A1(N1051), .A2(N1052), .ZN(n13398));
    NOR2X1 U527 (.A1(N1053), .A2(N1054), .ZN(n13399));
    NOR2X1 U528 (.A1(N1055), .A2(N1056), .ZN(n13400));
    NOR2X1 U529 (.A1(N1057), .A2(N1058), .ZN(n13401));
    NANDX1 U530 (.A1(N1059), .A2(N1060), .ZN(n13402));
    NOR2X1 U531 (.A1(N1061), .A2(N1062), .ZN(n13403));
    NOR2X1 U532 (.A1(N1063), .A2(N1064), .ZN(n13404));
    NANDX1 U533 (.A1(N1065), .A2(N1066), .ZN(n13405));
    NOR2X1 U534 (.A1(N1067), .A2(N1068), .ZN(n13406));
    NANDX1 U535 (.A1(N1069), .A2(N1070), .ZN(n13407));
    NOR2X1 U536 (.A1(N1071), .A2(N1072), .ZN(N13408));
    NANDX1 U537 (.A1(N1073), .A2(N1074), .ZN(n13409));
    NANDX1 U538 (.A1(N1075), .A2(N1076), .ZN(N13410));
    NANDX1 U539 (.A1(N1077), .A2(N1078), .ZN(n13411));
    NANDX1 U540 (.A1(N1079), .A2(N1080), .ZN(n13412));
    NOR2X1 U541 (.A1(N1081), .A2(N1082), .ZN(n13413));
    NOR2X1 U542 (.A1(N1083), .A2(N1084), .ZN(n13414));
    NOR2X1 U543 (.A1(N1085), .A2(N1086), .ZN(N13415));
    NANDX1 U544 (.A1(N1087), .A2(N1088), .ZN(n13416));
    NOR2X1 U545 (.A1(N1089), .A2(N1090), .ZN(n13417));
    NOR2X1 U546 (.A1(N1091), .A2(N1092), .ZN(n13418));
    NOR2X1 U547 (.A1(N1093), .A2(N1094), .ZN(n13419));
    NANDX1 U548 (.A1(N1095), .A2(N1096), .ZN(N13420));
    NOR2X1 U549 (.A1(N1097), .A2(N1098), .ZN(N13421));
    NANDX1 U550 (.A1(N1099), .A2(N1100), .ZN(n13422));
    NANDX1 U551 (.A1(N1101), .A2(N1102), .ZN(n13423));
    NOR2X1 U552 (.A1(N1103), .A2(N1104), .ZN(n13424));
    NANDX1 U553 (.A1(N1105), .A2(N1106), .ZN(n13425));
    NANDX1 U554 (.A1(N1107), .A2(N1108), .ZN(n13426));
    NOR2X1 U555 (.A1(N1109), .A2(N1110), .ZN(n13427));
    NANDX1 U556 (.A1(N1111), .A2(N1112), .ZN(n13428));
    NANDX1 U557 (.A1(N1113), .A2(N1114), .ZN(n13429));
    NOR2X1 U558 (.A1(N1115), .A2(N1116), .ZN(n13430));
    NOR2X1 U559 (.A1(N1117), .A2(N1118), .ZN(N13431));
    NOR2X1 U560 (.A1(N1119), .A2(N1120), .ZN(n13432));
    NOR2X1 U561 (.A1(N1121), .A2(N1122), .ZN(n13433));
    NOR2X1 U562 (.A1(N1123), .A2(N1124), .ZN(N13434));
    NOR2X1 U563 (.A1(N1125), .A2(N1126), .ZN(n13435));
    NANDX1 U564 (.A1(N1127), .A2(N1128), .ZN(n13436));
    NOR2X1 U565 (.A1(N1129), .A2(N1130), .ZN(n13437));
    NOR2X1 U566 (.A1(N1131), .A2(N1132), .ZN(n13438));
    NANDX1 U567 (.A1(N1133), .A2(N1134), .ZN(n13439));
    NANDX1 U568 (.A1(N1135), .A2(N1136), .ZN(n13440));
    NANDX1 U569 (.A1(N1137), .A2(N1138), .ZN(n13441));
    NANDX1 U570 (.A1(N1139), .A2(N1140), .ZN(N13442));
    NANDX1 U571 (.A1(N1141), .A2(N1142), .ZN(N13443));
    NOR2X1 U572 (.A1(N1143), .A2(N1144), .ZN(N13444));
    NANDX1 U573 (.A1(N1145), .A2(N1146), .ZN(n13445));
    NANDX1 U574 (.A1(N1147), .A2(N1148), .ZN(N13446));
    NANDX1 U575 (.A1(N1149), .A2(N1150), .ZN(n13447));
    NOR2X1 U576 (.A1(N1151), .A2(N1152), .ZN(N13448));
    NANDX1 U577 (.A1(N1153), .A2(N1154), .ZN(n13449));
    NANDX1 U578 (.A1(N1155), .A2(N1156), .ZN(n13450));
    NANDX1 U579 (.A1(N1157), .A2(N1158), .ZN(n13451));
    NANDX1 U580 (.A1(N1159), .A2(N1160), .ZN(n13452));
    NANDX1 U581 (.A1(N1161), .A2(N1162), .ZN(n13453));
    NOR2X1 U582 (.A1(N1163), .A2(N1164), .ZN(n13454));
    NANDX1 U583 (.A1(N1165), .A2(N1166), .ZN(n13455));
    NOR2X1 U584 (.A1(N1167), .A2(N1168), .ZN(N13456));
    NANDX1 U585 (.A1(N1169), .A2(N1170), .ZN(N13457));
    NANDX1 U586 (.A1(N1171), .A2(N1172), .ZN(N13458));
    NOR2X1 U587 (.A1(N1173), .A2(N1174), .ZN(n13459));
    NANDX1 U588 (.A1(N1175), .A2(N1176), .ZN(n13460));
    NOR2X1 U589 (.A1(N1177), .A2(N1178), .ZN(n13461));
    NOR2X1 U590 (.A1(N1179), .A2(N1180), .ZN(n13462));
    NANDX1 U591 (.A1(N1181), .A2(N1182), .ZN(n13463));
    NOR2X1 U592 (.A1(N1183), .A2(N1184), .ZN(n13464));
    NOR2X1 U593 (.A1(N1185), .A2(N1186), .ZN(N13465));
    NANDX1 U594 (.A1(N1187), .A2(N1188), .ZN(N13466));
    NANDX1 U595 (.A1(N1189), .A2(N1190), .ZN(n13467));
    NANDX1 U596 (.A1(N1191), .A2(N1192), .ZN(n13468));
    NANDX1 U597 (.A1(N1193), .A2(N1194), .ZN(n13469));
    NOR2X1 U598 (.A1(N1195), .A2(N1196), .ZN(n13470));
    NOR2X1 U599 (.A1(N1197), .A2(N1198), .ZN(n13471));
    NANDX1 U600 (.A1(N1199), .A2(N1200), .ZN(n13472));
    NANDX1 U601 (.A1(N1201), .A2(N1202), .ZN(n13473));
    NANDX1 U602 (.A1(N1203), .A2(N1204), .ZN(n13474));
    NANDX1 U603 (.A1(N1205), .A2(N1206), .ZN(n13475));
    NANDX1 U604 (.A1(N1207), .A2(N1208), .ZN(n13476));
    NOR2X1 U605 (.A1(N1209), .A2(N1210), .ZN(n13477));
    NOR2X1 U606 (.A1(N1211), .A2(N1212), .ZN(n13478));
    NANDX1 U607 (.A1(N1213), .A2(N1214), .ZN(n13479));
    NANDX1 U608 (.A1(N1215), .A2(N1216), .ZN(n13480));
    NANDX1 U609 (.A1(N1217), .A2(N1218), .ZN(n13481));
    NOR2X1 U610 (.A1(N1219), .A2(N1220), .ZN(N13482));
    NOR2X1 U611 (.A1(N1221), .A2(N1222), .ZN(N13483));
    NOR2X1 U612 (.A1(N1223), .A2(N1224), .ZN(n13484));
    NOR2X1 U613 (.A1(N1225), .A2(N1226), .ZN(n13485));
    NANDX1 U614 (.A1(N1227), .A2(N1228), .ZN(n13486));
    NANDX1 U615 (.A1(N1229), .A2(N1230), .ZN(n13487));
    NANDX1 U616 (.A1(N1231), .A2(N1232), .ZN(n13488));
    NANDX1 U617 (.A1(N1233), .A2(N1234), .ZN(n13489));
    NANDX1 U618 (.A1(N1235), .A2(N1236), .ZN(N13490));
    NOR2X1 U619 (.A1(N1237), .A2(N1238), .ZN(n13491));
    NANDX1 U620 (.A1(N1239), .A2(N1240), .ZN(N13492));
    NANDX1 U621 (.A1(N1241), .A2(N1242), .ZN(n13493));
    NANDX1 U622 (.A1(N1243), .A2(N1244), .ZN(n13494));
    NANDX1 U623 (.A1(N1245), .A2(N1246), .ZN(n13495));
    NANDX1 U624 (.A1(N1247), .A2(N1248), .ZN(n13496));
    NANDX1 U625 (.A1(N1249), .A2(N1250), .ZN(n13497));
    NOR2X1 U626 (.A1(N1251), .A2(N1252), .ZN(n13498));
    NOR2X1 U627 (.A1(N1253), .A2(N1254), .ZN(n13499));
    NOR2X1 U628 (.A1(N1255), .A2(N1256), .ZN(n13500));
    NOR2X1 U629 (.A1(N1257), .A2(N1258), .ZN(n13501));
    NANDX1 U630 (.A1(N1259), .A2(N1260), .ZN(n13502));
    NANDX1 U631 (.A1(N1261), .A2(N1262), .ZN(n13503));
    NOR2X1 U632 (.A1(N1263), .A2(N1264), .ZN(n13504));
    NOR2X1 U633 (.A1(N1265), .A2(N1266), .ZN(N13505));
    NOR2X1 U634 (.A1(N1267), .A2(N1268), .ZN(n13506));
    NANDX1 U635 (.A1(N1269), .A2(N1270), .ZN(n13507));
    NANDX1 U636 (.A1(N1271), .A2(N1272), .ZN(n13508));
    NOR2X1 U637 (.A1(N1273), .A2(N1274), .ZN(n13509));
    NOR2X1 U638 (.A1(N1275), .A2(N1276), .ZN(n13510));
    NOR2X1 U639 (.A1(N1277), .A2(N1278), .ZN(n13511));
    NOR2X1 U640 (.A1(N1279), .A2(N1280), .ZN(N13512));
    NOR2X1 U641 (.A1(N1281), .A2(N1282), .ZN(n13513));
    NANDX1 U642 (.A1(N1283), .A2(N1284), .ZN(N13514));
    NOR2X1 U643 (.A1(N1285), .A2(N1286), .ZN(n13515));
    NOR2X1 U644 (.A1(N1287), .A2(N1288), .ZN(n13516));
    NOR2X1 U645 (.A1(N1289), .A2(N1290), .ZN(N13517));
    NANDX1 U646 (.A1(N1291), .A2(N1292), .ZN(n13518));
    NANDX1 U647 (.A1(N1293), .A2(N1294), .ZN(n13519));
    NANDX1 U648 (.A1(N1295), .A2(N1296), .ZN(n13520));
    NOR2X1 U649 (.A1(N1297), .A2(N1298), .ZN(n13521));
    NOR2X1 U650 (.A1(N1299), .A2(N1300), .ZN(n13522));
    NOR2X1 U651 (.A1(N1301), .A2(N1302), .ZN(n13523));
    NANDX1 U652 (.A1(N1303), .A2(N1304), .ZN(N13524));
    NANDX1 U653 (.A1(N1305), .A2(N1306), .ZN(n13525));
    NANDX1 U654 (.A1(N1307), .A2(N1308), .ZN(n13526));
    NANDX1 U655 (.A1(N1309), .A2(N1310), .ZN(N13527));
    NOR2X1 U656 (.A1(N1311), .A2(N1312), .ZN(n13528));
    NANDX1 U657 (.A1(N1313), .A2(N1314), .ZN(n13529));
    NANDX1 U658 (.A1(N1315), .A2(N1316), .ZN(n13530));
    NANDX1 U659 (.A1(N1317), .A2(N1318), .ZN(n13531));
    NOR2X1 U660 (.A1(N1319), .A2(N1320), .ZN(n13532));
    NOR2X1 U661 (.A1(N1321), .A2(N1322), .ZN(N13533));
    NOR2X1 U662 (.A1(N1323), .A2(N1324), .ZN(n13534));
    NOR2X1 U663 (.A1(N1325), .A2(N1326), .ZN(n13535));
    NANDX1 U664 (.A1(N1327), .A2(N1328), .ZN(N13536));
    NANDX1 U665 (.A1(N1329), .A2(N1330), .ZN(n13537));
    NANDX1 U666 (.A1(N1331), .A2(N1332), .ZN(n13538));
    NOR2X1 U667 (.A1(N1333), .A2(N1334), .ZN(n13539));
    NANDX1 U668 (.A1(N1335), .A2(N1336), .ZN(n13540));
    NANDX1 U669 (.A1(N1337), .A2(N1338), .ZN(n13541));
    NOR2X1 U670 (.A1(N1339), .A2(N1340), .ZN(n13542));
    NANDX1 U671 (.A1(N1341), .A2(N1342), .ZN(n13543));
    NANDX1 U672 (.A1(N1343), .A2(N1344), .ZN(n13544));
    NANDX1 U673 (.A1(N1345), .A2(N1346), .ZN(n13545));
    NOR2X1 U674 (.A1(N1347), .A2(N1348), .ZN(n13546));
    NANDX1 U675 (.A1(N1349), .A2(N1350), .ZN(N13547));
    NOR2X1 U676 (.A1(N1351), .A2(N1352), .ZN(N13548));
    NANDX1 U677 (.A1(N1353), .A2(N1354), .ZN(n13549));
    NOR2X1 U678 (.A1(N1355), .A2(N1356), .ZN(n13550));
    NANDX1 U679 (.A1(N1357), .A2(N1358), .ZN(N13551));
    NOR2X1 U680 (.A1(N1359), .A2(N1360), .ZN(n13552));
    NOR2X1 U681 (.A1(N1361), .A2(N1362), .ZN(n13553));
    NOR2X1 U682 (.A1(N1363), .A2(N1364), .ZN(n13554));
    NANDX1 U683 (.A1(N1365), .A2(N1366), .ZN(n13555));
    NOR2X1 U684 (.A1(N1367), .A2(N1368), .ZN(N13556));
    NANDX1 U685 (.A1(N1369), .A2(N1370), .ZN(n13557));
    NOR2X1 U686 (.A1(N1371), .A2(N1372), .ZN(n13558));
    NOR2X1 U687 (.A1(N1373), .A2(N1374), .ZN(n13559));
    NANDX1 U688 (.A1(N1375), .A2(N1376), .ZN(n13560));
    NOR2X1 U689 (.A1(N1377), .A2(N1378), .ZN(n13561));
    NANDX1 U690 (.A1(N1379), .A2(N1380), .ZN(n13562));
    NANDX1 U691 (.A1(N1381), .A2(N1382), .ZN(N13563));
    NOR2X1 U692 (.A1(N1383), .A2(N1384), .ZN(n13564));
    NOR2X1 U693 (.A1(N1385), .A2(N1386), .ZN(n13565));
    NANDX1 U694 (.A1(N1387), .A2(N1388), .ZN(N13566));
    NANDX1 U695 (.A1(N1389), .A2(N1390), .ZN(n13567));
    NANDX1 U696 (.A1(N1391), .A2(N1392), .ZN(n13568));
    NOR2X1 U697 (.A1(N1393), .A2(N1394), .ZN(n13569));
    NANDX1 U698 (.A1(N1395), .A2(N1396), .ZN(n13570));
    NOR2X1 U699 (.A1(N1397), .A2(N1398), .ZN(n13571));
    NANDX1 U700 (.A1(N1399), .A2(N1400), .ZN(n13572));
    NOR2X1 U701 (.A1(N1401), .A2(N1402), .ZN(n13573));
    NOR2X1 U702 (.A1(N1403), .A2(N1404), .ZN(n13574));
    NOR2X1 U703 (.A1(N1405), .A2(N1406), .ZN(n13575));
    NANDX1 U704 (.A1(N1407), .A2(N1408), .ZN(n13576));
    NOR2X1 U705 (.A1(N1409), .A2(N1410), .ZN(N13577));
    NANDX1 U706 (.A1(N1411), .A2(N1412), .ZN(n13578));
    NANDX1 U707 (.A1(N1413), .A2(N1414), .ZN(n13579));
    NANDX1 U708 (.A1(N1415), .A2(N1416), .ZN(n13580));
    NANDX1 U709 (.A1(N1417), .A2(N1418), .ZN(n13581));
    NANDX1 U710 (.A1(N1419), .A2(N1420), .ZN(n13582));
    NANDX1 U711 (.A1(N1421), .A2(N1422), .ZN(n13583));
    NOR2X1 U712 (.A1(N1423), .A2(N1424), .ZN(n13584));
    NANDX1 U713 (.A1(N1425), .A2(N1426), .ZN(n13585));
    NANDX1 U714 (.A1(N1427), .A2(N1428), .ZN(n13586));
    NOR2X1 U715 (.A1(N1429), .A2(N1430), .ZN(n13587));
    NOR2X1 U716 (.A1(N1431), .A2(N1432), .ZN(n13588));
    NANDX1 U717 (.A1(N1433), .A2(N1434), .ZN(N13589));
    NOR2X1 U718 (.A1(N1435), .A2(N1436), .ZN(n13590));
    NANDX1 U719 (.A1(N1437), .A2(N1438), .ZN(n13591));
    NANDX1 U720 (.A1(N1439), .A2(N1440), .ZN(n13592));
    NOR2X1 U721 (.A1(N1441), .A2(N1442), .ZN(n13593));
    NOR2X1 U722 (.A1(N1443), .A2(N1444), .ZN(N13594));
    NOR2X1 U723 (.A1(N1445), .A2(N1446), .ZN(N13595));
    NOR2X1 U724 (.A1(N1447), .A2(N1448), .ZN(n13596));
    NANDX1 U725 (.A1(N1449), .A2(N1450), .ZN(n13597));
    NANDX1 U726 (.A1(N1451), .A2(N1452), .ZN(n13598));
    NANDX1 U727 (.A1(N1453), .A2(N1454), .ZN(n13599));
    NANDX1 U728 (.A1(N1455), .A2(N1456), .ZN(n13600));
    NANDX1 U729 (.A1(N1457), .A2(N1458), .ZN(n13601));
    NANDX1 U730 (.A1(N1459), .A2(N1460), .ZN(n13602));
    NOR2X1 U731 (.A1(N1461), .A2(N1462), .ZN(n13603));
    NANDX1 U732 (.A1(N1463), .A2(N1464), .ZN(n13604));
    NANDX1 U733 (.A1(N1465), .A2(N1466), .ZN(n13605));
    NOR2X1 U734 (.A1(N1467), .A2(N1468), .ZN(n13606));
    NOR2X1 U735 (.A1(N1469), .A2(N1470), .ZN(n13607));
    NANDX1 U736 (.A1(N1471), .A2(N1472), .ZN(N13608));
    NANDX1 U737 (.A1(N1473), .A2(N1474), .ZN(n13609));
    NOR2X1 U738 (.A1(N1475), .A2(N1476), .ZN(N13610));
    NANDX1 U739 (.A1(N1477), .A2(N1478), .ZN(N13611));
    NANDX1 U740 (.A1(N1479), .A2(N1480), .ZN(N13612));
    NANDX1 U741 (.A1(N1481), .A2(N1482), .ZN(n13613));
    NOR2X1 U742 (.A1(N1483), .A2(N1484), .ZN(n13614));
    NANDX1 U743 (.A1(N1485), .A2(N1486), .ZN(N13615));
    NOR2X1 U744 (.A1(N1487), .A2(N1488), .ZN(N13616));
    NANDX1 U745 (.A1(N1489), .A2(N1490), .ZN(n13617));
    NANDX1 U746 (.A1(N1491), .A2(N1492), .ZN(n13618));
    NOR2X1 U747 (.A1(N1493), .A2(N1494), .ZN(n13619));
    NANDX1 U748 (.A1(N1495), .A2(N1496), .ZN(n13620));
    NANDX1 U749 (.A1(N1497), .A2(N1498), .ZN(n13621));
    NOR2X1 U750 (.A1(N1499), .A2(N1500), .ZN(n13622));
    NOR2X1 U751 (.A1(N1501), .A2(N1502), .ZN(n13623));
    NANDX1 U752 (.A1(N1503), .A2(N1504), .ZN(n13624));
    NOR2X1 U753 (.A1(N1505), .A2(N1506), .ZN(n13625));
    NOR2X1 U754 (.A1(N1507), .A2(N1508), .ZN(n13626));
    NANDX1 U755 (.A1(N1509), .A2(N1510), .ZN(n13627));
    NOR2X1 U756 (.A1(N1511), .A2(N1512), .ZN(N13628));
    NOR2X1 U757 (.A1(N1513), .A2(N1514), .ZN(n13629));
    NOR2X1 U758 (.A1(N1515), .A2(N1516), .ZN(n13630));
    NANDX1 U759 (.A1(N1517), .A2(N1518), .ZN(n13631));
    NANDX1 U760 (.A1(N1519), .A2(N1520), .ZN(n13632));
    NOR2X1 U761 (.A1(N1521), .A2(N1522), .ZN(N13633));
    NOR2X1 U762 (.A1(N1523), .A2(N1524), .ZN(n13634));
    NOR2X1 U763 (.A1(N1525), .A2(N1526), .ZN(n13635));
    NANDX1 U764 (.A1(N1527), .A2(N1528), .ZN(n13636));
    NOR2X1 U765 (.A1(N1529), .A2(N1530), .ZN(n13637));
    NOR2X1 U766 (.A1(N1531), .A2(N1532), .ZN(n13638));
    NANDX1 U767 (.A1(N1533), .A2(N1534), .ZN(n13639));
    NOR2X1 U768 (.A1(N1535), .A2(N1536), .ZN(n13640));
    NOR2X1 U769 (.A1(N1537), .A2(N1538), .ZN(n13641));
    NOR2X1 U770 (.A1(N1539), .A2(N1540), .ZN(n13642));
    NANDX1 U771 (.A1(N1541), .A2(N1542), .ZN(n13643));
    NANDX1 U772 (.A1(N1543), .A2(N1544), .ZN(n13644));
    NOR2X1 U773 (.A1(N1545), .A2(N1546), .ZN(n13645));
    NOR2X1 U774 (.A1(N1547), .A2(N1548), .ZN(n13646));
    NANDX1 U775 (.A1(N1549), .A2(N1550), .ZN(N13647));
    NOR2X1 U776 (.A1(N1551), .A2(N1552), .ZN(n13648));
    NANDX1 U777 (.A1(N1553), .A2(N1554), .ZN(n13649));
    NOR2X1 U778 (.A1(N1555), .A2(N1556), .ZN(N13650));
    NANDX1 U779 (.A1(N1557), .A2(N1558), .ZN(N13651));
    NOR2X1 U780 (.A1(N1559), .A2(N1560), .ZN(n13652));
    NOR2X1 U781 (.A1(N1561), .A2(N1562), .ZN(n13653));
    NANDX1 U782 (.A1(N1563), .A2(N1564), .ZN(n13654));
    NOR2X1 U783 (.A1(N1565), .A2(N1566), .ZN(n13655));
    NOR2X1 U784 (.A1(N1567), .A2(N1568), .ZN(n13656));
    NOR2X1 U785 (.A1(N1569), .A2(N1570), .ZN(n13657));
    NANDX1 U786 (.A1(N1571), .A2(N1572), .ZN(n13658));
    NOR2X1 U787 (.A1(N1573), .A2(N1574), .ZN(n13659));
    NOR2X1 U788 (.A1(N1575), .A2(N1576), .ZN(n13660));
    NOR2X1 U789 (.A1(N1577), .A2(N1578), .ZN(n13661));
    NOR2X1 U790 (.A1(N1579), .A2(N1580), .ZN(n13662));
    NANDX1 U791 (.A1(N1581), .A2(N1582), .ZN(N13663));
    NOR2X1 U792 (.A1(N1583), .A2(N1584), .ZN(n13664));
    NOR2X1 U793 (.A1(N1585), .A2(N1586), .ZN(n13665));
    NANDX1 U794 (.A1(N1587), .A2(N1588), .ZN(N13666));
    NANDX1 U795 (.A1(N1589), .A2(N1590), .ZN(n13667));
    NOR2X1 U796 (.A1(N1591), .A2(N1592), .ZN(n13668));
    NANDX1 U797 (.A1(N1593), .A2(N1594), .ZN(n13669));
    NOR2X1 U798 (.A1(N1595), .A2(N1596), .ZN(n13670));
    NOR2X1 U799 (.A1(N1597), .A2(N1598), .ZN(n13671));
    NOR2X1 U800 (.A1(N1599), .A2(N1600), .ZN(n13672));
    NOR2X1 U801 (.A1(N1601), .A2(N1602), .ZN(N13673));
    NANDX1 U802 (.A1(N1603), .A2(N1604), .ZN(N13674));
    NANDX1 U803 (.A1(N1605), .A2(N1606), .ZN(n13675));
    NANDX1 U804 (.A1(N1607), .A2(N1608), .ZN(n13676));
    NANDX1 U805 (.A1(N1609), .A2(N1610), .ZN(n13677));
    NANDX1 U806 (.A1(N1611), .A2(N1612), .ZN(n13678));
    NANDX1 U807 (.A1(N1613), .A2(N1614), .ZN(N13679));
    NOR2X1 U808 (.A1(N1615), .A2(N1616), .ZN(n13680));
    NANDX1 U809 (.A1(N1617), .A2(N1618), .ZN(N13681));
    NOR2X1 U810 (.A1(N1619), .A2(N1620), .ZN(n13682));
    NANDX1 U811 (.A1(N1621), .A2(N1622), .ZN(n13683));
    NANDX1 U812 (.A1(N1623), .A2(N1624), .ZN(N13684));
    NANDX1 U813 (.A1(N1625), .A2(N1626), .ZN(n13685));
    NANDX1 U814 (.A1(N1627), .A2(N1628), .ZN(N13686));
    NANDX1 U815 (.A1(N1629), .A2(N1630), .ZN(n13687));
    NANDX1 U816 (.A1(N1631), .A2(N1632), .ZN(n13688));
    NOR2X1 U817 (.A1(N1633), .A2(N1634), .ZN(n13689));
    NOR2X1 U818 (.A1(N1635), .A2(N1636), .ZN(n13690));
    NANDX1 U819 (.A1(N1637), .A2(N1638), .ZN(N13691));
    NOR2X1 U820 (.A1(N1639), .A2(N1640), .ZN(n13692));
    NOR2X1 U821 (.A1(N1641), .A2(N1642), .ZN(n13693));
    NOR2X1 U822 (.A1(N1643), .A2(N1644), .ZN(n13694));
    NOR2X1 U823 (.A1(N1645), .A2(N1646), .ZN(n13695));
    NOR2X1 U824 (.A1(N1647), .A2(N1648), .ZN(n13696));
    NANDX1 U825 (.A1(N1649), .A2(N1650), .ZN(n13697));
    NOR2X1 U826 (.A1(N1651), .A2(N1652), .ZN(n13698));
    NOR2X1 U827 (.A1(N1653), .A2(N1654), .ZN(N13699));
    NANDX1 U828 (.A1(N1655), .A2(N1656), .ZN(N13700));
    NOR2X1 U829 (.A1(N1657), .A2(N1658), .ZN(n13701));
    NANDX1 U830 (.A1(N1659), .A2(N1660), .ZN(n13702));
    NANDX1 U831 (.A1(N1661), .A2(N1662), .ZN(n13703));
    NANDX1 U832 (.A1(N1663), .A2(N1664), .ZN(n13704));
    NOR2X1 U833 (.A1(N1665), .A2(N1666), .ZN(n13705));
    NOR2X1 U834 (.A1(N1667), .A2(N1668), .ZN(n13706));
    NOR2X1 U835 (.A1(N1669), .A2(N1670), .ZN(N13707));
    NOR2X1 U836 (.A1(N1671), .A2(N1672), .ZN(n13708));
    NANDX1 U837 (.A1(N1673), .A2(N1674), .ZN(n13709));
    NANDX1 U838 (.A1(N1675), .A2(N1676), .ZN(n13710));
    NOR2X1 U839 (.A1(N1677), .A2(N1678), .ZN(N13711));
    NOR2X1 U840 (.A1(N1679), .A2(N1680), .ZN(n13712));
    NANDX1 U841 (.A1(N1681), .A2(N1682), .ZN(n13713));
    NANDX1 U842 (.A1(N1683), .A2(N1684), .ZN(n13714));
    NANDX1 U843 (.A1(N1685), .A2(N1686), .ZN(n13715));
    NOR2X1 U844 (.A1(N1687), .A2(N1688), .ZN(n13716));
    NOR2X1 U845 (.A1(N1689), .A2(N1690), .ZN(n13717));
    NANDX1 U846 (.A1(N1691), .A2(N1692), .ZN(N13718));
    NOR2X1 U847 (.A1(N1693), .A2(N1694), .ZN(N13719));
    NANDX1 U848 (.A1(N1695), .A2(N1696), .ZN(n13720));
    NANDX1 U849 (.A1(N1697), .A2(N1698), .ZN(n13721));
    NANDX1 U850 (.A1(N1699), .A2(N1700), .ZN(n13722));
    NANDX1 U851 (.A1(N1701), .A2(N1702), .ZN(n13723));
    NANDX1 U852 (.A1(N1703), .A2(N1704), .ZN(n13724));
    NOR2X1 U853 (.A1(N1705), .A2(N1706), .ZN(n13725));
    NOR2X1 U854 (.A1(N1707), .A2(N1708), .ZN(n13726));
    NANDX1 U855 (.A1(N1709), .A2(N1710), .ZN(n13727));
    NANDX1 U856 (.A1(N1711), .A2(N1712), .ZN(n13728));
    NOR2X1 U857 (.A1(N1713), .A2(N1714), .ZN(n13729));
    NANDX1 U858 (.A1(N1715), .A2(N1716), .ZN(n13730));
    NOR2X1 U859 (.A1(N1717), .A2(N1718), .ZN(n13731));
    NOR2X1 U860 (.A1(N1719), .A2(N1720), .ZN(n13732));
    NOR2X1 U861 (.A1(N1721), .A2(N1722), .ZN(n13733));
    NANDX1 U862 (.A1(N1723), .A2(N1724), .ZN(N13734));
    NANDX1 U863 (.A1(N1725), .A2(N1726), .ZN(n13735));
    NANDX1 U864 (.A1(N1727), .A2(N1728), .ZN(n13736));
    NOR2X1 U865 (.A1(N1729), .A2(N1730), .ZN(N13737));
    NANDX1 U866 (.A1(N1731), .A2(N1732), .ZN(n13738));
    NANDX1 U867 (.A1(N1733), .A2(N1734), .ZN(n13739));
    NANDX1 U868 (.A1(N1735), .A2(N1736), .ZN(n13740));
    NOR2X1 U869 (.A1(N1737), .A2(N1738), .ZN(N13741));
    NANDX1 U870 (.A1(N1739), .A2(N1740), .ZN(N13742));
    NOR2X1 U871 (.A1(N1741), .A2(N1742), .ZN(n13743));
    NANDX1 U872 (.A1(N1743), .A2(N1744), .ZN(n13744));
    NANDX1 U873 (.A1(N1745), .A2(N1746), .ZN(n13745));
    NANDX1 U874 (.A1(N1747), .A2(N1748), .ZN(n13746));
    NOR2X1 U875 (.A1(N1749), .A2(N1750), .ZN(n13747));
    NANDX1 U876 (.A1(N1751), .A2(N1752), .ZN(n13748));
    NOR2X1 U877 (.A1(N1753), .A2(N1754), .ZN(n13749));
    NOR2X1 U878 (.A1(N1755), .A2(N1756), .ZN(n13750));
    NOR2X1 U879 (.A1(N1757), .A2(N1758), .ZN(n13751));
    NANDX1 U880 (.A1(N1759), .A2(N1760), .ZN(n13752));
    NANDX1 U881 (.A1(N1761), .A2(N1762), .ZN(n13753));
    NOR2X1 U882 (.A1(N1763), .A2(N1764), .ZN(n13754));
    NOR2X1 U883 (.A1(N1765), .A2(N1766), .ZN(n13755));
    NANDX1 U884 (.A1(N1767), .A2(N1768), .ZN(n13756));
    NOR2X1 U885 (.A1(N1769), .A2(N1770), .ZN(n13757));
    NANDX1 U886 (.A1(N1771), .A2(N1772), .ZN(n13758));
    NANDX1 U887 (.A1(N1773), .A2(N1774), .ZN(n13759));
    NOR2X1 U888 (.A1(N1775), .A2(N1776), .ZN(n13760));
    NANDX1 U889 (.A1(N1777), .A2(N1778), .ZN(N13761));
    NANDX1 U890 (.A1(N1779), .A2(N1780), .ZN(n13762));
    NOR2X1 U891 (.A1(N1781), .A2(N1782), .ZN(n13763));
    NANDX1 U892 (.A1(N1783), .A2(N1784), .ZN(n13764));
    NANDX1 U893 (.A1(N1785), .A2(N1786), .ZN(n13765));
    NOR2X1 U894 (.A1(N1787), .A2(N1788), .ZN(n13766));
    NOR2X1 U895 (.A1(N1789), .A2(N1790), .ZN(N13767));
    NANDX1 U896 (.A1(N1791), .A2(N1792), .ZN(n13768));
    NANDX1 U897 (.A1(N1793), .A2(N1794), .ZN(n13769));
    NANDX1 U898 (.A1(N1795), .A2(N1796), .ZN(N13770));
    NOR2X1 U899 (.A1(N1797), .A2(N1798), .ZN(n13771));
    NOR2X1 U900 (.A1(N1799), .A2(N1800), .ZN(n13772));
    NANDX1 U901 (.A1(N1801), .A2(N1802), .ZN(n13773));
    NOR2X1 U902 (.A1(N1803), .A2(N1804), .ZN(n13774));
    NANDX1 U903 (.A1(N1805), .A2(N1806), .ZN(N13775));
    NOR2X1 U904 (.A1(N1807), .A2(N1808), .ZN(N13776));
    NOR2X1 U905 (.A1(N1809), .A2(N1810), .ZN(n13777));
    NANDX1 U906 (.A1(N1811), .A2(N1812), .ZN(n13778));
    NANDX1 U907 (.A1(N1813), .A2(N1814), .ZN(n13779));
    NOR2X1 U908 (.A1(N1815), .A2(N1816), .ZN(n13780));
    NANDX1 U909 (.A1(N1817), .A2(N1818), .ZN(N13781));
    NOR2X1 U910 (.A1(N1819), .A2(N1820), .ZN(n13782));
    NOR2X1 U911 (.A1(N1821), .A2(N1822), .ZN(n13783));
    NANDX1 U912 (.A1(N1823), .A2(N1824), .ZN(n13784));
    NOR2X1 U913 (.A1(N1825), .A2(N1826), .ZN(N13785));
    NOR2X1 U914 (.A1(N1827), .A2(N1828), .ZN(n13786));
    NOR2X1 U915 (.A1(N1829), .A2(N1830), .ZN(n13787));
    NOR2X1 U916 (.A1(N1831), .A2(N1832), .ZN(n13788));
    NOR2X1 U917 (.A1(N1833), .A2(N1834), .ZN(N13789));
    NANDX1 U918 (.A1(N1835), .A2(N1836), .ZN(n13790));
    NOR2X1 U919 (.A1(N1837), .A2(N1838), .ZN(n13791));
    NANDX1 U920 (.A1(N1839), .A2(N1840), .ZN(n13792));
    NANDX1 U921 (.A1(N1841), .A2(N1842), .ZN(n13793));
    NOR2X1 U922 (.A1(N1843), .A2(N1844), .ZN(n13794));
    NOR2X1 U923 (.A1(N1845), .A2(N1846), .ZN(n13795));
    NOR2X1 U924 (.A1(N1847), .A2(N1848), .ZN(n13796));
    NOR2X1 U925 (.A1(N1849), .A2(N1850), .ZN(n13797));
    NANDX1 U926 (.A1(N1851), .A2(N1852), .ZN(n13798));
    NANDX1 U927 (.A1(N1853), .A2(N1854), .ZN(n13799));
    NOR2X1 U928 (.A1(N1855), .A2(N1856), .ZN(n13800));
    NOR2X1 U929 (.A1(N1857), .A2(N1858), .ZN(n13801));
    NANDX1 U930 (.A1(N1859), .A2(N1860), .ZN(n13802));
    NOR2X1 U931 (.A1(N1861), .A2(N1862), .ZN(N13803));
    NANDX1 U932 (.A1(N1863), .A2(N1864), .ZN(n13804));
    NOR2X1 U933 (.A1(N1865), .A2(N1866), .ZN(n13805));
    NANDX1 U934 (.A1(N1867), .A2(N1868), .ZN(N13806));
    NANDX1 U935 (.A1(N1869), .A2(N1870), .ZN(n13807));
    NOR2X1 U936 (.A1(N1871), .A2(N1872), .ZN(n13808));
    NANDX1 U937 (.A1(N1873), .A2(N1874), .ZN(N13809));
    NANDX1 U938 (.A1(N1875), .A2(N1876), .ZN(n13810));
    NOR2X1 U939 (.A1(N1877), .A2(N1878), .ZN(N13811));
    NOR2X1 U940 (.A1(N1879), .A2(N1880), .ZN(n13812));
    NANDX1 U941 (.A1(N1881), .A2(N1882), .ZN(n13813));
    NOR2X1 U942 (.A1(N1883), .A2(N1884), .ZN(n13814));
    NANDX1 U943 (.A1(N1885), .A2(N1886), .ZN(n13815));
    NANDX1 U944 (.A1(N1887), .A2(N1888), .ZN(n13816));
    NANDX1 U945 (.A1(N1889), .A2(N1890), .ZN(n13817));
    NOR2X1 U946 (.A1(N1891), .A2(N1892), .ZN(n13818));
    NANDX1 U947 (.A1(N1893), .A2(N1894), .ZN(N13819));
    NANDX1 U948 (.A1(N1895), .A2(N1896), .ZN(N13820));
    NANDX1 U949 (.A1(N1897), .A2(N1898), .ZN(n13821));
    NANDX1 U950 (.A1(N1899), .A2(N1900), .ZN(n13822));
    NOR2X1 U951 (.A1(N1901), .A2(N1902), .ZN(n13823));
    NOR2X1 U952 (.A1(N1903), .A2(N1904), .ZN(n13824));
    NANDX1 U953 (.A1(N1905), .A2(N1906), .ZN(n13825));
    NOR2X1 U954 (.A1(N1907), .A2(N1908), .ZN(n13826));
    NOR2X1 U955 (.A1(N1909), .A2(N1910), .ZN(n13827));
    NOR2X1 U956 (.A1(N1911), .A2(N1912), .ZN(N13828));
    NANDX1 U957 (.A1(N1913), .A2(N1914), .ZN(n13829));
    NANDX1 U958 (.A1(N1915), .A2(N1916), .ZN(n13830));
    NOR2X1 U959 (.A1(N1917), .A2(N1918), .ZN(n13831));
    NOR2X1 U960 (.A1(N1919), .A2(N1920), .ZN(n13832));
    NANDX1 U961 (.A1(N1921), .A2(N1922), .ZN(n13833));
    NOR2X1 U962 (.A1(N1923), .A2(N1924), .ZN(n13834));
    NANDX1 U963 (.A1(N1925), .A2(N1926), .ZN(n13835));
    NANDX1 U964 (.A1(N1927), .A2(N1928), .ZN(n13836));
    NANDX1 U965 (.A1(N1929), .A2(N1930), .ZN(n13837));
    NANDX1 U966 (.A1(N1931), .A2(N1932), .ZN(N13838));
    NANDX1 U967 (.A1(N1933), .A2(N1934), .ZN(n13839));
    NOR2X1 U968 (.A1(N1935), .A2(N1936), .ZN(n13840));
    NOR2X1 U969 (.A1(N1937), .A2(N1938), .ZN(n13841));
    NANDX1 U970 (.A1(N1939), .A2(N1940), .ZN(N13842));
    NANDX1 U971 (.A1(N1941), .A2(N1942), .ZN(n13843));
    NANDX1 U972 (.A1(N1943), .A2(N1944), .ZN(N13844));
    NOR2X1 U973 (.A1(N1945), .A2(N1946), .ZN(n13845));
    NOR2X1 U974 (.A1(N1947), .A2(N1948), .ZN(n13846));
    NOR2X1 U975 (.A1(N1949), .A2(N1950), .ZN(N13847));
    NANDX1 U976 (.A1(N1951), .A2(N1952), .ZN(n13848));
    NOR2X1 U977 (.A1(N1953), .A2(N1954), .ZN(n13849));
    NANDX1 U978 (.A1(N1955), .A2(N1956), .ZN(n13850));
    NOR2X1 U979 (.A1(N1957), .A2(N1958), .ZN(n13851));
    NOR2X1 U980 (.A1(N1959), .A2(N1960), .ZN(N13852));
    NOR2X1 U981 (.A1(N1961), .A2(N1962), .ZN(n13853));
    NOR2X1 U982 (.A1(N1963), .A2(N1964), .ZN(n13854));
    NOR2X1 U983 (.A1(N1965), .A2(N1966), .ZN(n13855));
    NANDX1 U984 (.A1(N1967), .A2(N1968), .ZN(n13856));
    NOR2X1 U985 (.A1(N1969), .A2(N1970), .ZN(n13857));
    NANDX1 U986 (.A1(N1971), .A2(N1972), .ZN(N13858));
    NANDX1 U987 (.A1(N1973), .A2(N1974), .ZN(n13859));
    NOR2X1 U988 (.A1(N1975), .A2(N1976), .ZN(n13860));
    NOR2X1 U989 (.A1(N1977), .A2(N1978), .ZN(n13861));
    NANDX1 U990 (.A1(N1979), .A2(N1980), .ZN(n13862));
    NOR2X1 U991 (.A1(N1981), .A2(N1982), .ZN(n13863));
    NANDX1 U992 (.A1(N1983), .A2(N1984), .ZN(n13864));
    NANDX1 U993 (.A1(N1985), .A2(N1986), .ZN(n13865));
    NANDX1 U994 (.A1(N1987), .A2(N1988), .ZN(n13866));
    NOR2X1 U995 (.A1(N1989), .A2(N1990), .ZN(N13867));
    NANDX1 U996 (.A1(N1991), .A2(N1992), .ZN(n13868));
    NOR2X1 U997 (.A1(N1993), .A2(N1994), .ZN(N13869));
    NANDX1 U998 (.A1(N1995), .A2(N1996), .ZN(N13870));
    NANDX1 U999 (.A1(N1997), .A2(N1998), .ZN(n13871));
    NOR2X1 U1000 (.A1(N1999), .A2(N2000), .ZN(n13872));
    NANDX1 U1001 (.A1(N2001), .A2(N2002), .ZN(N13873));
    NOR2X1 U1002 (.A1(N2003), .A2(N2004), .ZN(n13874));
    NANDX1 U1003 (.A1(N2005), .A2(N2006), .ZN(n13875));
    NANDX1 U1004 (.A1(N2007), .A2(N2008), .ZN(n13876));
    NANDX1 U1005 (.A1(N2009), .A2(N2010), .ZN(n13877));
    NANDX1 U1006 (.A1(N2011), .A2(N2012), .ZN(n13878));
    NOR2X1 U1007 (.A1(N2013), .A2(N2014), .ZN(n13879));
    NANDX1 U1008 (.A1(N2015), .A2(N2016), .ZN(N13880));
    NOR2X1 U1009 (.A1(N2017), .A2(N2018), .ZN(n13881));
    NOR2X1 U1010 (.A1(N2019), .A2(N2020), .ZN(n13882));
    NANDX1 U1011 (.A1(N2021), .A2(N2022), .ZN(n13883));
    NOR2X1 U1012 (.A1(N2023), .A2(N2024), .ZN(n13884));
    NOR2X1 U1013 (.A1(N2025), .A2(N2026), .ZN(N13885));
    NOR2X1 U1014 (.A1(N2027), .A2(N2028), .ZN(n13886));
    NOR2X1 U1015 (.A1(N2029), .A2(N2030), .ZN(n13887));
    NOR2X1 U1016 (.A1(N2031), .A2(N2032), .ZN(n13888));
    NANDX1 U1017 (.A1(N2033), .A2(N2034), .ZN(n13889));
    NANDX1 U1018 (.A1(N2035), .A2(N2036), .ZN(n13890));
    NOR2X1 U1019 (.A1(N2037), .A2(N2038), .ZN(n13891));
    NANDX1 U1020 (.A1(N2039), .A2(N2040), .ZN(n13892));
    NANDX1 U1021 (.A1(N2041), .A2(N2042), .ZN(N13893));
    NOR2X1 U1022 (.A1(N2043), .A2(N2044), .ZN(n13894));
    NANDX1 U1023 (.A1(N2045), .A2(N2046), .ZN(n13895));
    NOR2X1 U1024 (.A1(N2047), .A2(N2048), .ZN(N13896));
    NOR2X1 U1025 (.A1(N2049), .A2(N2050), .ZN(n13897));
    NANDX1 U1026 (.A1(N2051), .A2(N2052), .ZN(n13898));
    NANDX1 U1027 (.A1(N2053), .A2(N2054), .ZN(n13899));
    NOR2X1 U1028 (.A1(N2055), .A2(N2056), .ZN(n13900));
    NANDX1 U1029 (.A1(N2057), .A2(N2058), .ZN(N13901));
    NANDX1 U1030 (.A1(N2059), .A2(N2060), .ZN(n13902));
    NANDX1 U1031 (.A1(N2061), .A2(N2062), .ZN(n13903));
    NOR2X1 U1032 (.A1(N2063), .A2(N2064), .ZN(n13904));
    NANDX1 U1033 (.A1(N2065), .A2(N2066), .ZN(N13905));
    NOR2X1 U1034 (.A1(N2067), .A2(N2068), .ZN(N13906));
    NANDX1 U1035 (.A1(N2069), .A2(N2070), .ZN(n13907));
    NOR2X1 U1036 (.A1(N2071), .A2(N2072), .ZN(n13908));
    NOR2X1 U1037 (.A1(N2073), .A2(N2074), .ZN(n13909));
    NANDX1 U1038 (.A1(N2075), .A2(N2076), .ZN(N13910));
    NOR2X1 U1039 (.A1(N2077), .A2(N2078), .ZN(n13911));
    NOR2X1 U1040 (.A1(N2079), .A2(N2080), .ZN(n13912));
    NANDX1 U1041 (.A1(N2081), .A2(N2082), .ZN(n13913));
    NANDX1 U1042 (.A1(N2083), .A2(N2084), .ZN(n13914));
    NANDX1 U1043 (.A1(N2085), .A2(N2086), .ZN(N13915));
    NANDX1 U1044 (.A1(N2087), .A2(N2088), .ZN(n13916));
    NANDX1 U1045 (.A1(N2089), .A2(N2090), .ZN(n13917));
    NANDX1 U1046 (.A1(N2091), .A2(N2092), .ZN(n13918));
    NANDX1 U1047 (.A1(N2093), .A2(N2094), .ZN(n13919));
    NOR2X1 U1048 (.A1(N2095), .A2(N2096), .ZN(N13920));
    NOR2X1 U1049 (.A1(N2097), .A2(N2098), .ZN(N13921));
    NOR2X1 U1050 (.A1(N2099), .A2(N2100), .ZN(n13922));
    NOR2X1 U1051 (.A1(N2101), .A2(N2102), .ZN(n13923));
    NANDX1 U1052 (.A1(N2103), .A2(N2104), .ZN(n13924));
    NOR2X1 U1053 (.A1(N2105), .A2(N2106), .ZN(n13925));
    NANDX1 U1054 (.A1(N2107), .A2(N2108), .ZN(n13926));
    NOR2X1 U1055 (.A1(N2109), .A2(N2110), .ZN(n13927));
    NOR2X1 U1056 (.A1(N2111), .A2(N2112), .ZN(n13928));
    NOR2X1 U1057 (.A1(N2113), .A2(N2114), .ZN(N13929));
    NANDX1 U1058 (.A1(N2115), .A2(N2116), .ZN(n13930));
    NANDX1 U1059 (.A1(N2117), .A2(N2118), .ZN(n13931));
    NANDX1 U1060 (.A1(N2119), .A2(N2120), .ZN(N13932));
    NOR2X1 U1061 (.A1(N2121), .A2(N2122), .ZN(n13933));
    NOR2X1 U1062 (.A1(N2123), .A2(N2124), .ZN(N13934));
    NANDX1 U1063 (.A1(N2125), .A2(N2126), .ZN(n13935));
    NOR2X1 U1064 (.A1(N2127), .A2(N2128), .ZN(n13936));
    NOR2X1 U1065 (.A1(N2129), .A2(N2130), .ZN(n13937));
    NOR2X1 U1066 (.A1(N2131), .A2(N2132), .ZN(n13938));
    NOR2X1 U1067 (.A1(N2133), .A2(N2134), .ZN(n13939));
    NOR2X1 U1068 (.A1(N2135), .A2(N2136), .ZN(n13940));
    NANDX1 U1069 (.A1(N2137), .A2(N2138), .ZN(N13941));
    NOR2X1 U1070 (.A1(N2139), .A2(N2140), .ZN(n13942));
    NANDX1 U1071 (.A1(N2141), .A2(N2142), .ZN(n13943));
    NOR2X1 U1072 (.A1(N2143), .A2(N2144), .ZN(n13944));
    NOR2X1 U1073 (.A1(N2145), .A2(N2146), .ZN(n13945));
    NOR2X1 U1074 (.A1(N2147), .A2(N2148), .ZN(n13946));
    NANDX1 U1075 (.A1(N2149), .A2(N2150), .ZN(n13947));
    NANDX1 U1076 (.A1(N2151), .A2(N2152), .ZN(n13948));
    NANDX1 U1077 (.A1(N2153), .A2(N2154), .ZN(n13949));
    NANDX1 U1078 (.A1(N2155), .A2(N2156), .ZN(n13950));
    NOR2X1 U1079 (.A1(N2157), .A2(N2158), .ZN(n13951));
    NANDX1 U1080 (.A1(N2159), .A2(N2160), .ZN(n13952));
    NANDX1 U1081 (.A1(N2161), .A2(N2162), .ZN(n13953));
    NOR2X1 U1082 (.A1(N2163), .A2(N2164), .ZN(n13954));
    NANDX1 U1083 (.A1(N2165), .A2(N2166), .ZN(n13955));
    NANDX1 U1084 (.A1(N2167), .A2(N2168), .ZN(N13956));
    NANDX1 U1085 (.A1(N2169), .A2(N2170), .ZN(n13957));
    NANDX1 U1086 (.A1(N2171), .A2(N2172), .ZN(n13958));
    NOR2X1 U1087 (.A1(N2173), .A2(N2174), .ZN(N13959));
    NANDX1 U1088 (.A1(N2175), .A2(N2176), .ZN(n13960));
    NOR2X1 U1089 (.A1(N2177), .A2(N2178), .ZN(n13961));
    NANDX1 U1090 (.A1(N2179), .A2(N2180), .ZN(n13962));
    NANDX1 U1091 (.A1(N2181), .A2(N2182), .ZN(n13963));
    NANDX1 U1092 (.A1(N2183), .A2(N2184), .ZN(n13964));
    NANDX1 U1093 (.A1(N2185), .A2(N2186), .ZN(N13965));
    NOR2X1 U1094 (.A1(N2187), .A2(N2188), .ZN(n13966));
    NANDX1 U1095 (.A1(N2189), .A2(N2190), .ZN(n13967));
    NANDX1 U1096 (.A1(N2191), .A2(N2192), .ZN(n13968));
    NANDX1 U1097 (.A1(N2193), .A2(N2194), .ZN(N13969));
    NANDX1 U1098 (.A1(N2195), .A2(N2196), .ZN(n13970));
    NOR2X1 U1099 (.A1(N2197), .A2(N2198), .ZN(n13971));
    NOR2X1 U1100 (.A1(N2199), .A2(N2200), .ZN(N13972));
    NOR2X1 U1101 (.A1(N2201), .A2(N2202), .ZN(n13973));
    NANDX1 U1102 (.A1(N2203), .A2(N2204), .ZN(n13974));
    NANDX1 U1103 (.A1(N2205), .A2(N2206), .ZN(n13975));
    NOR2X1 U1104 (.A1(N2207), .A2(N2208), .ZN(n13976));
    NANDX1 U1105 (.A1(N2209), .A2(N2210), .ZN(n13977));
    NOR2X1 U1106 (.A1(N2211), .A2(N2212), .ZN(n13978));
    NANDX1 U1107 (.A1(N2213), .A2(N2214), .ZN(n13979));
    NOR2X1 U1108 (.A1(N2215), .A2(N2216), .ZN(n13980));
    NANDX1 U1109 (.A1(N2217), .A2(N2218), .ZN(n13981));
    NANDX1 U1110 (.A1(N2219), .A2(N2220), .ZN(n13982));
    NANDX1 U1111 (.A1(N2221), .A2(N2222), .ZN(n13983));
    NOR2X1 U1112 (.A1(N2223), .A2(N2224), .ZN(n13984));
    NANDX1 U1113 (.A1(N2225), .A2(N2226), .ZN(n13985));
    NOR2X1 U1114 (.A1(N2227), .A2(N2228), .ZN(n13986));
    NOR2X1 U1115 (.A1(N2229), .A2(N2230), .ZN(n13987));
    NOR2X1 U1116 (.A1(N2231), .A2(N2232), .ZN(n13988));
    NANDX1 U1117 (.A1(N2233), .A2(N2234), .ZN(n13989));
    NOR2X1 U1118 (.A1(N2235), .A2(N2236), .ZN(n13990));
    NOR2X1 U1119 (.A1(N2237), .A2(N2238), .ZN(N13991));
    NOR2X1 U1120 (.A1(N2239), .A2(N2240), .ZN(n13992));
    NANDX1 U1121 (.A1(N2241), .A2(N2242), .ZN(n13993));
    NANDX1 U1122 (.A1(N2243), .A2(N2244), .ZN(n13994));
    NANDX1 U1123 (.A1(N2245), .A2(N2246), .ZN(n13995));
    NOR2X1 U1124 (.A1(N2247), .A2(N2248), .ZN(n13996));
    NANDX1 U1125 (.A1(N2249), .A2(N2250), .ZN(n13997));
    NOR2X1 U1126 (.A1(N2251), .A2(N2252), .ZN(n13998));
    NANDX1 U1127 (.A1(N2253), .A2(N2254), .ZN(n13999));
    NOR2X1 U1128 (.A1(N2255), .A2(N2256), .ZN(N14000));
    NANDX1 U1129 (.A1(N2257), .A2(N2258), .ZN(n14001));
    NANDX1 U1130 (.A1(N2259), .A2(N2260), .ZN(n14002));
    NANDX1 U1131 (.A1(N2261), .A2(N2262), .ZN(n14003));
    NANDX1 U1132 (.A1(N2263), .A2(N2264), .ZN(n14004));
    NOR2X1 U1133 (.A1(N2265), .A2(N2266), .ZN(N14005));
    NOR2X1 U1134 (.A1(N2267), .A2(N2268), .ZN(n14006));
    NANDX1 U1135 (.A1(N2269), .A2(N2270), .ZN(n14007));
    NANDX1 U1136 (.A1(N2271), .A2(N2272), .ZN(n14008));
    NOR2X1 U1137 (.A1(N2273), .A2(N2274), .ZN(n14009));
    NANDX1 U1138 (.A1(N2275), .A2(N2276), .ZN(n14010));
    NANDX1 U1139 (.A1(N2277), .A2(N2278), .ZN(n14011));
    NOR2X1 U1140 (.A1(N2279), .A2(N2280), .ZN(n14012));
    NOR2X1 U1141 (.A1(N2281), .A2(N2282), .ZN(n14013));
    NANDX1 U1142 (.A1(N2283), .A2(N2284), .ZN(n14014));
    NOR2X1 U1143 (.A1(N2285), .A2(N2286), .ZN(n14015));
    NOR2X1 U1144 (.A1(N2287), .A2(N2288), .ZN(n14016));
    NANDX1 U1145 (.A1(N2289), .A2(N2290), .ZN(n14017));
    NOR2X1 U1146 (.A1(N2291), .A2(N2292), .ZN(N14018));
    NOR2X1 U1147 (.A1(N2293), .A2(N2294), .ZN(N14019));
    NANDX1 U1148 (.A1(N2295), .A2(N2296), .ZN(n14020));
    NOR2X1 U1149 (.A1(N2297), .A2(N2298), .ZN(n14021));
    NOR2X1 U1150 (.A1(N2299), .A2(N2300), .ZN(n14022));
    NANDX1 U1151 (.A1(N2301), .A2(N2302), .ZN(n14023));
    NANDX1 U1152 (.A1(N2303), .A2(N2304), .ZN(n14024));
    NANDX1 U1153 (.A1(N2305), .A2(N2306), .ZN(n14025));
    NOR2X1 U1154 (.A1(N2307), .A2(N2308), .ZN(n14026));
    NANDX1 U1155 (.A1(N2309), .A2(N2310), .ZN(n14027));
    NANDX1 U1156 (.A1(N2311), .A2(N2312), .ZN(n14028));
    NOR2X1 U1157 (.A1(N2313), .A2(N2314), .ZN(n14029));
    NANDX1 U1158 (.A1(N2315), .A2(N2316), .ZN(n14030));
    NANDX1 U1159 (.A1(N2317), .A2(N2318), .ZN(n14031));
    NANDX1 U1160 (.A1(N2319), .A2(N2320), .ZN(n14032));
    NOR2X1 U1161 (.A1(N2321), .A2(N2322), .ZN(N14033));
    NOR2X1 U1162 (.A1(N2323), .A2(N2324), .ZN(N14034));
    NANDX1 U1163 (.A1(N2325), .A2(N2326), .ZN(n14035));
    NANDX1 U1164 (.A1(N2327), .A2(N2328), .ZN(n14036));
    NOR2X1 U1165 (.A1(N2329), .A2(N2330), .ZN(N14037));
    NOR2X1 U1166 (.A1(N2331), .A2(N2332), .ZN(n14038));
    NOR2X1 U1167 (.A1(N2333), .A2(N2334), .ZN(n14039));
    NANDX1 U1168 (.A1(N2335), .A2(N2336), .ZN(N14040));
    NANDX1 U1169 (.A1(N2337), .A2(N2338), .ZN(n14041));
    NOR2X1 U1170 (.A1(N2339), .A2(N2340), .ZN(n14042));
    NANDX1 U1171 (.A1(N2341), .A2(N2342), .ZN(n14043));
    NOR2X1 U1172 (.A1(N2343), .A2(N2344), .ZN(n14044));
    NANDX1 U1173 (.A1(N2345), .A2(N2346), .ZN(N14045));
    NANDX1 U1174 (.A1(N2347), .A2(N2348), .ZN(n14046));
    NOR2X1 U1175 (.A1(N2349), .A2(N2350), .ZN(n14047));
    NOR2X1 U1176 (.A1(N2351), .A2(N2352), .ZN(n14048));
    NOR2X1 U1177 (.A1(N2353), .A2(N2354), .ZN(n14049));
    NOR2X1 U1178 (.A1(N2355), .A2(N2356), .ZN(n14050));
    NANDX1 U1179 (.A1(N2357), .A2(N2358), .ZN(n14051));
    NOR2X1 U1180 (.A1(N2359), .A2(N2360), .ZN(N14052));
    NANDX1 U1181 (.A1(N2361), .A2(N2362), .ZN(n14053));
    NOR2X1 U1182 (.A1(N2363), .A2(N2364), .ZN(n14054));
    NOR2X1 U1183 (.A1(N2365), .A2(N2366), .ZN(n14055));
    NOR2X1 U1184 (.A1(N2367), .A2(N2368), .ZN(N14056));
    NOR2X1 U1185 (.A1(N2369), .A2(N2370), .ZN(n14057));
    NANDX1 U1186 (.A1(N2371), .A2(N2372), .ZN(n14058));
    NANDX1 U1187 (.A1(N2373), .A2(N2374), .ZN(n14059));
    NOR2X1 U1188 (.A1(N2375), .A2(N2376), .ZN(N14060));
    NOR2X1 U1189 (.A1(N2377), .A2(N2378), .ZN(n14061));
    NANDX1 U1190 (.A1(N2379), .A2(N2380), .ZN(n14062));
    NOR2X1 U1191 (.A1(N2381), .A2(N2382), .ZN(n14063));
    NANDX1 U1192 (.A1(N2383), .A2(N2384), .ZN(n14064));
    NANDX1 U1193 (.A1(N2385), .A2(N2386), .ZN(n14065));
    NANDX1 U1194 (.A1(N2387), .A2(N2388), .ZN(n14066));
    NOR2X1 U1195 (.A1(N2389), .A2(N2390), .ZN(n14067));
    NOR2X1 U1196 (.A1(N2391), .A2(N2392), .ZN(n14068));
    NANDX1 U1197 (.A1(N2393), .A2(N2394), .ZN(n14069));
    NOR2X1 U1198 (.A1(N2395), .A2(N2396), .ZN(n14070));
    NANDX1 U1199 (.A1(N2397), .A2(N2398), .ZN(n14071));
    NANDX1 U1200 (.A1(N2399), .A2(N2400), .ZN(n14072));
    NOR2X1 U1201 (.A1(N2401), .A2(N2402), .ZN(n14073));
    NOR2X1 U1202 (.A1(N2403), .A2(N2404), .ZN(n14074));
    NANDX1 U1203 (.A1(N2405), .A2(N2406), .ZN(n14075));
    NANDX1 U1204 (.A1(N2407), .A2(N2408), .ZN(n14076));
    NANDX1 U1205 (.A1(N2409), .A2(N2410), .ZN(n14077));
    NANDX1 U1206 (.A1(N2411), .A2(N2412), .ZN(n14078));
    NOR2X1 U1207 (.A1(N2413), .A2(N2414), .ZN(N14079));
    NANDX1 U1208 (.A1(N2415), .A2(N2416), .ZN(n14080));
    NANDX1 U1209 (.A1(N2417), .A2(N2418), .ZN(n14081));
    NANDX1 U1210 (.A1(N2419), .A2(N2420), .ZN(n14082));
    NOR2X1 U1211 (.A1(N2421), .A2(N2422), .ZN(n14083));
    NOR2X1 U1212 (.A1(N2423), .A2(N2424), .ZN(N14084));
    NOR2X1 U1213 (.A1(N2425), .A2(N2426), .ZN(n14085));
    NOR2X1 U1214 (.A1(N2427), .A2(N2428), .ZN(n14086));
    NANDX1 U1215 (.A1(N2429), .A2(N2430), .ZN(N14087));
    NOR2X1 U1216 (.A1(N2431), .A2(N2432), .ZN(n14088));
    NANDX1 U1217 (.A1(N2433), .A2(N2434), .ZN(n14089));
    NOR2X1 U1218 (.A1(N2435), .A2(N2436), .ZN(n14090));
    NANDX1 U1219 (.A1(N2437), .A2(N2438), .ZN(n14091));
    NOR2X1 U1220 (.A1(N2439), .A2(N2440), .ZN(n14092));
    NANDX1 U1221 (.A1(N2441), .A2(N2442), .ZN(n14093));
    NANDX1 U1222 (.A1(N2443), .A2(N2444), .ZN(n14094));
    NANDX1 U1223 (.A1(N2445), .A2(N2446), .ZN(n14095));
    NANDX1 U1224 (.A1(N2447), .A2(N2448), .ZN(n14096));
    NOR2X1 U1225 (.A1(N2449), .A2(N2450), .ZN(n14097));
    NANDX1 U1226 (.A1(N2451), .A2(N2452), .ZN(n14098));
    NANDX1 U1227 (.A1(N2453), .A2(N2454), .ZN(n14099));
    NANDX1 U1228 (.A1(N2455), .A2(N2456), .ZN(N14100));
    NANDX1 U1229 (.A1(N2457), .A2(N2458), .ZN(N14101));
    NOR2X1 U1230 (.A1(N2459), .A2(N2460), .ZN(n14102));
    NOR2X1 U1231 (.A1(N2461), .A2(N2462), .ZN(n14103));
    NOR2X1 U1232 (.A1(N2463), .A2(N2464), .ZN(N14104));
    NOR2X1 U1233 (.A1(N2465), .A2(N2466), .ZN(n14105));
    NANDX1 U1234 (.A1(N2467), .A2(N2468), .ZN(n14106));
    NANDX1 U1235 (.A1(N2469), .A2(N2470), .ZN(N14107));
    NANDX1 U1236 (.A1(N2471), .A2(N2472), .ZN(n14108));
    NOR2X1 U1237 (.A1(N2473), .A2(N2474), .ZN(n14109));
    NANDX1 U1238 (.A1(N2475), .A2(N2476), .ZN(n14110));
    NANDX1 U1239 (.A1(N2477), .A2(N2478), .ZN(n14111));
    NOR2X1 U1240 (.A1(N2479), .A2(N2480), .ZN(n14112));
    NANDX1 U1241 (.A1(N2481), .A2(N2482), .ZN(N14113));
    NANDX1 U1242 (.A1(N2483), .A2(N2484), .ZN(n14114));
    NOR2X1 U1243 (.A1(N2485), .A2(N2486), .ZN(n14115));
    NANDX1 U1244 (.A1(N2487), .A2(N2488), .ZN(n14116));
    NANDX1 U1245 (.A1(N2489), .A2(N2490), .ZN(n14117));
    NANDX1 U1246 (.A1(N2491), .A2(N2492), .ZN(n14118));
    NANDX1 U1247 (.A1(N2493), .A2(N2494), .ZN(N14119));
    NOR2X1 U1248 (.A1(N2495), .A2(N2496), .ZN(n14120));
    NOR2X1 U1249 (.A1(N2497), .A2(N2498), .ZN(n14121));
    NOR2X1 U1250 (.A1(N2499), .A2(N2500), .ZN(n14122));
    NOR2X1 U1251 (.A1(N2501), .A2(N2502), .ZN(n14123));
    NANDX1 U1252 (.A1(N2503), .A2(N2504), .ZN(N14124));
    NANDX1 U1253 (.A1(N2505), .A2(N2506), .ZN(N14125));
    NANDX1 U1254 (.A1(N2507), .A2(N2508), .ZN(N14126));
    NOR2X1 U1255 (.A1(N2509), .A2(N2510), .ZN(n14127));
    NANDX1 U1256 (.A1(N2511), .A2(N2512), .ZN(n14128));
    NOR2X1 U1257 (.A1(N2513), .A2(N2514), .ZN(n14129));
    NANDX1 U1258 (.A1(N2515), .A2(N2516), .ZN(n14130));
    NANDX1 U1259 (.A1(N2517), .A2(N2518), .ZN(n14131));
    NOR2X1 U1260 (.A1(N2519), .A2(N2520), .ZN(n14132));
    NANDX1 U1261 (.A1(N2521), .A2(N2522), .ZN(n14133));
    NANDX1 U1262 (.A1(N2523), .A2(N2524), .ZN(n14134));
    NOR2X1 U1263 (.A1(N2525), .A2(N2526), .ZN(n14135));
    NANDX1 U1264 (.A1(N2527), .A2(N2528), .ZN(n14136));
    NANDX1 U1265 (.A1(N2529), .A2(N2530), .ZN(n14137));
    NANDX1 U1266 (.A1(N2531), .A2(N2532), .ZN(n14138));
    NANDX1 U1267 (.A1(N2533), .A2(N2534), .ZN(n14139));
    NANDX1 U1268 (.A1(N2535), .A2(N2536), .ZN(n14140));
    NANDX1 U1269 (.A1(N2537), .A2(N2538), .ZN(n14141));
    NOR2X1 U1270 (.A1(N2539), .A2(N2540), .ZN(n14142));
    NANDX1 U1271 (.A1(N2541), .A2(N2542), .ZN(n14143));
    NOR2X1 U1272 (.A1(N2543), .A2(N2544), .ZN(n14144));
    NANDX1 U1273 (.A1(N2545), .A2(N2546), .ZN(n14145));
    NOR2X1 U1274 (.A1(N2547), .A2(N2548), .ZN(n14146));
    NANDX1 U1275 (.A1(N2549), .A2(N2550), .ZN(N14147));
    NOR2X1 U1276 (.A1(N2551), .A2(N2552), .ZN(n14148));
    NANDX1 U1277 (.A1(N2553), .A2(N2554), .ZN(n14149));
    NOR2X1 U1278 (.A1(N2555), .A2(N2556), .ZN(n14150));
    NOR2X1 U1279 (.A1(N2557), .A2(N2558), .ZN(N14151));
    NANDX1 U1280 (.A1(N2559), .A2(N2560), .ZN(n14152));
    NANDX1 U1281 (.A1(N2561), .A2(N2562), .ZN(n14153));
    NANDX1 U1282 (.A1(N2563), .A2(N2564), .ZN(n14154));
    NANDX1 U1283 (.A1(N2565), .A2(N2566), .ZN(n14155));
    NOR2X1 U1284 (.A1(N2567), .A2(N2568), .ZN(n14156));
    NOR2X1 U1285 (.A1(N2569), .A2(N2570), .ZN(n14157));
    NANDX1 U1286 (.A1(N2571), .A2(N2572), .ZN(N14158));
    NOR2X1 U1287 (.A1(N2573), .A2(N2574), .ZN(N14159));
    NANDX1 U1288 (.A1(N2575), .A2(N2576), .ZN(n14160));
    NANDX1 U1289 (.A1(N2577), .A2(N2578), .ZN(N14161));
    NANDX1 U1290 (.A1(N2579), .A2(N2580), .ZN(n14162));
    NANDX1 U1291 (.A1(N2581), .A2(N2582), .ZN(n14163));
    NOR2X1 U1292 (.A1(N2583), .A2(N2584), .ZN(n14164));
    NOR2X1 U1293 (.A1(N2585), .A2(N2586), .ZN(N14165));
    NANDX1 U1294 (.A1(N2587), .A2(N2588), .ZN(n14166));
    NOR2X1 U1295 (.A1(N2589), .A2(N2590), .ZN(n14167));
    NANDX1 U1296 (.A1(N2591), .A2(N2592), .ZN(n14168));
    NOR2X1 U1297 (.A1(N2593), .A2(N2594), .ZN(n14169));
    NANDX1 U1298 (.A1(N2595), .A2(N2596), .ZN(n14170));
    NANDX1 U1299 (.A1(N2597), .A2(N2598), .ZN(N14171));
    NANDX1 U1300 (.A1(N2599), .A2(N2600), .ZN(n14172));
    NANDX1 U1301 (.A1(N2601), .A2(N2602), .ZN(n14173));
    NOR2X1 U1302 (.A1(N2603), .A2(N2604), .ZN(N14174));
    NANDX1 U1303 (.A1(N2605), .A2(N2606), .ZN(n14175));
    NOR2X1 U1304 (.A1(N2607), .A2(N2608), .ZN(n14176));
    NOR2X1 U1305 (.A1(N2609), .A2(N2610), .ZN(n14177));
    NOR2X1 U1306 (.A1(N2611), .A2(N2612), .ZN(n14178));
    NOR2X1 U1307 (.A1(N2613), .A2(N2614), .ZN(n14179));
    NOR2X1 U1308 (.A1(N2615), .A2(N2616), .ZN(N14180));
    NANDX1 U1309 (.A1(N2617), .A2(N2618), .ZN(n14181));
    NOR2X1 U1310 (.A1(N2619), .A2(N2620), .ZN(n14182));
    NANDX1 U1311 (.A1(N2621), .A2(N2622), .ZN(n14183));
    NOR2X1 U1312 (.A1(N2623), .A2(N2624), .ZN(n14184));
    NANDX1 U1313 (.A1(N2625), .A2(N2626), .ZN(N14185));
    NOR2X1 U1314 (.A1(N2627), .A2(N2628), .ZN(N14186));
    NOR2X1 U1315 (.A1(N2629), .A2(N2630), .ZN(N14187));
    NOR2X1 U1316 (.A1(N2631), .A2(N2632), .ZN(n14188));
    NOR2X1 U1317 (.A1(N2633), .A2(N2634), .ZN(n14189));
    NOR2X1 U1318 (.A1(N2635), .A2(N2636), .ZN(n14190));
    NANDX1 U1319 (.A1(N2637), .A2(N2638), .ZN(n14191));
    NANDX1 U1320 (.A1(N2639), .A2(N2640), .ZN(n14192));
    NANDX1 U1321 (.A1(N2641), .A2(N2642), .ZN(n14193));
    NOR2X1 U1322 (.A1(N2643), .A2(N2644), .ZN(n14194));
    NANDX1 U1323 (.A1(N2645), .A2(N2646), .ZN(n14195));
    NOR2X1 U1324 (.A1(N2647), .A2(N2648), .ZN(n14196));
    NANDX1 U1325 (.A1(N2649), .A2(N2650), .ZN(n14197));
    NANDX1 U1326 (.A1(N2651), .A2(N2652), .ZN(n14198));
    NANDX1 U1327 (.A1(N2653), .A2(N2654), .ZN(n14199));
    NANDX1 U1328 (.A1(N2655), .A2(N2656), .ZN(n14200));
    NOR2X1 U1329 (.A1(N2657), .A2(N2658), .ZN(n14201));
    NOR2X1 U1330 (.A1(N2659), .A2(N2660), .ZN(n14202));
    NANDX1 U1331 (.A1(N2661), .A2(N2662), .ZN(N14203));
    NANDX1 U1332 (.A1(N2663), .A2(N2664), .ZN(n14204));
    NANDX1 U1333 (.A1(N2665), .A2(N2666), .ZN(N14205));
    NOR2X1 U1334 (.A1(N2667), .A2(N2668), .ZN(n14206));
    NANDX1 U1335 (.A1(N2669), .A2(N2670), .ZN(N14207));
    NANDX1 U1336 (.A1(N2671), .A2(N2672), .ZN(N14208));
    NANDX1 U1337 (.A1(N2673), .A2(N2674), .ZN(n14209));
    NANDX1 U1338 (.A1(N2675), .A2(N2676), .ZN(n14210));
    NANDX1 U1339 (.A1(N2677), .A2(N2678), .ZN(n14211));
    NOR2X1 U1340 (.A1(N2679), .A2(N2680), .ZN(N14212));
    NOR2X1 U1341 (.A1(N2681), .A2(N2682), .ZN(n14213));
    NANDX1 U1342 (.A1(N2683), .A2(N2684), .ZN(N14214));
    NOR2X1 U1343 (.A1(N2685), .A2(N2686), .ZN(N14215));
    NANDX1 U1344 (.A1(N2687), .A2(N2688), .ZN(N14216));
    NANDX1 U1345 (.A1(N2689), .A2(N2690), .ZN(N14217));
    NOR2X1 U1346 (.A1(N2691), .A2(N2692), .ZN(n14218));
    NANDX1 U1347 (.A1(N2693), .A2(N2694), .ZN(N14219));
    NANDX1 U1348 (.A1(N2695), .A2(N2696), .ZN(n14220));
    NANDX1 U1349 (.A1(N2697), .A2(N2698), .ZN(n14221));
    NOR2X1 U1350 (.A1(N2699), .A2(N2700), .ZN(N14222));
    NOR2X1 U1351 (.A1(N2701), .A2(N2702), .ZN(n14223));
    NOR2X1 U1352 (.A1(N2703), .A2(N2704), .ZN(n14224));
    NOR2X1 U1353 (.A1(N2705), .A2(N2706), .ZN(n14225));
    NOR2X1 U1354 (.A1(N2707), .A2(N2708), .ZN(n14226));
    NOR2X1 U1355 (.A1(N2709), .A2(N2710), .ZN(n14227));
    NANDX1 U1356 (.A1(N2711), .A2(N2712), .ZN(n14228));
    NANDX1 U1357 (.A1(N2713), .A2(N2714), .ZN(n14229));
    NOR2X1 U1358 (.A1(N2715), .A2(N2716), .ZN(n14230));
    NANDX1 U1359 (.A1(N2717), .A2(N2718), .ZN(n14231));
    NOR2X1 U1360 (.A1(N2719), .A2(N2720), .ZN(n14232));
    NOR2X1 U1361 (.A1(N2721), .A2(N2722), .ZN(n14233));
    NOR2X1 U1362 (.A1(N2723), .A2(N2724), .ZN(N14234));
    NANDX1 U1363 (.A1(N2725), .A2(N2726), .ZN(n14235));
    NANDX1 U1364 (.A1(N2727), .A2(N2728), .ZN(n14236));
    NOR2X1 U1365 (.A1(N2729), .A2(N2730), .ZN(n14237));
    NANDX1 U1366 (.A1(N2731), .A2(N2732), .ZN(n14238));
    NANDX1 U1367 (.A1(N2733), .A2(N2734), .ZN(n14239));
    NANDX1 U1368 (.A1(N2735), .A2(N2736), .ZN(n14240));
    NOR2X1 U1369 (.A1(N2737), .A2(N2738), .ZN(n14241));
    NOR2X1 U1370 (.A1(N2739), .A2(N2740), .ZN(n14242));
    NANDX1 U1371 (.A1(N2741), .A2(N2742), .ZN(N14243));
    NOR2X1 U1372 (.A1(N2743), .A2(N2744), .ZN(n14244));
    NANDX1 U1373 (.A1(N2745), .A2(N2746), .ZN(n14245));
    NANDX1 U1374 (.A1(N2747), .A2(N2748), .ZN(n14246));
    NOR2X1 U1375 (.A1(N2749), .A2(N2750), .ZN(n14247));
    NANDX1 U1376 (.A1(N2751), .A2(N2752), .ZN(n14248));
    NOR2X1 U1377 (.A1(N2753), .A2(N2754), .ZN(n14249));
    NANDX1 U1378 (.A1(N2755), .A2(N2756), .ZN(n14250));
    NOR2X1 U1379 (.A1(N2757), .A2(N2758), .ZN(n14251));
    NANDX1 U1380 (.A1(N2759), .A2(N2760), .ZN(n14252));
    NOR2X1 U1381 (.A1(N2761), .A2(N2762), .ZN(n14253));
    NANDX1 U1382 (.A1(N2763), .A2(N2764), .ZN(n14254));
    NANDX1 U1383 (.A1(N2765), .A2(N2766), .ZN(n14255));
    NOR2X1 U1384 (.A1(N2767), .A2(N2768), .ZN(n14256));
    NANDX1 U1385 (.A1(N2769), .A2(N2770), .ZN(n14257));
    NOR2X1 U1386 (.A1(N2771), .A2(N2772), .ZN(n14258));
    NOR2X1 U1387 (.A1(N2773), .A2(N2774), .ZN(n14259));
    NOR2X1 U1388 (.A1(N2775), .A2(N2776), .ZN(n14260));
    NOR2X1 U1389 (.A1(N2777), .A2(N2778), .ZN(n14261));
    NANDX1 U1390 (.A1(N2779), .A2(N2780), .ZN(n14262));
    NOR2X1 U1391 (.A1(N2781), .A2(N2782), .ZN(n14263));
    NOR2X1 U1392 (.A1(N2783), .A2(N2784), .ZN(n14264));
    NANDX1 U1393 (.A1(N2785), .A2(N2786), .ZN(n14265));
    NOR2X1 U1394 (.A1(N2787), .A2(N2788), .ZN(n14266));
    NOR2X1 U1395 (.A1(N2789), .A2(N2790), .ZN(n14267));
    NANDX1 U1396 (.A1(N2791), .A2(N2792), .ZN(n14268));
    NANDX1 U1397 (.A1(N2793), .A2(N2794), .ZN(N14269));
    NANDX1 U1398 (.A1(N2795), .A2(N2796), .ZN(n14270));
    NANDX1 U1399 (.A1(N2797), .A2(N2798), .ZN(n14271));
    NANDX1 U1400 (.A1(N2799), .A2(N2800), .ZN(n14272));
    NANDX1 U1401 (.A1(N2801), .A2(N2802), .ZN(n14273));
    NOR2X1 U1402 (.A1(N2803), .A2(N2804), .ZN(N14274));
    NOR2X1 U1403 (.A1(N2805), .A2(N2806), .ZN(N14275));
    NANDX1 U1404 (.A1(N2807), .A2(N2808), .ZN(n14276));
    NOR2X1 U1405 (.A1(N2809), .A2(N2810), .ZN(n14277));
    NOR2X1 U1406 (.A1(N2811), .A2(N2812), .ZN(n14278));
    NOR2X1 U1407 (.A1(N2813), .A2(N2814), .ZN(n14279));
    NOR2X1 U1408 (.A1(N2815), .A2(N2816), .ZN(N14280));
    NANDX1 U1409 (.A1(N2817), .A2(N2818), .ZN(n14281));
    NOR2X1 U1410 (.A1(N2819), .A2(N2820), .ZN(n14282));
    NANDX1 U1411 (.A1(N2821), .A2(N2822), .ZN(n14283));
    NANDX1 U1412 (.A1(N2823), .A2(N2824), .ZN(n14284));
    NANDX1 U1413 (.A1(N2825), .A2(N2826), .ZN(n14285));
    NOR2X1 U1414 (.A1(N2827), .A2(N2828), .ZN(n14286));
    NOR2X1 U1415 (.A1(N2829), .A2(N2830), .ZN(n14287));
    NOR2X1 U1416 (.A1(N2831), .A2(N2832), .ZN(N14288));
    NOR2X1 U1417 (.A1(N2833), .A2(N2834), .ZN(N14289));
    NOR2X1 U1418 (.A1(N2835), .A2(N2836), .ZN(n14290));
    NANDX1 U1419 (.A1(N2837), .A2(N2838), .ZN(N14291));
    NOR2X1 U1420 (.A1(N2839), .A2(N2840), .ZN(n14292));
    NANDX1 U1421 (.A1(N2841), .A2(N2842), .ZN(n14293));
    NANDX1 U1422 (.A1(N2843), .A2(N2844), .ZN(n14294));
    NANDX1 U1423 (.A1(N2845), .A2(N2846), .ZN(n14295));
    NOR2X1 U1424 (.A1(N2847), .A2(N2848), .ZN(N14296));
    NANDX1 U1425 (.A1(N2849), .A2(N2850), .ZN(n14297));
    NANDX1 U1426 (.A1(N2851), .A2(N2852), .ZN(N14298));
    NANDX1 U1427 (.A1(N2853), .A2(N2854), .ZN(n14299));
    NOR2X1 U1428 (.A1(N2855), .A2(N2856), .ZN(n14300));
    NOR2X1 U1429 (.A1(N2857), .A2(N2858), .ZN(n14301));
    NOR2X1 U1430 (.A1(N2859), .A2(N2860), .ZN(n14302));
    NOR2X1 U1431 (.A1(N2861), .A2(N2862), .ZN(n14303));
    NANDX1 U1432 (.A1(N2863), .A2(N2864), .ZN(n14304));
    NANDX1 U1433 (.A1(N2865), .A2(N2866), .ZN(n14305));
    NOR2X1 U1434 (.A1(N2867), .A2(N2868), .ZN(n14306));
    NOR2X1 U1435 (.A1(N2869), .A2(N2870), .ZN(n14307));
    NANDX1 U1436 (.A1(N2871), .A2(N2872), .ZN(n14308));
    NOR2X1 U1437 (.A1(N2873), .A2(N2874), .ZN(n14309));
    NOR2X1 U1438 (.A1(N2875), .A2(N2876), .ZN(n14310));
    NANDX1 U1439 (.A1(N2877), .A2(N2878), .ZN(N14311));
    NANDX1 U1440 (.A1(N2879), .A2(N2880), .ZN(n14312));
    NANDX1 U1441 (.A1(N2881), .A2(N2882), .ZN(n14313));
    NOR2X1 U1442 (.A1(N2883), .A2(N2884), .ZN(n14314));
    NANDX1 U1443 (.A1(N2885), .A2(N2886), .ZN(n14315));
    NOR2X1 U1444 (.A1(N2887), .A2(N2888), .ZN(n14316));
    NOR2X1 U1445 (.A1(N2889), .A2(N2890), .ZN(n14317));
    NANDX1 U1446 (.A1(N2891), .A2(N2892), .ZN(N14318));
    NANDX1 U1447 (.A1(N2893), .A2(N2894), .ZN(n14319));
    NANDX1 U1448 (.A1(N2895), .A2(N2896), .ZN(n14320));
    NANDX1 U1449 (.A1(N2897), .A2(N2898), .ZN(N14321));
    NOR2X1 U1450 (.A1(N2899), .A2(N2900), .ZN(n14322));
    NANDX1 U1451 (.A1(N2901), .A2(N2902), .ZN(n14323));
    NOR2X1 U1452 (.A1(N2903), .A2(N2904), .ZN(n14324));
    NANDX1 U1453 (.A1(N2905), .A2(N2906), .ZN(n14325));
    NOR2X1 U1454 (.A1(N2907), .A2(N2908), .ZN(n14326));
    NOR2X1 U1455 (.A1(N2909), .A2(N2910), .ZN(n14327));
    NANDX1 U1456 (.A1(N2911), .A2(N2912), .ZN(n14328));
    NANDX1 U1457 (.A1(N2913), .A2(N2914), .ZN(n14329));
    NANDX1 U1458 (.A1(N2915), .A2(N2916), .ZN(n14330));
    NANDX1 U1459 (.A1(N2917), .A2(N2918), .ZN(n14331));
    NANDX1 U1460 (.A1(N2919), .A2(N2920), .ZN(n14332));
    NOR2X1 U1461 (.A1(N2921), .A2(N2922), .ZN(n14333));
    NANDX1 U1462 (.A1(N2923), .A2(N2924), .ZN(n14334));
    NANDX1 U1463 (.A1(N2925), .A2(N2926), .ZN(n14335));
    NANDX1 U1464 (.A1(N2927), .A2(N2928), .ZN(n14336));
    NANDX1 U1465 (.A1(N2929), .A2(N2930), .ZN(N14337));
    NANDX1 U1466 (.A1(N2931), .A2(N2932), .ZN(n14338));
    NOR2X1 U1467 (.A1(N2933), .A2(N2934), .ZN(n14339));
    NANDX1 U1468 (.A1(N2935), .A2(N2936), .ZN(n14340));
    NOR2X1 U1469 (.A1(N2937), .A2(N2938), .ZN(n14341));
    NANDX1 U1470 (.A1(N2939), .A2(N2940), .ZN(n14342));
    NANDX1 U1471 (.A1(N2941), .A2(N2942), .ZN(n14343));
    NANDX1 U1472 (.A1(N2943), .A2(N2944), .ZN(n14344));
    NANDX1 U1473 (.A1(N2945), .A2(N2946), .ZN(n14345));
    NOR2X1 U1474 (.A1(N2947), .A2(N2948), .ZN(n14346));
    NANDX1 U1475 (.A1(N2949), .A2(N2950), .ZN(N14347));
    NANDX1 U1476 (.A1(N2951), .A2(N2952), .ZN(n14348));
    NANDX1 U1477 (.A1(N2953), .A2(N2954), .ZN(n14349));
    NOR2X1 U1478 (.A1(N2955), .A2(N2956), .ZN(n14350));
    NOR2X1 U1479 (.A1(N2957), .A2(N2958), .ZN(n14351));
    NOR2X1 U1480 (.A1(N2959), .A2(N2960), .ZN(N14352));
    NOR2X1 U1481 (.A1(N2961), .A2(N2962), .ZN(n14353));
    NOR2X1 U1482 (.A1(N2963), .A2(N2964), .ZN(N14354));
    NOR2X1 U1483 (.A1(N2965), .A2(N2966), .ZN(N14355));
    NOR2X1 U1484 (.A1(N2967), .A2(N2968), .ZN(n14356));
    NOR2X1 U1485 (.A1(N2969), .A2(N2970), .ZN(n14357));
    NOR2X1 U1486 (.A1(N2971), .A2(N2972), .ZN(n14358));
    NANDX1 U1487 (.A1(N2973), .A2(N2974), .ZN(N14359));
    NOR2X1 U1488 (.A1(N2975), .A2(N2976), .ZN(n14360));
    NANDX1 U1489 (.A1(N2977), .A2(N2978), .ZN(N14361));
    NOR2X1 U1490 (.A1(N2979), .A2(N2980), .ZN(n14362));
    NANDX1 U1491 (.A1(N2981), .A2(N2982), .ZN(n14363));
    NANDX1 U1492 (.A1(N2983), .A2(N2984), .ZN(n14364));
    NOR2X1 U1493 (.A1(N2985), .A2(N2986), .ZN(n14365));
    NOR2X1 U1494 (.A1(N2987), .A2(N2988), .ZN(n14366));
    NOR2X1 U1495 (.A1(N2989), .A2(N2990), .ZN(n14367));
    NANDX1 U1496 (.A1(N2991), .A2(N2992), .ZN(N14368));
    NOR2X1 U1497 (.A1(N2993), .A2(N2994), .ZN(n14369));
    NOR2X1 U1498 (.A1(N2995), .A2(N2996), .ZN(n14370));
    NANDX1 U1499 (.A1(N2997), .A2(N2998), .ZN(n14371));
    NOR2X1 U1500 (.A1(N2999), .A2(N3000), .ZN(n14372));
    NANDX1 U1501 (.A1(N3001), .A2(N3002), .ZN(n14373));
    NOR2X1 U1502 (.A1(N3003), .A2(N3004), .ZN(n14374));
    NANDX1 U1503 (.A1(N3005), .A2(N3006), .ZN(n14375));
    NOR2X1 U1504 (.A1(N3007), .A2(N3008), .ZN(n14376));
    NOR2X1 U1505 (.A1(N3009), .A2(N3010), .ZN(n14377));
    NOR2X1 U1506 (.A1(N3011), .A2(N3012), .ZN(n14378));
    NOR2X1 U1507 (.A1(N3013), .A2(N3014), .ZN(n14379));
    NANDX1 U1508 (.A1(N3015), .A2(N3016), .ZN(n14380));
    NANDX1 U1509 (.A1(N3017), .A2(N3018), .ZN(n14381));
    NOR2X1 U1510 (.A1(N3019), .A2(N3020), .ZN(N14382));
    NANDX1 U1511 (.A1(N3021), .A2(N3022), .ZN(n14383));
    NANDX1 U1512 (.A1(N3023), .A2(N3024), .ZN(n14384));
    NOR2X1 U1513 (.A1(N3025), .A2(N3026), .ZN(N14385));
    NANDX1 U1514 (.A1(N3027), .A2(N3028), .ZN(n14386));
    NANDX1 U1515 (.A1(N3029), .A2(N3030), .ZN(n14387));
    NANDX1 U1516 (.A1(N3031), .A2(N3032), .ZN(n14388));
    NANDX1 U1517 (.A1(N3033), .A2(N3034), .ZN(n14389));
    NOR2X1 U1518 (.A1(N3035), .A2(N3036), .ZN(n14390));
    NANDX1 U1519 (.A1(N3037), .A2(N3038), .ZN(n14391));
    NOR2X1 U1520 (.A1(N3039), .A2(N3040), .ZN(n14392));
    NANDX1 U1521 (.A1(N3041), .A2(N3042), .ZN(n14393));
    NOR2X1 U1522 (.A1(N3043), .A2(N3044), .ZN(n14394));
    NOR2X1 U1523 (.A1(N3045), .A2(N3046), .ZN(n14395));
    NANDX1 U1524 (.A1(N3047), .A2(N3048), .ZN(n14396));
    NANDX1 U1525 (.A1(N3049), .A2(N3050), .ZN(n14397));
    NOR2X1 U1526 (.A1(N3051), .A2(N3052), .ZN(n14398));
    NOR2X1 U1527 (.A1(N3053), .A2(N3054), .ZN(n14399));
    NANDX1 U1528 (.A1(N3055), .A2(N3056), .ZN(n14400));
    NANDX1 U1529 (.A1(N3057), .A2(N3058), .ZN(n14401));
    NANDX1 U1530 (.A1(N3059), .A2(N3060), .ZN(n14402));
    NANDX1 U1531 (.A1(N3061), .A2(N3062), .ZN(n14403));
    NOR2X1 U1532 (.A1(N3063), .A2(N3064), .ZN(n14404));
    NANDX1 U1533 (.A1(N3065), .A2(N3066), .ZN(n14405));
    NOR2X1 U1534 (.A1(N3067), .A2(N3068), .ZN(n14406));
    NANDX1 U1535 (.A1(N3069), .A2(N3070), .ZN(n14407));
    NANDX1 U1536 (.A1(N3071), .A2(N3072), .ZN(n14408));
    NOR2X1 U1537 (.A1(N3073), .A2(N3074), .ZN(n14409));
    NANDX1 U1538 (.A1(N3075), .A2(N3076), .ZN(n14410));
    NOR2X1 U1539 (.A1(N3077), .A2(N3078), .ZN(n14411));
    NANDX1 U1540 (.A1(N3079), .A2(N3080), .ZN(n14412));
    NANDX1 U1541 (.A1(N3081), .A2(N3082), .ZN(n14413));
    NANDX1 U1542 (.A1(N3083), .A2(N3084), .ZN(n14414));
    NANDX1 U1543 (.A1(N3085), .A2(N3086), .ZN(n14415));
    NOR2X1 U1544 (.A1(N3087), .A2(N3088), .ZN(N14416));
    NOR2X1 U1545 (.A1(N3089), .A2(N3090), .ZN(N14417));
    NOR2X1 U1546 (.A1(N3091), .A2(N3092), .ZN(n14418));
    NANDX1 U1547 (.A1(N3093), .A2(N3094), .ZN(n14419));
    NANDX1 U1548 (.A1(N3095), .A2(N3096), .ZN(n14420));
    NANDX1 U1549 (.A1(N3097), .A2(N3098), .ZN(n14421));
    NOR2X1 U1550 (.A1(N3099), .A2(N3100), .ZN(n14422));
    NOR2X1 U1551 (.A1(N3101), .A2(N3102), .ZN(n14423));
    NOR2X1 U1552 (.A1(N3103), .A2(N3104), .ZN(N14424));
    NOR2X1 U1553 (.A1(N3105), .A2(N3106), .ZN(n14425));
    NOR2X1 U1554 (.A1(N3107), .A2(N3108), .ZN(n14426));
    NANDX1 U1555 (.A1(N3109), .A2(N3110), .ZN(n14427));
    NANDX1 U1556 (.A1(N3111), .A2(N3112), .ZN(N14428));
    NOR2X1 U1557 (.A1(N3113), .A2(N3114), .ZN(N14429));
    NANDX1 U1558 (.A1(N3115), .A2(N3116), .ZN(n14430));
    NOR2X1 U1559 (.A1(N3117), .A2(N3118), .ZN(n14431));
    NANDX1 U1560 (.A1(N3119), .A2(N3120), .ZN(n14432));
    NANDX1 U1561 (.A1(N3121), .A2(N3122), .ZN(N14433));
    NANDX1 U1562 (.A1(N3123), .A2(N3124), .ZN(n14434));
    NOR2X1 U1563 (.A1(N3125), .A2(N3126), .ZN(n14435));
    NOR2X1 U1564 (.A1(N3127), .A2(N3128), .ZN(N14436));
    NANDX1 U1565 (.A1(N3129), .A2(N3130), .ZN(n14437));
    NANDX1 U1566 (.A1(N3131), .A2(N3132), .ZN(n14438));
    NOR2X1 U1567 (.A1(N3133), .A2(N3134), .ZN(n14439));
    NOR2X1 U1568 (.A1(N3135), .A2(N3136), .ZN(n14440));
    NOR2X1 U1569 (.A1(N3137), .A2(N3138), .ZN(N14441));
    NOR2X1 U1570 (.A1(N3139), .A2(N3140), .ZN(n14442));
    NANDX1 U1571 (.A1(N3141), .A2(N3142), .ZN(N14443));
    NANDX1 U1572 (.A1(N3143), .A2(N3144), .ZN(N14444));
    NOR2X1 U1573 (.A1(N3145), .A2(N3146), .ZN(n14445));
    NOR2X1 U1574 (.A1(N3147), .A2(N3148), .ZN(n14446));
    NANDX1 U1575 (.A1(N3149), .A2(N3150), .ZN(n14447));
    NOR2X1 U1576 (.A1(N3151), .A2(N3152), .ZN(n14448));
    NANDX1 U1577 (.A1(N3153), .A2(N3154), .ZN(n14449));
    NOR2X1 U1578 (.A1(N3155), .A2(N3156), .ZN(n14450));
    NOR2X1 U1579 (.A1(N3157), .A2(N3158), .ZN(n14451));
    NOR2X1 U1580 (.A1(N3159), .A2(N3160), .ZN(n14452));
    NOR2X1 U1581 (.A1(N3161), .A2(N3162), .ZN(N14453));
    NOR2X1 U1582 (.A1(N3163), .A2(N3164), .ZN(n14454));
    NOR2X1 U1583 (.A1(N3165), .A2(N3166), .ZN(N14455));
    NANDX1 U1584 (.A1(N3167), .A2(N3168), .ZN(n14456));
    NOR2X1 U1585 (.A1(N3169), .A2(N3170), .ZN(n14457));
    NANDX1 U1586 (.A1(N3171), .A2(N3172), .ZN(n14458));
    NOR2X1 U1587 (.A1(N3173), .A2(N3174), .ZN(n14459));
    NOR2X1 U1588 (.A1(N3175), .A2(N3176), .ZN(n14460));
    NOR2X1 U1589 (.A1(N3177), .A2(N3178), .ZN(n14461));
    NANDX1 U1590 (.A1(N3179), .A2(N3180), .ZN(N14462));
    NOR2X1 U1591 (.A1(N3181), .A2(N3182), .ZN(n14463));
    NANDX1 U1592 (.A1(N3183), .A2(N3184), .ZN(n14464));
    NOR2X1 U1593 (.A1(N3185), .A2(N3186), .ZN(n14465));
    NOR2X1 U1594 (.A1(N3187), .A2(N3188), .ZN(n14466));
    NOR2X1 U1595 (.A1(N3189), .A2(N3190), .ZN(n14467));
    NOR2X1 U1596 (.A1(N3191), .A2(N3192), .ZN(n14468));
    NANDX1 U1597 (.A1(N3193), .A2(N3194), .ZN(N14469));
    NOR2X1 U1598 (.A1(N3195), .A2(N3196), .ZN(n14470));
    NOR2X1 U1599 (.A1(N3197), .A2(N3198), .ZN(N14471));
    NANDX1 U1600 (.A1(N3199), .A2(N3200), .ZN(n14472));
    NOR2X1 U1601 (.A1(N3201), .A2(N3202), .ZN(n14473));
    NANDX1 U1602 (.A1(N3203), .A2(N3204), .ZN(n14474));
    NOR2X1 U1603 (.A1(N3205), .A2(N3206), .ZN(n14475));
    NOR2X1 U1604 (.A1(N3207), .A2(N3208), .ZN(n14476));
    NOR2X1 U1605 (.A1(N3209), .A2(N3210), .ZN(n14477));
    NOR2X1 U1606 (.A1(N3211), .A2(N3212), .ZN(n14478));
    NANDX1 U1607 (.A1(N3213), .A2(N3214), .ZN(n14479));
    NANDX1 U1608 (.A1(N3215), .A2(N3216), .ZN(N14480));
    NOR2X1 U1609 (.A1(N3217), .A2(N3218), .ZN(N14481));
    NANDX1 U1610 (.A1(N3219), .A2(N3220), .ZN(n14482));
    NANDX1 U1611 (.A1(N3221), .A2(N3222), .ZN(n14483));
    NANDX1 U1612 (.A1(N3223), .A2(N3224), .ZN(n14484));
    NANDX1 U1613 (.A1(N3225), .A2(N3226), .ZN(n14485));
    NANDX1 U1614 (.A1(N3227), .A2(N3228), .ZN(n14486));
    NOR2X1 U1615 (.A1(N3229), .A2(N3230), .ZN(n14487));
    NANDX1 U1616 (.A1(N3231), .A2(N3232), .ZN(n14488));
    NOR2X1 U1617 (.A1(N3233), .A2(N3234), .ZN(n14489));
    NOR2X1 U1618 (.A1(N3235), .A2(N3236), .ZN(N14490));
    NANDX1 U1619 (.A1(N3237), .A2(N3238), .ZN(n14491));
    NOR2X1 U1620 (.A1(N3239), .A2(N3240), .ZN(n14492));
    NANDX1 U1621 (.A1(N3241), .A2(N3242), .ZN(n14493));
    NANDX1 U1622 (.A1(N3243), .A2(N3244), .ZN(n14494));
    NOR2X1 U1623 (.A1(N3245), .A2(N3246), .ZN(n14495));
    NOR2X1 U1624 (.A1(N3247), .A2(N3248), .ZN(n14496));
    NANDX1 U1625 (.A1(N3249), .A2(N3250), .ZN(n14497));
    NOR2X1 U1626 (.A1(N3251), .A2(N3252), .ZN(n14498));
    NOR2X1 U1627 (.A1(N3253), .A2(N3254), .ZN(N14499));
    NOR2X1 U1628 (.A1(N3255), .A2(N3256), .ZN(n14500));
    NOR2X1 U1629 (.A1(N3257), .A2(N3258), .ZN(n14501));
    NOR2X1 U1630 (.A1(N3259), .A2(N3260), .ZN(N14502));
    NANDX1 U1631 (.A1(N3261), .A2(N3262), .ZN(n14503));
    NOR2X1 U1632 (.A1(N3263), .A2(N3264), .ZN(n14504));
    NANDX1 U1633 (.A1(N3265), .A2(N3266), .ZN(n14505));
    NOR2X1 U1634 (.A1(N3267), .A2(N3268), .ZN(n14506));
    NANDX1 U1635 (.A1(N3269), .A2(N3270), .ZN(N14507));
    NANDX1 U1636 (.A1(N3271), .A2(N3272), .ZN(n14508));
    NOR2X1 U1637 (.A1(N3273), .A2(N3274), .ZN(n14509));
    NOR2X1 U1638 (.A1(N3275), .A2(N3276), .ZN(n14510));
    NOR2X1 U1639 (.A1(N3277), .A2(N3278), .ZN(n14511));
    NOR2X1 U1640 (.A1(N3279), .A2(N3280), .ZN(n14512));
    NANDX1 U1641 (.A1(N3281), .A2(N3282), .ZN(n14513));
    NANDX1 U1642 (.A1(N3283), .A2(N3284), .ZN(n14514));
    NANDX1 U1643 (.A1(N3285), .A2(N3286), .ZN(N14515));
    NOR2X1 U1644 (.A1(N3287), .A2(N3288), .ZN(n14516));
    NOR2X1 U1645 (.A1(N3289), .A2(N3290), .ZN(n14517));
    NANDX1 U1646 (.A1(N3291), .A2(N3292), .ZN(N14518));
    NANDX1 U1647 (.A1(N3293), .A2(N3294), .ZN(N14519));
    NOR2X1 U1648 (.A1(N3295), .A2(N3296), .ZN(n14520));
    NOR2X1 U1649 (.A1(N3297), .A2(N3298), .ZN(n14521));
    NOR2X1 U1650 (.A1(N3299), .A2(N3300), .ZN(n14522));
    NANDX1 U1651 (.A1(N3301), .A2(N3302), .ZN(n14523));
    NANDX1 U1652 (.A1(N3303), .A2(N3304), .ZN(n14524));
    NOR2X1 U1653 (.A1(N3305), .A2(N3306), .ZN(n14525));
    NANDX1 U1654 (.A1(N3307), .A2(N3308), .ZN(n14526));
    NANDX1 U1655 (.A1(N3309), .A2(N3310), .ZN(n14527));
    NANDX1 U1656 (.A1(N3311), .A2(N3312), .ZN(N14528));
    NANDX1 U1657 (.A1(N3313), .A2(N3314), .ZN(n14529));
    NANDX1 U1658 (.A1(N3315), .A2(N3316), .ZN(n14530));
    NOR2X1 U1659 (.A1(N3317), .A2(N3318), .ZN(n14531));
    NANDX1 U1660 (.A1(N3319), .A2(N3320), .ZN(n14532));
    NANDX1 U1661 (.A1(N3321), .A2(N3322), .ZN(n14533));
    NANDX1 U1662 (.A1(N3323), .A2(N3324), .ZN(n14534));
    NANDX1 U1663 (.A1(N3325), .A2(N3326), .ZN(n14535));
    NANDX1 U1664 (.A1(N3327), .A2(N3328), .ZN(n14536));
    NANDX1 U1665 (.A1(N3329), .A2(N3330), .ZN(n14537));
    NOR2X1 U1666 (.A1(N3331), .A2(N3332), .ZN(n14538));
    NOR2X1 U1667 (.A1(N3333), .A2(N3334), .ZN(n14539));
    NANDX1 U1668 (.A1(N3335), .A2(N3336), .ZN(n14540));
    NOR2X1 U1669 (.A1(N3337), .A2(N3338), .ZN(n14541));
    NANDX1 U1670 (.A1(N3339), .A2(N3340), .ZN(n14542));
    NOR2X1 U1671 (.A1(N3341), .A2(N3342), .ZN(n14543));
    NANDX1 U1672 (.A1(N3343), .A2(N3344), .ZN(n14544));
    NOR2X1 U1673 (.A1(N3345), .A2(N3346), .ZN(n14545));
    NANDX1 U1674 (.A1(N3347), .A2(N3348), .ZN(N14546));
    NANDX1 U1675 (.A1(N3349), .A2(N3350), .ZN(n14547));
    NANDX1 U1676 (.A1(N3351), .A2(N3352), .ZN(n14548));
    NANDX1 U1677 (.A1(N3353), .A2(N3354), .ZN(n14549));
    NOR2X1 U1678 (.A1(N3355), .A2(N3356), .ZN(n14550));
    NANDX1 U1679 (.A1(N3357), .A2(N3358), .ZN(n14551));
    NANDX1 U1680 (.A1(N3359), .A2(N3360), .ZN(n14552));
    NANDX1 U1681 (.A1(N3361), .A2(N3362), .ZN(N14553));
    NOR2X1 U1682 (.A1(N3363), .A2(N3364), .ZN(n14554));
    NOR2X1 U1683 (.A1(N3365), .A2(N3366), .ZN(n14555));
    NANDX1 U1684 (.A1(N3367), .A2(N3368), .ZN(n14556));
    NANDX1 U1685 (.A1(N3369), .A2(N3370), .ZN(n14557));
    NOR2X1 U1686 (.A1(N3371), .A2(N3372), .ZN(n14558));
    NOR2X1 U1687 (.A1(N3373), .A2(N3374), .ZN(n14559));
    NOR2X1 U1688 (.A1(N3375), .A2(N3376), .ZN(n14560));
    NANDX1 U1689 (.A1(N3377), .A2(N3378), .ZN(n14561));
    NOR2X1 U1690 (.A1(N3379), .A2(N3380), .ZN(n14562));
    NANDX1 U1691 (.A1(N3381), .A2(N3382), .ZN(N14563));
    NANDX1 U1692 (.A1(N3383), .A2(N3384), .ZN(n14564));
    NOR2X1 U1693 (.A1(N3385), .A2(N3386), .ZN(n14565));
    NANDX1 U1694 (.A1(N3387), .A2(N3388), .ZN(n14566));
    NOR2X1 U1695 (.A1(N3389), .A2(N3390), .ZN(n14567));
    NANDX1 U1696 (.A1(N3391), .A2(N3392), .ZN(N14568));
    NANDX1 U1697 (.A1(N3393), .A2(N3394), .ZN(n14569));
    NOR2X1 U1698 (.A1(N3395), .A2(N3396), .ZN(N14570));
    NANDX1 U1699 (.A1(N3397), .A2(N3398), .ZN(n14571));
    NOR2X1 U1700 (.A1(N3399), .A2(N3400), .ZN(n14572));
    NANDX1 U1701 (.A1(N3401), .A2(N3402), .ZN(n14573));
    NANDX1 U1702 (.A1(N3403), .A2(N3404), .ZN(n14574));
    NANDX1 U1703 (.A1(N3405), .A2(N3406), .ZN(n14575));
    NOR2X1 U1704 (.A1(N3407), .A2(N3408), .ZN(n14576));
    NOR2X1 U1705 (.A1(N3409), .A2(N3410), .ZN(N14577));
    NANDX1 U1706 (.A1(N3411), .A2(N3412), .ZN(N14578));
    NANDX1 U1707 (.A1(N3413), .A2(N3414), .ZN(n14579));
    NANDX1 U1708 (.A1(N3415), .A2(N3416), .ZN(n14580));
    NANDX1 U1709 (.A1(N3417), .A2(N3418), .ZN(n14581));
    NOR2X1 U1710 (.A1(N3419), .A2(N3420), .ZN(n14582));
    NOR2X1 U1711 (.A1(N3421), .A2(N3422), .ZN(n14583));
    NOR2X1 U1712 (.A1(N3423), .A2(N3424), .ZN(n14584));
    NANDX1 U1713 (.A1(N3425), .A2(N3426), .ZN(n14585));
    NANDX1 U1714 (.A1(N3427), .A2(N3428), .ZN(n14586));
    NANDX1 U1715 (.A1(N3429), .A2(N3430), .ZN(n14587));
    NOR2X1 U1716 (.A1(N3431), .A2(N3432), .ZN(n14588));
    NANDX1 U1717 (.A1(N3433), .A2(N3434), .ZN(n14589));
    NOR2X1 U1718 (.A1(N3435), .A2(N3436), .ZN(n14590));
    NANDX1 U1719 (.A1(N3437), .A2(N3438), .ZN(n14591));
    NOR2X1 U1720 (.A1(N3439), .A2(N3440), .ZN(n14592));
    NOR2X1 U1721 (.A1(N3441), .A2(N3442), .ZN(n14593));
    NOR2X1 U1722 (.A1(N3443), .A2(N3444), .ZN(N14594));
    NANDX1 U1723 (.A1(N3445), .A2(N3446), .ZN(n14595));
    NOR2X1 U1724 (.A1(N3447), .A2(N3448), .ZN(n14596));
    NANDX1 U1725 (.A1(N3449), .A2(N3450), .ZN(n14597));
    NANDX1 U1726 (.A1(N3451), .A2(N3452), .ZN(n14598));
    NOR2X1 U1727 (.A1(N3453), .A2(N3454), .ZN(n14599));
    NANDX1 U1728 (.A1(N3455), .A2(N3456), .ZN(N14600));
    NOR2X1 U1729 (.A1(N3457), .A2(N3458), .ZN(n14601));
    NANDX1 U1730 (.A1(N3459), .A2(N3460), .ZN(n14602));
    NANDX1 U1731 (.A1(N3461), .A2(N3462), .ZN(N14603));
    NANDX1 U1732 (.A1(N3463), .A2(N3464), .ZN(N14604));
    NOR2X1 U1733 (.A1(N3465), .A2(N3466), .ZN(n14605));
    NOR2X1 U1734 (.A1(N3467), .A2(N3468), .ZN(N14606));
    NANDX1 U1735 (.A1(N3469), .A2(N3470), .ZN(n14607));
    NOR2X1 U1736 (.A1(N3471), .A2(N3472), .ZN(N14608));
    NANDX1 U1737 (.A1(N3473), .A2(N3474), .ZN(n14609));
    NOR2X1 U1738 (.A1(N3475), .A2(N3476), .ZN(n14610));
    NOR2X1 U1739 (.A1(N3477), .A2(N3478), .ZN(n14611));
    NANDX1 U1740 (.A1(N3479), .A2(N3480), .ZN(n14612));
    NANDX1 U1741 (.A1(N3481), .A2(N3482), .ZN(N14613));
    NOR2X1 U1742 (.A1(N3483), .A2(N3484), .ZN(n14614));
    NANDX1 U1743 (.A1(N3485), .A2(N3486), .ZN(n14615));
    NOR2X1 U1744 (.A1(N3487), .A2(N3488), .ZN(n14616));
    NANDX1 U1745 (.A1(N3489), .A2(N3490), .ZN(n14617));
    NANDX1 U1746 (.A1(N3491), .A2(N3492), .ZN(n14618));
    NOR2X1 U1747 (.A1(N3493), .A2(N3494), .ZN(n14619));
    NOR2X1 U1748 (.A1(N3495), .A2(N3496), .ZN(n14620));
    NANDX1 U1749 (.A1(N3497), .A2(N3498), .ZN(n14621));
    NANDX1 U1750 (.A1(N3499), .A2(N3500), .ZN(n14622));
    NANDX1 U1751 (.A1(N3501), .A2(N3502), .ZN(N14623));
    NANDX1 U1752 (.A1(N3503), .A2(N3504), .ZN(n14624));
    NOR2X1 U1753 (.A1(N3505), .A2(N3506), .ZN(n14625));
    NOR2X1 U1754 (.A1(N3507), .A2(N3508), .ZN(n14626));
    NOR2X1 U1755 (.A1(N3509), .A2(N3510), .ZN(n14627));
    NANDX1 U1756 (.A1(N3511), .A2(N3512), .ZN(n14628));
    NOR2X1 U1757 (.A1(N3513), .A2(N3514), .ZN(n14629));
    NOR2X1 U1758 (.A1(N3515), .A2(N3516), .ZN(n14630));
    NOR2X1 U1759 (.A1(N3517), .A2(N3518), .ZN(n14631));
    NOR2X1 U1760 (.A1(N3519), .A2(N3520), .ZN(n14632));
    NANDX1 U1761 (.A1(N3521), .A2(N3522), .ZN(n14633));
    NANDX1 U1762 (.A1(N3523), .A2(N3524), .ZN(n14634));
    NANDX1 U1763 (.A1(N3525), .A2(N3526), .ZN(n14635));
    NANDX1 U1764 (.A1(N3527), .A2(N3528), .ZN(n14636));
    NOR2X1 U1765 (.A1(N3529), .A2(N3530), .ZN(N14637));
    NANDX1 U1766 (.A1(N3531), .A2(N3532), .ZN(N14638));
    NANDX1 U1767 (.A1(N3533), .A2(N3534), .ZN(n14639));
    NANDX1 U1768 (.A1(N3535), .A2(N3536), .ZN(n14640));
    NANDX1 U1769 (.A1(N3537), .A2(N3538), .ZN(n14641));
    NANDX1 U1770 (.A1(N3539), .A2(N3540), .ZN(n14642));
    NOR2X1 U1771 (.A1(N3541), .A2(N3542), .ZN(n14643));
    NOR2X1 U1772 (.A1(N3543), .A2(N3544), .ZN(n14644));
    NOR2X1 U1773 (.A1(N3545), .A2(N3546), .ZN(n14645));
    NOR2X1 U1774 (.A1(N3547), .A2(N3548), .ZN(n14646));
    NOR2X1 U1775 (.A1(N3549), .A2(N3550), .ZN(n14647));
    NANDX1 U1776 (.A1(N3551), .A2(N3552), .ZN(n14648));
    NANDX1 U1777 (.A1(N3553), .A2(N3554), .ZN(n14649));
    NANDX1 U1778 (.A1(N3555), .A2(N3556), .ZN(n14650));
    NOR2X1 U1779 (.A1(N3557), .A2(N3558), .ZN(n14651));
    NOR2X1 U1780 (.A1(N3559), .A2(N3560), .ZN(n14652));
    NOR2X1 U1781 (.A1(N3561), .A2(N3562), .ZN(N14653));
    NANDX1 U1782 (.A1(N3563), .A2(N3564), .ZN(n14654));
    NANDX1 U1783 (.A1(N3565), .A2(N3566), .ZN(n14655));
    NOR2X1 U1784 (.A1(N3567), .A2(N3568), .ZN(n14656));
    NANDX1 U1785 (.A1(N3569), .A2(N3570), .ZN(n14657));
    NANDX1 U1786 (.A1(N3571), .A2(N3572), .ZN(n14658));
    NOR2X1 U1787 (.A1(N3573), .A2(N3574), .ZN(n14659));
    NANDX1 U1788 (.A1(N3575), .A2(N3576), .ZN(n14660));
    NANDX1 U1789 (.A1(N3577), .A2(N3578), .ZN(n14661));
    NOR2X1 U1790 (.A1(N3579), .A2(N3580), .ZN(n14662));
    NANDX1 U1791 (.A1(N3581), .A2(N3582), .ZN(N14663));
    NOR2X1 U1792 (.A1(N3583), .A2(N3584), .ZN(n14664));
    NOR2X1 U1793 (.A1(N3585), .A2(N3586), .ZN(n14665));
    NANDX1 U1794 (.A1(N3587), .A2(N3588), .ZN(N14666));
    NANDX1 U1795 (.A1(N3589), .A2(N3590), .ZN(n14667));
    NOR2X1 U1796 (.A1(N3591), .A2(N3592), .ZN(n14668));
    NOR2X1 U1797 (.A1(N3593), .A2(N3594), .ZN(n14669));
    NANDX1 U1798 (.A1(N3595), .A2(N3596), .ZN(n14670));
    NANDX1 U1799 (.A1(N3597), .A2(N3598), .ZN(N14671));
    NANDX1 U1800 (.A1(N3599), .A2(N3600), .ZN(n14672));
    NOR2X1 U1801 (.A1(N3601), .A2(N3602), .ZN(n14673));
    NOR2X1 U1802 (.A1(N3603), .A2(N3604), .ZN(n14674));
    NOR2X1 U1803 (.A1(N3605), .A2(N3606), .ZN(n14675));
    NOR2X1 U1804 (.A1(N3607), .A2(N3608), .ZN(n14676));
    NOR2X1 U1805 (.A1(N3609), .A2(N3610), .ZN(n14677));
    NOR2X1 U1806 (.A1(N3611), .A2(N3612), .ZN(n14678));
    NOR2X1 U1807 (.A1(N3613), .A2(N3614), .ZN(N14679));
    NANDX1 U1808 (.A1(N3615), .A2(N3616), .ZN(N14680));
    NANDX1 U1809 (.A1(N3617), .A2(N3618), .ZN(n14681));
    NOR2X1 U1810 (.A1(N3619), .A2(N3620), .ZN(n14682));
    NANDX1 U1811 (.A1(N3621), .A2(N3622), .ZN(n14683));
    NOR2X1 U1812 (.A1(N3623), .A2(N3624), .ZN(n14684));
    NANDX1 U1813 (.A1(N3625), .A2(N3626), .ZN(N14685));
    NOR2X1 U1814 (.A1(N3627), .A2(N3628), .ZN(n14686));
    NOR2X1 U1815 (.A1(N3629), .A2(N3630), .ZN(n14687));
    NOR2X1 U1816 (.A1(N3631), .A2(N3632), .ZN(n14688));
    NOR2X1 U1817 (.A1(N3633), .A2(N3634), .ZN(n14689));
    NOR2X1 U1818 (.A1(N3635), .A2(N3636), .ZN(n14690));
    NOR2X1 U1819 (.A1(N3637), .A2(N3638), .ZN(N14691));
    NANDX1 U1820 (.A1(N3639), .A2(N3640), .ZN(n14692));
    NANDX1 U1821 (.A1(N3641), .A2(N3642), .ZN(n14693));
    NANDX1 U1822 (.A1(N3643), .A2(N3644), .ZN(N14694));
    NOR2X1 U1823 (.A1(N3645), .A2(N3646), .ZN(n14695));
    NANDX1 U1824 (.A1(N3647), .A2(N3648), .ZN(n14696));
    NOR2X1 U1825 (.A1(N3649), .A2(N3650), .ZN(n14697));
    NANDX1 U1826 (.A1(N3651), .A2(N3652), .ZN(N14698));
    NANDX1 U1827 (.A1(N3653), .A2(N3654), .ZN(n14699));
    NOR2X1 U1828 (.A1(N3655), .A2(N3656), .ZN(n14700));
    NOR2X1 U1829 (.A1(N3657), .A2(N3658), .ZN(n14701));
    NOR2X1 U1830 (.A1(N3659), .A2(N3660), .ZN(n14702));
    NOR2X1 U1831 (.A1(N3661), .A2(N3662), .ZN(n14703));
    NANDX1 U1832 (.A1(N3663), .A2(N3664), .ZN(n14704));
    NOR2X1 U1833 (.A1(N3665), .A2(N3666), .ZN(n14705));
    NOR2X1 U1834 (.A1(N3667), .A2(N3668), .ZN(n14706));
    NANDX1 U1835 (.A1(N3669), .A2(N3670), .ZN(n14707));
    NOR2X1 U1836 (.A1(N3671), .A2(N3672), .ZN(n14708));
    NOR2X1 U1837 (.A1(N3673), .A2(N3674), .ZN(N14709));
    NANDX1 U1838 (.A1(N3675), .A2(N3676), .ZN(n14710));
    NANDX1 U1839 (.A1(N3677), .A2(N3678), .ZN(n14711));
    NOR2X1 U1840 (.A1(N3679), .A2(N3680), .ZN(n14712));
    NANDX1 U1841 (.A1(N3681), .A2(N3682), .ZN(n14713));
    NOR2X1 U1842 (.A1(N3683), .A2(N3684), .ZN(n14714));
    NOR2X1 U1843 (.A1(N3685), .A2(N3686), .ZN(N14715));
    NOR2X1 U1844 (.A1(N3687), .A2(N3688), .ZN(n14716));
    NANDX1 U1845 (.A1(N3689), .A2(N3690), .ZN(n14717));
    NOR2X1 U1846 (.A1(N3691), .A2(N3692), .ZN(n14718));
    NANDX1 U1847 (.A1(N3693), .A2(N3694), .ZN(n14719));
    NANDX1 U1848 (.A1(N3695), .A2(N3696), .ZN(n14720));
    NANDX1 U1849 (.A1(N3697), .A2(N3698), .ZN(n14721));
    NANDX1 U1850 (.A1(N3699), .A2(N3700), .ZN(n14722));
    NOR2X1 U1851 (.A1(N3701), .A2(N3702), .ZN(n14723));
    NOR2X1 U1852 (.A1(N3703), .A2(N3704), .ZN(n14724));
    NOR2X1 U1853 (.A1(N3705), .A2(N3706), .ZN(N14725));
    NOR2X1 U1854 (.A1(N3707), .A2(N3708), .ZN(n14726));
    NANDX1 U1855 (.A1(N3709), .A2(N3710), .ZN(n14727));
    NANDX1 U1856 (.A1(N3711), .A2(N3712), .ZN(n14728));
    NOR2X1 U1857 (.A1(N3713), .A2(N3714), .ZN(n14729));
    NOR2X1 U1858 (.A1(N3715), .A2(N3716), .ZN(n14730));
    NANDX1 U1859 (.A1(N3717), .A2(N3718), .ZN(n14731));
    NOR2X1 U1860 (.A1(N3719), .A2(N3720), .ZN(n14732));
    NOR2X1 U1861 (.A1(N3721), .A2(N3722), .ZN(N14733));
    NANDX1 U1862 (.A1(N3723), .A2(N3724), .ZN(n14734));
    NANDX1 U1863 (.A1(N3725), .A2(N3726), .ZN(n14735));
    NANDX1 U1864 (.A1(N3727), .A2(N3728), .ZN(N14736));
    NANDX1 U1865 (.A1(N3729), .A2(N3730), .ZN(n14737));
    NANDX1 U1866 (.A1(N3731), .A2(N3732), .ZN(n14738));
    NANDX1 U1867 (.A1(N3733), .A2(N3734), .ZN(n14739));
    NOR2X1 U1868 (.A1(N3735), .A2(N3736), .ZN(n14740));
    NOR2X1 U1869 (.A1(N3737), .A2(N3738), .ZN(n14741));
    NANDX1 U1870 (.A1(N3739), .A2(N3740), .ZN(n14742));
    NOR2X1 U1871 (.A1(N3741), .A2(N3742), .ZN(n14743));
    NOR2X1 U1872 (.A1(N3743), .A2(N3744), .ZN(N14744));
    NANDX1 U1873 (.A1(N3745), .A2(N3746), .ZN(n14745));
    NOR2X1 U1874 (.A1(N3747), .A2(N3748), .ZN(n14746));
    NOR2X1 U1875 (.A1(N3749), .A2(N3750), .ZN(n14747));
    NOR2X1 U1876 (.A1(N3751), .A2(N3752), .ZN(n14748));
    NOR2X1 U1877 (.A1(N3753), .A2(N3754), .ZN(n14749));
    NANDX1 U1878 (.A1(N3755), .A2(N3756), .ZN(n14750));
    NANDX1 U1879 (.A1(N3757), .A2(N3758), .ZN(n14751));
    NANDX1 U1880 (.A1(N3759), .A2(N3760), .ZN(N14752));
    NOR2X1 U1881 (.A1(N3761), .A2(N3762), .ZN(n14753));
    NOR2X1 U1882 (.A1(N3763), .A2(N3764), .ZN(n14754));
    NANDX1 U1883 (.A1(N3765), .A2(N3766), .ZN(N14755));
    NANDX1 U1884 (.A1(N3767), .A2(N3768), .ZN(N14756));
    NOR2X1 U1885 (.A1(N3769), .A2(N3770), .ZN(n14757));
    NOR2X1 U1886 (.A1(N3771), .A2(N3772), .ZN(n14758));
    NOR2X1 U1887 (.A1(N3773), .A2(N3774), .ZN(n14759));
    NOR2X1 U1888 (.A1(N3775), .A2(N3776), .ZN(n14760));
    NOR2X1 U1889 (.A1(N3777), .A2(N3778), .ZN(n14761));
    NANDX1 U1890 (.A1(N3779), .A2(N3780), .ZN(n14762));
    NANDX1 U1891 (.A1(N3781), .A2(N3782), .ZN(n14763));
    NANDX1 U1892 (.A1(N3783), .A2(N3784), .ZN(n14764));
    NANDX1 U1893 (.A1(N3785), .A2(N3786), .ZN(n14765));
    NOR2X1 U1894 (.A1(N3787), .A2(N3788), .ZN(n14766));
    NOR2X1 U1895 (.A1(N3789), .A2(N3790), .ZN(N14767));
    NOR2X1 U1896 (.A1(N3791), .A2(N3792), .ZN(n14768));
    NANDX1 U1897 (.A1(N3793), .A2(N3794), .ZN(n14769));
    NANDX1 U1898 (.A1(N3795), .A2(N3796), .ZN(n14770));
    NOR2X1 U1899 (.A1(N3797), .A2(N3798), .ZN(n14771));
    NOR2X1 U1900 (.A1(N3799), .A2(N3800), .ZN(n14772));
    NOR2X1 U1901 (.A1(N3801), .A2(N3802), .ZN(n14773));
    NOR2X1 U1902 (.A1(N3803), .A2(N3804), .ZN(n14774));
    NOR2X1 U1903 (.A1(N3805), .A2(N3806), .ZN(N14775));
    NOR2X1 U1904 (.A1(N3807), .A2(N3808), .ZN(n14776));
    NOR2X1 U1905 (.A1(N3809), .A2(N3810), .ZN(n14777));
    NOR2X1 U1906 (.A1(N3811), .A2(N3812), .ZN(n14778));
    NOR2X1 U1907 (.A1(N3813), .A2(N3814), .ZN(n14779));
    NANDX1 U1908 (.A1(N3815), .A2(N3816), .ZN(n14780));
    NOR2X1 U1909 (.A1(N3817), .A2(N3818), .ZN(n14781));
    NOR2X1 U1910 (.A1(N3819), .A2(N3820), .ZN(n14782));
    NOR2X1 U1911 (.A1(N3821), .A2(N3822), .ZN(N14783));
    NOR2X1 U1912 (.A1(N3823), .A2(N3824), .ZN(n14784));
    NOR2X1 U1913 (.A1(N3825), .A2(N3826), .ZN(N14785));
    NOR2X1 U1914 (.A1(N3827), .A2(N3828), .ZN(n14786));
    NANDX1 U1915 (.A1(N3829), .A2(N3830), .ZN(n14787));
    NOR2X1 U1916 (.A1(N3831), .A2(N3832), .ZN(n14788));
    NOR2X1 U1917 (.A1(N3833), .A2(N3834), .ZN(n14789));
    NANDX1 U1918 (.A1(N3835), .A2(N3836), .ZN(n14790));
    NANDX1 U1919 (.A1(N3837), .A2(N3838), .ZN(N14791));
    NANDX1 U1920 (.A1(N3839), .A2(N3840), .ZN(n14792));
    NANDX1 U1921 (.A1(N3841), .A2(N3842), .ZN(n14793));
    NOR2X1 U1922 (.A1(N3843), .A2(N3844), .ZN(n14794));
    NOR2X1 U1923 (.A1(N3845), .A2(N3846), .ZN(n14795));
    NOR2X1 U1924 (.A1(N3847), .A2(N3848), .ZN(n14796));
    NOR2X1 U1925 (.A1(N3849), .A2(N3850), .ZN(n14797));
    NOR2X1 U1926 (.A1(N3851), .A2(N3852), .ZN(n14798));
    NOR2X1 U1927 (.A1(N3853), .A2(N3854), .ZN(n14799));
    NOR2X1 U1928 (.A1(N3855), .A2(N3856), .ZN(n14800));
    NANDX1 U1929 (.A1(N3857), .A2(N3858), .ZN(n14801));
    NANDX1 U1930 (.A1(N3859), .A2(N3860), .ZN(n14802));
    NOR2X1 U1931 (.A1(N3861), .A2(N3862), .ZN(n14803));
    NOR2X1 U1932 (.A1(N3863), .A2(N3864), .ZN(n14804));
    NANDX1 U1933 (.A1(N3865), .A2(N3866), .ZN(n14805));
    NOR2X1 U1934 (.A1(N3867), .A2(N3868), .ZN(n14806));
    NOR2X1 U1935 (.A1(N3869), .A2(N3870), .ZN(n14807));
    NOR2X1 U1936 (.A1(N3871), .A2(N3872), .ZN(n14808));
    NOR2X1 U1937 (.A1(N3873), .A2(N3874), .ZN(n14809));
    NOR2X1 U1938 (.A1(N3875), .A2(N3876), .ZN(n14810));
    NANDX1 U1939 (.A1(N3877), .A2(N3878), .ZN(n14811));
    NOR2X1 U1940 (.A1(N3879), .A2(N3880), .ZN(N14812));
    NOR2X1 U1941 (.A1(N3881), .A2(N3882), .ZN(n14813));
    NANDX1 U1942 (.A1(N3883), .A2(N3884), .ZN(n14814));
    NANDX1 U1943 (.A1(N3885), .A2(N3886), .ZN(n14815));
    NOR2X1 U1944 (.A1(N3887), .A2(N3888), .ZN(n14816));
    NANDX1 U1945 (.A1(N3889), .A2(N3890), .ZN(n14817));
    NOR2X1 U1946 (.A1(N3891), .A2(N3892), .ZN(n14818));
    NANDX1 U1947 (.A1(N3893), .A2(N3894), .ZN(n14819));
    NOR2X1 U1948 (.A1(N3895), .A2(N3896), .ZN(n14820));
    NOR2X1 U1949 (.A1(N3897), .A2(N3898), .ZN(n14821));
    NOR2X1 U1950 (.A1(N3899), .A2(N3900), .ZN(n14822));
    NANDX1 U1951 (.A1(N3901), .A2(N3902), .ZN(n14823));
    NANDX1 U1952 (.A1(N3903), .A2(N3904), .ZN(N14824));
    NOR2X1 U1953 (.A1(N3905), .A2(N3906), .ZN(n14825));
    NANDX1 U1954 (.A1(N3907), .A2(N3908), .ZN(N14826));
    NANDX1 U1955 (.A1(N3909), .A2(N3910), .ZN(n14827));
    NOR2X1 U1956 (.A1(N3911), .A2(N3912), .ZN(n14828));
    NANDX1 U1957 (.A1(N3913), .A2(N3914), .ZN(n14829));
    NANDX1 U1958 (.A1(N3915), .A2(N3916), .ZN(n14830));
    NOR2X1 U1959 (.A1(N3917), .A2(N3918), .ZN(N14831));
    NOR2X1 U1960 (.A1(N3919), .A2(N3920), .ZN(n14832));
    NOR2X1 U1961 (.A1(N3921), .A2(N3922), .ZN(n14833));
    NOR2X1 U1962 (.A1(N3923), .A2(N3924), .ZN(n14834));
    NOR2X1 U1963 (.A1(N3925), .A2(N3926), .ZN(n14835));
    NOR2X1 U1964 (.A1(N3927), .A2(N3928), .ZN(n14836));
    NOR2X1 U1965 (.A1(N3929), .A2(N3930), .ZN(N14837));
    NOR2X1 U1966 (.A1(N3931), .A2(N3932), .ZN(n14838));
    NOR2X1 U1967 (.A1(N3933), .A2(N3934), .ZN(N14839));
    NANDX1 U1968 (.A1(N3935), .A2(N3936), .ZN(N14840));
    NANDX1 U1969 (.A1(N3937), .A2(N3938), .ZN(n14841));
    NANDX1 U1970 (.A1(N3939), .A2(N3940), .ZN(n14842));
    NANDX1 U1971 (.A1(N3941), .A2(N3942), .ZN(n14843));
    NANDX1 U1972 (.A1(N3943), .A2(N3944), .ZN(n14844));
    NOR2X1 U1973 (.A1(N3945), .A2(N3946), .ZN(n14845));
    NOR2X1 U1974 (.A1(N3947), .A2(N3948), .ZN(n14846));
    NOR2X1 U1975 (.A1(N3949), .A2(N3950), .ZN(n14847));
    NOR2X1 U1976 (.A1(N3951), .A2(N3952), .ZN(N14848));
    NANDX1 U1977 (.A1(N3953), .A2(N3954), .ZN(N14849));
    NANDX1 U1978 (.A1(N3955), .A2(N3956), .ZN(N14850));
    NOR2X1 U1979 (.A1(N3957), .A2(N3958), .ZN(n14851));
    NANDX1 U1980 (.A1(N3959), .A2(N3960), .ZN(n14852));
    NANDX1 U1981 (.A1(N3961), .A2(N3962), .ZN(n14853));
    NANDX1 U1982 (.A1(N3963), .A2(N3964), .ZN(n14854));
    NOR2X1 U1983 (.A1(N3965), .A2(N3966), .ZN(n14855));
    NANDX1 U1984 (.A1(N3967), .A2(N3968), .ZN(n14856));
    NOR2X1 U1985 (.A1(N3969), .A2(N3970), .ZN(n14857));
    NANDX1 U1986 (.A1(N3971), .A2(N3972), .ZN(n14858));
    NANDX1 U1987 (.A1(N3973), .A2(N3974), .ZN(n14859));
    NANDX1 U1988 (.A1(N3975), .A2(N3976), .ZN(n14860));
    NOR2X1 U1989 (.A1(N3977), .A2(N3978), .ZN(n14861));
    NOR2X1 U1990 (.A1(N3979), .A2(N3980), .ZN(n14862));
    NANDX1 U1991 (.A1(N3981), .A2(N3982), .ZN(N14863));
    NANDX1 U1992 (.A1(N3983), .A2(N3984), .ZN(n14864));
    NOR2X1 U1993 (.A1(N3985), .A2(N3986), .ZN(n14865));
    NOR2X1 U1994 (.A1(N3987), .A2(N3988), .ZN(n14866));
    NANDX1 U1995 (.A1(N3989), .A2(N3990), .ZN(N14867));
    NANDX1 U1996 (.A1(N3991), .A2(N3992), .ZN(n14868));
    NOR2X1 U1997 (.A1(N3993), .A2(N3994), .ZN(n14869));
    NANDX1 U1998 (.A1(N3995), .A2(N3996), .ZN(n14870));
    NOR2X1 U1999 (.A1(N3997), .A2(N3998), .ZN(n14871));
    NANDX1 U2000 (.A1(N3999), .A2(N4000), .ZN(n14872));
    NOR2X1 U2001 (.A1(N4001), .A2(N4002), .ZN(n14873));
    NANDX1 U2002 (.A1(N4003), .A2(N4004), .ZN(n14874));
    NANDX1 U2003 (.A1(N4005), .A2(N4006), .ZN(n14875));
    NOR2X1 U2004 (.A1(N4007), .A2(N4008), .ZN(N14876));
    NOR2X1 U2005 (.A1(N4009), .A2(N4010), .ZN(n14877));
    NANDX1 U2006 (.A1(N4011), .A2(N4012), .ZN(n14878));
    NOR2X1 U2007 (.A1(N4013), .A2(N4014), .ZN(n14879));
    NANDX1 U2008 (.A1(N4015), .A2(N4016), .ZN(n14880));
    NOR2X1 U2009 (.A1(N4017), .A2(N4018), .ZN(N14881));
    NOR2X1 U2010 (.A1(N4019), .A2(N4020), .ZN(n14882));
    NOR2X1 U2011 (.A1(N4021), .A2(N4022), .ZN(n14883));
    NANDX1 U2012 (.A1(N4023), .A2(N4024), .ZN(n14884));
    NANDX1 U2013 (.A1(N4025), .A2(N4026), .ZN(n14885));
    NOR2X1 U2014 (.A1(N4027), .A2(N4028), .ZN(n14886));
    NOR2X1 U2015 (.A1(N4029), .A2(N4030), .ZN(n14887));
    NANDX1 U2016 (.A1(N4031), .A2(N4032), .ZN(n14888));
    NANDX1 U2017 (.A1(N4033), .A2(N4034), .ZN(n14889));
    NANDX1 U2018 (.A1(N4035), .A2(N4036), .ZN(N14890));
    NOR2X1 U2019 (.A1(N4037), .A2(N4038), .ZN(n14891));
    NANDX1 U2020 (.A1(N4039), .A2(N4040), .ZN(n14892));
    NANDX1 U2021 (.A1(N4041), .A2(N4042), .ZN(n14893));
    NOR2X1 U2022 (.A1(N4043), .A2(N4044), .ZN(n14894));
    NOR2X1 U2023 (.A1(N4045), .A2(N4046), .ZN(n14895));
    NOR2X1 U2024 (.A1(N4047), .A2(N4048), .ZN(n14896));
    NOR2X1 U2025 (.A1(N4049), .A2(N4050), .ZN(n14897));
    NANDX1 U2026 (.A1(N4051), .A2(N4052), .ZN(N14898));
    NANDX1 U2027 (.A1(N4053), .A2(N4054), .ZN(N14899));
    NOR2X1 U2028 (.A1(N4055), .A2(N4056), .ZN(n14900));
    NOR2X1 U2029 (.A1(N4057), .A2(N4058), .ZN(n14901));
    NANDX1 U2030 (.A1(N4059), .A2(N4060), .ZN(n14902));
    NOR2X1 U2031 (.A1(N4061), .A2(N4062), .ZN(n14903));
    NOR2X1 U2032 (.A1(N4063), .A2(N4064), .ZN(n14904));
    NOR2X1 U2033 (.A1(N4065), .A2(N4066), .ZN(n14905));
    NANDX1 U2034 (.A1(N4067), .A2(N4068), .ZN(n14906));
    NANDX1 U2035 (.A1(N4069), .A2(N4070), .ZN(n14907));
    NOR2X1 U2036 (.A1(N4071), .A2(N4072), .ZN(n14908));
    NOR2X1 U2037 (.A1(N4073), .A2(N4074), .ZN(n14909));
    NANDX1 U2038 (.A1(N4075), .A2(N4076), .ZN(n14910));
    NANDX1 U2039 (.A1(N4077), .A2(N4078), .ZN(n14911));
    NOR2X1 U2040 (.A1(N4079), .A2(N4080), .ZN(n14912));
    NOR2X1 U2041 (.A1(N4081), .A2(N4082), .ZN(n14913));
    NANDX1 U2042 (.A1(N4083), .A2(N4084), .ZN(n14914));
    NANDX1 U2043 (.A1(N4085), .A2(N4086), .ZN(n14915));
    NANDX1 U2044 (.A1(N4087), .A2(N4088), .ZN(n14916));
    NANDX1 U2045 (.A1(N4089), .A2(N4090), .ZN(n14917));
    NANDX1 U2046 (.A1(N4091), .A2(N4092), .ZN(n14918));
    NANDX1 U2047 (.A1(N4093), .A2(N4094), .ZN(n14919));
    NOR2X1 U2048 (.A1(N4095), .A2(N4096), .ZN(N14920));
    NOR2X1 U2049 (.A1(N4097), .A2(N4098), .ZN(n14921));
    NANDX1 U2050 (.A1(N4099), .A2(N4100), .ZN(N14922));
    NOR2X1 U2051 (.A1(N4101), .A2(N4102), .ZN(n14923));
    NOR2X1 U2052 (.A1(N4103), .A2(N4104), .ZN(n14924));
    NANDX1 U2053 (.A1(N4105), .A2(N4106), .ZN(n14925));
    NOR2X1 U2054 (.A1(N4107), .A2(N4108), .ZN(n14926));
    NOR2X1 U2055 (.A1(N4109), .A2(N4110), .ZN(n14927));
    NANDX1 U2056 (.A1(N4111), .A2(N4112), .ZN(n14928));
    NOR2X1 U2057 (.A1(N4113), .A2(N4114), .ZN(n14929));
    NANDX1 U2058 (.A1(N4115), .A2(N4116), .ZN(n14930));
    NOR2X1 U2059 (.A1(N4117), .A2(N4118), .ZN(N14931));
    NOR2X1 U2060 (.A1(N4119), .A2(N4120), .ZN(n14932));
    NOR2X1 U2061 (.A1(N4121), .A2(N4122), .ZN(n14933));
    NOR2X1 U2062 (.A1(N4123), .A2(N4124), .ZN(n14934));
    NANDX1 U2063 (.A1(N4125), .A2(N4126), .ZN(n14935));
    NOR2X1 U2064 (.A1(N4127), .A2(N4128), .ZN(N14936));
    NANDX1 U2065 (.A1(N4129), .A2(N4130), .ZN(n14937));
    NOR2X1 U2066 (.A1(N4131), .A2(N4132), .ZN(n14938));
    NANDX1 U2067 (.A1(N4133), .A2(N4134), .ZN(N14939));
    NANDX1 U2068 (.A1(N4135), .A2(N4136), .ZN(n14940));
    NANDX1 U2069 (.A1(N4137), .A2(N4138), .ZN(n14941));
    NOR2X1 U2070 (.A1(N4139), .A2(N4140), .ZN(n14942));
    NANDX1 U2071 (.A1(N4141), .A2(N4142), .ZN(n14943));
    NANDX1 U2072 (.A1(N4143), .A2(N4144), .ZN(n14944));
    NOR2X1 U2073 (.A1(N4145), .A2(N4146), .ZN(n14945));
    NOR2X1 U2074 (.A1(N4147), .A2(N4148), .ZN(n14946));
    NANDX1 U2075 (.A1(N4149), .A2(N4150), .ZN(N14947));
    NANDX1 U2076 (.A1(N4151), .A2(N4152), .ZN(n14948));
    NANDX1 U2077 (.A1(N4153), .A2(N4154), .ZN(n14949));
    NOR2X1 U2078 (.A1(N4155), .A2(N4156), .ZN(n14950));
    NOR2X1 U2079 (.A1(N4157), .A2(N4158), .ZN(n14951));
    NANDX1 U2080 (.A1(N4159), .A2(N4160), .ZN(n14952));
    NANDX1 U2081 (.A1(N4161), .A2(N4162), .ZN(N14953));
    NOR2X1 U2082 (.A1(N4163), .A2(N4164), .ZN(n14954));
    NANDX1 U2083 (.A1(N4165), .A2(N4166), .ZN(n14955));
    NANDX1 U2084 (.A1(N4167), .A2(N4168), .ZN(n14956));
    NOR2X1 U2085 (.A1(N4169), .A2(N4170), .ZN(n14957));
    NANDX1 U2086 (.A1(N4171), .A2(N4172), .ZN(N14958));
    NOR2X1 U2087 (.A1(N4173), .A2(N4174), .ZN(n14959));
    NOR2X1 U2088 (.A1(N4175), .A2(N4176), .ZN(n14960));
    NOR2X1 U2089 (.A1(N4177), .A2(N4178), .ZN(N14961));
    NOR2X1 U2090 (.A1(N4179), .A2(N4180), .ZN(n14962));
    NANDX1 U2091 (.A1(N4181), .A2(N4182), .ZN(n14963));
    NOR2X1 U2092 (.A1(N4183), .A2(N4184), .ZN(n14964));
    NOR2X1 U2093 (.A1(N4185), .A2(N4186), .ZN(n14965));
    NOR2X1 U2094 (.A1(N4187), .A2(N4188), .ZN(n14966));
    NANDX1 U2095 (.A1(N4189), .A2(N4190), .ZN(n14967));
    NANDX1 U2096 (.A1(N4191), .A2(N4192), .ZN(N14968));
    NOR2X1 U2097 (.A1(N4193), .A2(N4194), .ZN(N14969));
    NOR2X1 U2098 (.A1(N4195), .A2(N4196), .ZN(n14970));
    NOR2X1 U2099 (.A1(N4197), .A2(N4198), .ZN(N14971));
    NANDX1 U2100 (.A1(N4199), .A2(N4200), .ZN(n14972));
    NOR2X1 U2101 (.A1(N4201), .A2(N4202), .ZN(n14973));
    NANDX1 U2102 (.A1(N4203), .A2(N4204), .ZN(n14974));
    NANDX1 U2103 (.A1(N4205), .A2(N4206), .ZN(n14975));
    NOR2X1 U2104 (.A1(N4207), .A2(N4208), .ZN(n14976));
    NANDX1 U2105 (.A1(N4209), .A2(N4210), .ZN(n14977));
    NOR2X1 U2106 (.A1(N4211), .A2(N4212), .ZN(N14978));
    NOR2X1 U2107 (.A1(N4213), .A2(N4214), .ZN(n14979));
    NOR2X1 U2108 (.A1(N4215), .A2(N4216), .ZN(n14980));
    NOR2X1 U2109 (.A1(N4217), .A2(N4218), .ZN(n14981));
    NOR2X1 U2110 (.A1(N4219), .A2(N4220), .ZN(n14982));
    NOR2X1 U2111 (.A1(N4221), .A2(N4222), .ZN(n14983));
    NANDX1 U2112 (.A1(N4223), .A2(N4224), .ZN(n14984));
    NOR2X1 U2113 (.A1(N4225), .A2(N4226), .ZN(n14985));
    NANDX1 U2114 (.A1(N4227), .A2(N4228), .ZN(n14986));
    NOR2X1 U2115 (.A1(N4229), .A2(N4230), .ZN(n14987));
    NOR2X1 U2116 (.A1(N4231), .A2(N4232), .ZN(n14988));
    NANDX1 U2117 (.A1(N4233), .A2(N4234), .ZN(n14989));
    NANDX1 U2118 (.A1(N4235), .A2(N4236), .ZN(n14990));
    NANDX1 U2119 (.A1(N4237), .A2(N4238), .ZN(N14991));
    NANDX1 U2120 (.A1(N4239), .A2(N4240), .ZN(N14992));
    NANDX1 U2121 (.A1(N4241), .A2(N4242), .ZN(n14993));
    NOR2X1 U2122 (.A1(N4243), .A2(N4244), .ZN(n14994));
    NOR2X1 U2123 (.A1(N4245), .A2(N4246), .ZN(n14995));
    NOR2X1 U2124 (.A1(N4247), .A2(N4248), .ZN(n14996));
    NOR2X1 U2125 (.A1(N4249), .A2(N4250), .ZN(n14997));
    NANDX1 U2126 (.A1(N4251), .A2(N4252), .ZN(n14998));
    NANDX1 U2127 (.A1(N4253), .A2(N4254), .ZN(n14999));
    NOR2X1 U2128 (.A1(N4255), .A2(N4256), .ZN(n15000));
    NANDX1 U2129 (.A1(N4257), .A2(N4258), .ZN(n15001));
    NOR2X1 U2130 (.A1(N4259), .A2(N4260), .ZN(N15002));
    NANDX1 U2131 (.A1(N4261), .A2(N4262), .ZN(n15003));
    NANDX1 U2132 (.A1(N4263), .A2(N4264), .ZN(n15004));
    NANDX1 U2133 (.A1(N4265), .A2(N4266), .ZN(N15005));
    NOR2X1 U2134 (.A1(N4267), .A2(N4268), .ZN(N15006));
    NOR2X1 U2135 (.A1(N4269), .A2(N4270), .ZN(n15007));
    NANDX1 U2136 (.A1(N4271), .A2(N4272), .ZN(n15008));
    NOR2X1 U2137 (.A1(N4273), .A2(N4274), .ZN(n15009));
    NOR2X1 U2138 (.A1(N4275), .A2(N4276), .ZN(n15010));
    NANDX1 U2139 (.A1(N4277), .A2(N4278), .ZN(n15011));
    NOR2X1 U2140 (.A1(N4279), .A2(N4280), .ZN(n15012));
    NOR2X1 U2141 (.A1(N4281), .A2(N4282), .ZN(N15013));
    NANDX1 U2142 (.A1(N4283), .A2(N4284), .ZN(n15014));
    NOR2X1 U2143 (.A1(N4285), .A2(N4286), .ZN(N15015));
    NOR2X1 U2144 (.A1(N4287), .A2(N4288), .ZN(n15016));
    NANDX1 U2145 (.A1(N4289), .A2(N4290), .ZN(n15017));
    NOR2X1 U2146 (.A1(N4291), .A2(N4292), .ZN(N15018));
    NOR2X1 U2147 (.A1(N4293), .A2(N4294), .ZN(n15019));
    NOR2X1 U2148 (.A1(N4295), .A2(N4296), .ZN(n15020));
    NANDX1 U2149 (.A1(N4297), .A2(N4298), .ZN(n15021));
    NANDX1 U2150 (.A1(N4299), .A2(N4300), .ZN(n15022));
    NANDX1 U2151 (.A1(N4301), .A2(N4302), .ZN(n15023));
    NANDX1 U2152 (.A1(N4303), .A2(N4304), .ZN(n15024));
    NANDX1 U2153 (.A1(N4305), .A2(N4306), .ZN(n15025));
    NANDX1 U2154 (.A1(N4307), .A2(N4308), .ZN(n15026));
    NANDX1 U2155 (.A1(N4309), .A2(N4310), .ZN(n15027));
    NANDX1 U2156 (.A1(N4311), .A2(N4312), .ZN(n15028));
    NOR2X1 U2157 (.A1(N4313), .A2(N4314), .ZN(n15029));
    NOR2X1 U2158 (.A1(N4315), .A2(N4316), .ZN(n15030));
    NANDX1 U2159 (.A1(N4317), .A2(N4318), .ZN(n15031));
    NANDX1 U2160 (.A1(N4319), .A2(N4320), .ZN(N15032));
    NOR2X1 U2161 (.A1(N4321), .A2(N4322), .ZN(n15033));
    NANDX1 U2162 (.A1(N4323), .A2(N4324), .ZN(n15034));
    NANDX1 U2163 (.A1(N4325), .A2(N4326), .ZN(N15035));
    NOR2X1 U2164 (.A1(N4327), .A2(N4328), .ZN(n15036));
    NANDX1 U2165 (.A1(N4329), .A2(N4330), .ZN(n15037));
    NANDX1 U2166 (.A1(N4331), .A2(N4332), .ZN(N15038));
    NANDX1 U2167 (.A1(N4333), .A2(N4334), .ZN(n15039));
    NOR2X1 U2168 (.A1(N4335), .A2(N4336), .ZN(n15040));
    NANDX1 U2169 (.A1(N4337), .A2(N4338), .ZN(n15041));
    NOR2X1 U2170 (.A1(N4339), .A2(N4340), .ZN(n15042));
    NOR2X1 U2171 (.A1(N4341), .A2(N4342), .ZN(n15043));
    NANDX1 U2172 (.A1(N4343), .A2(N4344), .ZN(n15044));
    NOR2X1 U2173 (.A1(N4345), .A2(N4346), .ZN(n15045));
    NOR2X1 U2174 (.A1(N4347), .A2(N4348), .ZN(n15046));
    NANDX1 U2175 (.A1(N4349), .A2(N4350), .ZN(n15047));
    NANDX1 U2176 (.A1(N4351), .A2(N4352), .ZN(n15048));
    NANDX1 U2177 (.A1(N4353), .A2(N4354), .ZN(n15049));
    NANDX1 U2178 (.A1(N4355), .A2(N4356), .ZN(n15050));
    NANDX1 U2179 (.A1(N4357), .A2(N4358), .ZN(n15051));
    NOR2X1 U2180 (.A1(N4359), .A2(N4360), .ZN(n15052));
    NANDX1 U2181 (.A1(N4361), .A2(N4362), .ZN(n15053));
    NOR2X1 U2182 (.A1(N4363), .A2(N4364), .ZN(n15054));
    NANDX1 U2183 (.A1(N4365), .A2(N4366), .ZN(n15055));
    NOR2X1 U2184 (.A1(N4367), .A2(N4368), .ZN(n15056));
    NOR2X1 U2185 (.A1(N4369), .A2(N4370), .ZN(n15057));
    NOR2X1 U2186 (.A1(N4371), .A2(N4372), .ZN(n15058));
    NOR2X1 U2187 (.A1(N4373), .A2(N4374), .ZN(n15059));
    NOR2X1 U2188 (.A1(N4375), .A2(N4376), .ZN(n15060));
    NANDX1 U2189 (.A1(N4377), .A2(N4378), .ZN(n15061));
    NANDX1 U2190 (.A1(N4379), .A2(N4380), .ZN(n15062));
    NOR2X1 U2191 (.A1(N4381), .A2(N4382), .ZN(n15063));
    NANDX1 U2192 (.A1(N4383), .A2(N4384), .ZN(n15064));
    NOR2X1 U2193 (.A1(N4385), .A2(N4386), .ZN(n15065));
    NANDX1 U2194 (.A1(N4387), .A2(N4388), .ZN(n15066));
    NANDX1 U2195 (.A1(N4389), .A2(N4390), .ZN(n15067));
    NOR2X1 U2196 (.A1(N4391), .A2(N4392), .ZN(n15068));
    NOR2X1 U2197 (.A1(N4393), .A2(N4394), .ZN(n15069));
    NOR2X1 U2198 (.A1(N4395), .A2(N4396), .ZN(n15070));
    NOR2X1 U2199 (.A1(N4397), .A2(N4398), .ZN(N15071));
    NANDX1 U2200 (.A1(N4399), .A2(N4400), .ZN(n15072));
    NANDX1 U2201 (.A1(N4401), .A2(N4402), .ZN(n15073));
    NOR2X1 U2202 (.A1(N4403), .A2(N4404), .ZN(n15074));
    NOR2X1 U2203 (.A1(N4405), .A2(N4406), .ZN(N15075));
    NANDX1 U2204 (.A1(N4407), .A2(N4408), .ZN(n15076));
    NANDX1 U2205 (.A1(N4409), .A2(N4410), .ZN(n15077));
    NANDX1 U2206 (.A1(N4411), .A2(N4412), .ZN(N15078));
    NOR2X1 U2207 (.A1(N4413), .A2(N4414), .ZN(n15079));
    NOR2X1 U2208 (.A1(N4415), .A2(N4416), .ZN(n15080));
    NOR2X1 U2209 (.A1(N4417), .A2(N4418), .ZN(n15081));
    NANDX1 U2210 (.A1(N4419), .A2(N4420), .ZN(n15082));
    NOR2X1 U2211 (.A1(N4421), .A2(N4422), .ZN(n15083));
    NANDX1 U2212 (.A1(N4423), .A2(N4424), .ZN(n15084));
    NANDX1 U2213 (.A1(N4425), .A2(N4426), .ZN(N15085));
    NOR2X1 U2214 (.A1(N4427), .A2(N4428), .ZN(n15086));
    NOR2X1 U2215 (.A1(N4429), .A2(N4430), .ZN(n15087));
    NANDX1 U2216 (.A1(N4431), .A2(N4432), .ZN(n15088));
    NOR2X1 U2217 (.A1(N4433), .A2(N4434), .ZN(n15089));
    NOR2X1 U2218 (.A1(N4435), .A2(N4436), .ZN(N15090));
    NOR2X1 U2219 (.A1(N4437), .A2(N4438), .ZN(n15091));
    NANDX1 U2220 (.A1(N4439), .A2(N4440), .ZN(n15092));
    NANDX1 U2221 (.A1(N4441), .A2(N4442), .ZN(n15093));
    NOR2X1 U2222 (.A1(N4443), .A2(N4444), .ZN(n15094));
    NANDX1 U2223 (.A1(N4445), .A2(N4446), .ZN(n15095));
    NOR2X1 U2224 (.A1(N4447), .A2(N4448), .ZN(n15096));
    NANDX1 U2225 (.A1(N4449), .A2(N4450), .ZN(n15097));
    NOR2X1 U2226 (.A1(N4451), .A2(N4452), .ZN(n15098));
    NOR2X1 U2227 (.A1(N4453), .A2(N4454), .ZN(n15099));
    NANDX1 U2228 (.A1(N4455), .A2(N4456), .ZN(N15100));
    NANDX1 U2229 (.A1(N4457), .A2(N4458), .ZN(N15101));
    NOR2X1 U2230 (.A1(N4459), .A2(N4460), .ZN(n15102));
    NOR2X1 U2231 (.A1(N4461), .A2(N4462), .ZN(n15103));
    NOR2X1 U2232 (.A1(N4463), .A2(N4464), .ZN(N15104));
    NOR2X1 U2233 (.A1(N4465), .A2(N4466), .ZN(N15105));
    NOR2X1 U2234 (.A1(N4467), .A2(N4468), .ZN(n15106));
    NANDX1 U2235 (.A1(N4469), .A2(N4470), .ZN(N15107));
    NANDX1 U2236 (.A1(N4471), .A2(N4472), .ZN(n15108));
    NANDX1 U2237 (.A1(N4473), .A2(N4474), .ZN(n15109));
    NANDX1 U2238 (.A1(N4475), .A2(N4476), .ZN(N15110));
    NANDX1 U2239 (.A1(N4477), .A2(N4478), .ZN(N15111));
    NANDX1 U2240 (.A1(N4479), .A2(N4480), .ZN(n15112));
    NOR2X1 U2241 (.A1(N4481), .A2(N4482), .ZN(n15113));
    NOR2X1 U2242 (.A1(N4483), .A2(N4484), .ZN(N15114));
    NANDX1 U2243 (.A1(N4485), .A2(N4486), .ZN(n15115));
    NANDX1 U2244 (.A1(N4487), .A2(N4488), .ZN(n15116));
    NOR2X1 U2245 (.A1(N4489), .A2(N4490), .ZN(n15117));
    NANDX1 U2246 (.A1(N4491), .A2(N4492), .ZN(n15118));
    NANDX1 U2247 (.A1(N4493), .A2(N4494), .ZN(n15119));
    NOR2X1 U2248 (.A1(N4495), .A2(N4496), .ZN(n15120));
    NANDX1 U2249 (.A1(N4497), .A2(N4498), .ZN(n15121));
    NANDX1 U2250 (.A1(N4499), .A2(N4500), .ZN(n15122));
    NOR2X1 U2251 (.A1(N4501), .A2(N4502), .ZN(n15123));
    NOR2X1 U2252 (.A1(N4503), .A2(N4504), .ZN(n15124));
    NANDX1 U2253 (.A1(N4505), .A2(N4506), .ZN(n15125));
    NANDX1 U2254 (.A1(N4507), .A2(N4508), .ZN(N15126));
    NOR2X1 U2255 (.A1(N4509), .A2(N4510), .ZN(n15127));
    NOR2X1 U2256 (.A1(N4511), .A2(N4512), .ZN(n15128));
    NANDX1 U2257 (.A1(N4513), .A2(N4514), .ZN(n15129));
    NOR2X1 U2258 (.A1(N4515), .A2(N4516), .ZN(n15130));
    NANDX1 U2259 (.A1(N4517), .A2(N4518), .ZN(n15131));
    NOR2X1 U2260 (.A1(N4519), .A2(N4520), .ZN(n15132));
    NOR2X1 U2261 (.A1(N4521), .A2(N4522), .ZN(n15133));
    NANDX1 U2262 (.A1(N4523), .A2(N4524), .ZN(N15134));
    NOR2X1 U2263 (.A1(N4525), .A2(N4526), .ZN(n15135));
    NANDX1 U2264 (.A1(N4527), .A2(N4528), .ZN(n15136));
    NANDX1 U2265 (.A1(N4529), .A2(N4530), .ZN(n15137));
    NANDX1 U2266 (.A1(N4531), .A2(N4532), .ZN(n15138));
    NOR2X1 U2267 (.A1(N4533), .A2(N4534), .ZN(n15139));
    NOR2X1 U2268 (.A1(N4535), .A2(N4536), .ZN(n15140));
    NOR2X1 U2269 (.A1(N4537), .A2(N4538), .ZN(n15141));
    NOR2X1 U2270 (.A1(N4539), .A2(N4540), .ZN(n15142));
    NANDX1 U2271 (.A1(N4541), .A2(N4542), .ZN(n15143));
    NOR2X1 U2272 (.A1(N4543), .A2(N4544), .ZN(N15144));
    NOR2X1 U2273 (.A1(N4545), .A2(N4546), .ZN(n15145));
    NOR2X1 U2274 (.A1(N4547), .A2(N4548), .ZN(n15146));
    NOR2X1 U2275 (.A1(N4549), .A2(N4550), .ZN(n15147));
    NOR2X1 U2276 (.A1(N4551), .A2(N4552), .ZN(N15148));
    NANDX1 U2277 (.A1(N4553), .A2(N4554), .ZN(n15149));
    NANDX1 U2278 (.A1(N4555), .A2(N4556), .ZN(n15150));
    NOR2X1 U2279 (.A1(N4557), .A2(N4558), .ZN(n15151));
    NOR2X1 U2280 (.A1(N4559), .A2(N4560), .ZN(N15152));
    NOR2X1 U2281 (.A1(N4561), .A2(N4562), .ZN(n15153));
    NOR2X1 U2282 (.A1(N4563), .A2(N4564), .ZN(n15154));
    NANDX1 U2283 (.A1(N4565), .A2(N4566), .ZN(n15155));
    NANDX1 U2284 (.A1(N4567), .A2(N4568), .ZN(N15156));
    NANDX1 U2285 (.A1(N4569), .A2(N4570), .ZN(n15157));
    NANDX1 U2286 (.A1(N4571), .A2(N4572), .ZN(N15158));
    NANDX1 U2287 (.A1(N4573), .A2(N4574), .ZN(n15159));
    NANDX1 U2288 (.A1(N4575), .A2(N4576), .ZN(n15160));
    NOR2X1 U2289 (.A1(N4577), .A2(N4578), .ZN(n15161));
    NOR2X1 U2290 (.A1(N4579), .A2(N4580), .ZN(n15162));
    NANDX1 U2291 (.A1(N4581), .A2(N4582), .ZN(n15163));
    NOR2X1 U2292 (.A1(N4583), .A2(N4584), .ZN(n15164));
    NANDX1 U2293 (.A1(N4585), .A2(N4586), .ZN(n15165));
    NOR2X1 U2294 (.A1(N4587), .A2(N4588), .ZN(n15166));
    NANDX1 U2295 (.A1(N4589), .A2(N4590), .ZN(n15167));
    NOR2X1 U2296 (.A1(N4591), .A2(N4592), .ZN(n15168));
    NANDX1 U2297 (.A1(N4593), .A2(N4594), .ZN(N15169));
    NOR2X1 U2298 (.A1(N4595), .A2(N4596), .ZN(N15170));
    NOR2X1 U2299 (.A1(N4597), .A2(N4598), .ZN(N15171));
    NOR2X1 U2300 (.A1(N4599), .A2(N4600), .ZN(n15172));
    NOR2X1 U2301 (.A1(N4601), .A2(N4602), .ZN(N15173));
    NANDX1 U2302 (.A1(N4603), .A2(N4604), .ZN(N15174));
    NOR2X1 U2303 (.A1(N4605), .A2(N4606), .ZN(n15175));
    NOR2X1 U2304 (.A1(N4607), .A2(N4608), .ZN(n15176));
    NOR2X1 U2305 (.A1(N4609), .A2(N4610), .ZN(n15177));
    NOR2X1 U2306 (.A1(N4611), .A2(N4612), .ZN(n15178));
    NOR2X1 U2307 (.A1(N4613), .A2(N4614), .ZN(n15179));
    NANDX1 U2308 (.A1(N4615), .A2(N4616), .ZN(n15180));
    NANDX1 U2309 (.A1(N4617), .A2(N4618), .ZN(n15181));
    NOR2X1 U2310 (.A1(N4619), .A2(N4620), .ZN(n15182));
    NOR2X1 U2311 (.A1(N4621), .A2(N4622), .ZN(N15183));
    NANDX1 U2312 (.A1(N4623), .A2(N4624), .ZN(n15184));
    NANDX1 U2313 (.A1(N4625), .A2(N4626), .ZN(N15185));
    NANDX1 U2314 (.A1(N4627), .A2(N4628), .ZN(n15186));
    NOR2X1 U2315 (.A1(N4629), .A2(N4630), .ZN(n15187));
    NOR2X1 U2316 (.A1(N4631), .A2(N4632), .ZN(n15188));
    NOR2X1 U2317 (.A1(N4633), .A2(N4634), .ZN(n15189));
    NANDX1 U2318 (.A1(N4635), .A2(N4636), .ZN(n15190));
    NANDX1 U2319 (.A1(N4637), .A2(N4638), .ZN(n15191));
    NOR2X1 U2320 (.A1(N4639), .A2(N4640), .ZN(n15192));
    NANDX1 U2321 (.A1(N4641), .A2(N4642), .ZN(n15193));
    NANDX1 U2322 (.A1(N4643), .A2(N4644), .ZN(n15194));
    NANDX1 U2323 (.A1(N4645), .A2(N4646), .ZN(n15195));
    NOR2X1 U2324 (.A1(N4647), .A2(N4648), .ZN(n15196));
    NANDX1 U2325 (.A1(N4649), .A2(N4650), .ZN(n15197));
    NOR2X1 U2326 (.A1(N4651), .A2(N4652), .ZN(n15198));
    NOR2X1 U2327 (.A1(N4653), .A2(N4654), .ZN(N15199));
    NOR2X1 U2328 (.A1(N4655), .A2(N4656), .ZN(n15200));
    NOR2X1 U2329 (.A1(N4657), .A2(N4658), .ZN(N15201));
    NOR2X1 U2330 (.A1(N4659), .A2(N4660), .ZN(n15202));
    NOR2X1 U2331 (.A1(N4661), .A2(N4662), .ZN(n15203));
    NOR2X1 U2332 (.A1(N4663), .A2(N4664), .ZN(n15204));
    NOR2X1 U2333 (.A1(N4665), .A2(N4666), .ZN(n15205));
    NANDX1 U2334 (.A1(N4667), .A2(N4668), .ZN(n15206));
    NOR2X1 U2335 (.A1(N4669), .A2(N4670), .ZN(n15207));
    NOR2X1 U2336 (.A1(N4671), .A2(N4672), .ZN(n15208));
    NANDX1 U2337 (.A1(N4673), .A2(N4674), .ZN(N15209));
    NOR2X1 U2338 (.A1(N4675), .A2(N4676), .ZN(n15210));
    NANDX1 U2339 (.A1(N4677), .A2(N4678), .ZN(n15211));
    NANDX1 U2340 (.A1(N4679), .A2(N4680), .ZN(n15212));
    NANDX1 U2341 (.A1(N4681), .A2(N4682), .ZN(n15213));
    NANDX1 U2342 (.A1(N4683), .A2(N4684), .ZN(N15214));
    NOR2X1 U2343 (.A1(N4685), .A2(N4686), .ZN(n15215));
    NOR2X1 U2344 (.A1(N4687), .A2(N4688), .ZN(n15216));
    NOR2X1 U2345 (.A1(N4689), .A2(N4690), .ZN(N15217));
    NANDX1 U2346 (.A1(N4691), .A2(N4692), .ZN(n15218));
    NOR2X1 U2347 (.A1(N4693), .A2(N4694), .ZN(n15219));
    NANDX1 U2348 (.A1(N4695), .A2(N4696), .ZN(n15220));
    NOR2X1 U2349 (.A1(N4697), .A2(N4698), .ZN(n15221));
    NOR2X1 U2350 (.A1(N4699), .A2(N4700), .ZN(n15222));
    NANDX1 U2351 (.A1(N4701), .A2(N4702), .ZN(n15223));
    NOR2X1 U2352 (.A1(N4703), .A2(N4704), .ZN(N15224));
    NANDX1 U2353 (.A1(N4705), .A2(N4706), .ZN(n15225));
    NOR2X1 U2354 (.A1(N4707), .A2(N4708), .ZN(n15226));
    NOR2X1 U2355 (.A1(N4709), .A2(N4710), .ZN(n15227));
    NOR2X1 U2356 (.A1(N4711), .A2(N4712), .ZN(N15228));
    NANDX1 U2357 (.A1(N4713), .A2(N4714), .ZN(n15229));
    NANDX1 U2358 (.A1(N4715), .A2(N4716), .ZN(n15230));
    NOR2X1 U2359 (.A1(N4717), .A2(N4718), .ZN(n15231));
    NANDX1 U2360 (.A1(N4719), .A2(N4720), .ZN(n15232));
    NANDX1 U2361 (.A1(N4721), .A2(N4722), .ZN(N15233));
    NANDX1 U2362 (.A1(N4723), .A2(N4724), .ZN(n15234));
    NOR2X1 U2363 (.A1(N4725), .A2(N4726), .ZN(n15235));
    NANDX1 U2364 (.A1(N4727), .A2(N4728), .ZN(n15236));
    NOR2X1 U2365 (.A1(N4729), .A2(N4730), .ZN(n15237));
    NOR2X1 U2366 (.A1(N4731), .A2(N4732), .ZN(n15238));
    NANDX1 U2367 (.A1(N4733), .A2(N4734), .ZN(n15239));
    NANDX1 U2368 (.A1(N4735), .A2(N4736), .ZN(n15240));
    NANDX1 U2369 (.A1(N4737), .A2(N4738), .ZN(n15241));
    NANDX1 U2370 (.A1(N4739), .A2(N4740), .ZN(n15242));
    NOR2X1 U2371 (.A1(N4741), .A2(N4742), .ZN(n15243));
    NOR2X1 U2372 (.A1(N4743), .A2(N4744), .ZN(n15244));
    NOR2X1 U2373 (.A1(N4745), .A2(N4746), .ZN(n15245));
    NANDX1 U2374 (.A1(N4747), .A2(N4748), .ZN(n15246));
    NOR2X1 U2375 (.A1(N4749), .A2(N4750), .ZN(n15247));
    NANDX1 U2376 (.A1(N4751), .A2(N4752), .ZN(n15248));
    NOR2X1 U2377 (.A1(N4753), .A2(N4754), .ZN(N15249));
    NOR2X1 U2378 (.A1(N4755), .A2(N4756), .ZN(n15250));
    NOR2X1 U2379 (.A1(N4757), .A2(N4758), .ZN(n15251));
    NOR2X1 U2380 (.A1(N4759), .A2(N4760), .ZN(n15252));
    NOR2X1 U2381 (.A1(N4761), .A2(N4762), .ZN(n15253));
    NANDX1 U2382 (.A1(N4763), .A2(N4764), .ZN(N15254));
    NOR2X1 U2383 (.A1(N4765), .A2(N4766), .ZN(N15255));
    NANDX1 U2384 (.A1(N4767), .A2(N4768), .ZN(n15256));
    NOR2X1 U2385 (.A1(N4769), .A2(N4770), .ZN(N15257));
    NANDX1 U2386 (.A1(N4771), .A2(N4772), .ZN(n15258));
    NANDX1 U2387 (.A1(N4773), .A2(N4774), .ZN(N15259));
    NANDX1 U2388 (.A1(N4775), .A2(N4776), .ZN(N15260));
    NOR2X1 U2389 (.A1(N4777), .A2(N4778), .ZN(n15261));
    NOR2X1 U2390 (.A1(N4779), .A2(N4780), .ZN(n15262));
    NOR2X1 U2391 (.A1(N4781), .A2(N4782), .ZN(n15263));
    NANDX1 U2392 (.A1(N4783), .A2(N4784), .ZN(n15264));
    NANDX1 U2393 (.A1(N4785), .A2(N4786), .ZN(n15265));
    NOR2X1 U2394 (.A1(N4787), .A2(N4788), .ZN(n15266));
    NANDX1 U2395 (.A1(N4789), .A2(N4790), .ZN(n15267));
    NANDX1 U2396 (.A1(N4791), .A2(N4792), .ZN(n15268));
    NANDX1 U2397 (.A1(N4793), .A2(N4794), .ZN(n15269));
    NOR2X1 U2398 (.A1(N4795), .A2(N4796), .ZN(n15270));
    NOR2X1 U2399 (.A1(N4797), .A2(N4798), .ZN(n15271));
    NOR2X1 U2400 (.A1(N4799), .A2(N4800), .ZN(n15272));
    NANDX1 U2401 (.A1(N4801), .A2(N4802), .ZN(n15273));
    NANDX1 U2402 (.A1(N4803), .A2(N4804), .ZN(N15274));
    NOR2X1 U2403 (.A1(N4805), .A2(N4806), .ZN(n15275));
    NOR2X1 U2404 (.A1(N4807), .A2(N4808), .ZN(n15276));
    NOR2X1 U2405 (.A1(N4809), .A2(N4810), .ZN(n15277));
    NOR2X1 U2406 (.A1(N4811), .A2(N4812), .ZN(N15278));
    NANDX1 U2407 (.A1(N4813), .A2(N4814), .ZN(n15279));
    NOR2X1 U2408 (.A1(N4815), .A2(N4816), .ZN(n15280));
    NOR2X1 U2409 (.A1(N4817), .A2(N4818), .ZN(n15281));
    NANDX1 U2410 (.A1(N4819), .A2(N4820), .ZN(n15282));
    NOR2X1 U2411 (.A1(N4821), .A2(N4822), .ZN(n15283));
    NANDX1 U2412 (.A1(N4823), .A2(N4824), .ZN(n15284));
    NOR2X1 U2413 (.A1(N4825), .A2(N4826), .ZN(n15285));
    NANDX1 U2414 (.A1(N4827), .A2(N4828), .ZN(n15286));
    NOR2X1 U2415 (.A1(N4829), .A2(N4830), .ZN(n15287));
    NOR2X1 U2416 (.A1(N4831), .A2(N4832), .ZN(n15288));
    NOR2X1 U2417 (.A1(N4833), .A2(N4834), .ZN(n15289));
    NOR2X1 U2418 (.A1(N4835), .A2(N4836), .ZN(n15290));
    NANDX1 U2419 (.A1(N4837), .A2(N4838), .ZN(N15291));
    NOR2X1 U2420 (.A1(N4839), .A2(N4840), .ZN(n15292));
    NOR2X1 U2421 (.A1(N4841), .A2(N4842), .ZN(n15293));
    NOR2X1 U2422 (.A1(N4843), .A2(N4844), .ZN(N15294));
    NANDX1 U2423 (.A1(N4845), .A2(N4846), .ZN(n15295));
    NANDX1 U2424 (.A1(N4847), .A2(N4848), .ZN(N15296));
    NOR2X1 U2425 (.A1(N4849), .A2(N4850), .ZN(n15297));
    NOR2X1 U2426 (.A1(N4851), .A2(N4852), .ZN(n15298));
    NOR2X1 U2427 (.A1(N4853), .A2(N4854), .ZN(n15299));
    NANDX1 U2428 (.A1(N4855), .A2(N4856), .ZN(n15300));
    NANDX1 U2429 (.A1(N4857), .A2(N4858), .ZN(n15301));
    NOR2X1 U2430 (.A1(N4859), .A2(N4860), .ZN(n15302));
    NANDX1 U2431 (.A1(N4861), .A2(N4862), .ZN(N15303));
    NOR2X1 U2432 (.A1(N4863), .A2(N4864), .ZN(N15304));
    NANDX1 U2433 (.A1(N4865), .A2(N4866), .ZN(n15305));
    NANDX1 U2434 (.A1(N4867), .A2(N4868), .ZN(n15306));
    NOR2X1 U2435 (.A1(N4869), .A2(N4870), .ZN(N15307));
    NANDX1 U2436 (.A1(N4871), .A2(N4872), .ZN(N15308));
    NANDX1 U2437 (.A1(N4873), .A2(N4874), .ZN(n15309));
    NANDX1 U2438 (.A1(N4875), .A2(N4876), .ZN(N15310));
    NANDX1 U2439 (.A1(N4877), .A2(N4878), .ZN(n15311));
    NOR2X1 U2440 (.A1(N4879), .A2(N4880), .ZN(n15312));
    NOR2X1 U2441 (.A1(N4881), .A2(N4882), .ZN(N15313));
    NOR2X1 U2442 (.A1(N4883), .A2(N4884), .ZN(n15314));
    NANDX1 U2443 (.A1(N4885), .A2(N4886), .ZN(n15315));
    NANDX1 U2444 (.A1(N4887), .A2(N4888), .ZN(n15316));
    NANDX1 U2445 (.A1(N4889), .A2(N4890), .ZN(N15317));
    NANDX1 U2446 (.A1(N4891), .A2(N4892), .ZN(n15318));
    NANDX1 U2447 (.A1(N4893), .A2(N4894), .ZN(N15319));
    NANDX1 U2448 (.A1(N4895), .A2(N4896), .ZN(n15320));
    NANDX1 U2449 (.A1(N4897), .A2(N4898), .ZN(n15321));
    NANDX1 U2450 (.A1(N4899), .A2(N4900), .ZN(n15322));
    NANDX1 U2451 (.A1(N4901), .A2(N4902), .ZN(N15323));
    NANDX1 U2452 (.A1(N4903), .A2(N4904), .ZN(n15324));
    NANDX1 U2453 (.A1(N4905), .A2(N4906), .ZN(n15325));
    NOR2X1 U2454 (.A1(N4907), .A2(N4908), .ZN(n15326));
    NOR2X1 U2455 (.A1(N4909), .A2(N4910), .ZN(n15327));
    NANDX1 U2456 (.A1(N4911), .A2(N4912), .ZN(n15328));
    NANDX1 U2457 (.A1(N4913), .A2(N4914), .ZN(n15329));
    NOR2X1 U2458 (.A1(N4915), .A2(N4916), .ZN(n15330));
    NANDX1 U2459 (.A1(N4917), .A2(N4918), .ZN(N15331));
    NOR2X1 U2460 (.A1(N4919), .A2(N4920), .ZN(n15332));
    NANDX1 U2461 (.A1(N4921), .A2(N4922), .ZN(n15333));
    NOR2X1 U2462 (.A1(N4923), .A2(N4924), .ZN(n15334));
    NOR2X1 U2463 (.A1(N4925), .A2(N4926), .ZN(n15335));
    NOR2X1 U2464 (.A1(N4927), .A2(N4928), .ZN(n15336));
    NOR2X1 U2465 (.A1(N4929), .A2(N4930), .ZN(n15337));
    NANDX1 U2466 (.A1(N4931), .A2(N4932), .ZN(n15338));
    NOR2X1 U2467 (.A1(N4933), .A2(N4934), .ZN(n15339));
    NANDX1 U2468 (.A1(N4935), .A2(N4936), .ZN(n15340));
    NOR2X1 U2469 (.A1(N4937), .A2(N4938), .ZN(n15341));
    NANDX1 U2470 (.A1(N4939), .A2(N4940), .ZN(n15342));
    NANDX1 U2471 (.A1(N4941), .A2(N4942), .ZN(n15343));
    NANDX1 U2472 (.A1(N4943), .A2(N4944), .ZN(n15344));
    NANDX1 U2473 (.A1(N4945), .A2(N4946), .ZN(n15345));
    NOR2X1 U2474 (.A1(N4947), .A2(N4948), .ZN(N15346));
    NOR2X1 U2475 (.A1(N4949), .A2(N4950), .ZN(n15347));
    NOR2X1 U2476 (.A1(N4951), .A2(N4952), .ZN(n15348));
    NOR2X1 U2477 (.A1(N4953), .A2(N4954), .ZN(n15349));
    NANDX1 U2478 (.A1(N4955), .A2(N4956), .ZN(n15350));
    NANDX1 U2479 (.A1(N4957), .A2(N4958), .ZN(n15351));
    NANDX1 U2480 (.A1(N4959), .A2(N4960), .ZN(n15352));
    NOR2X1 U2481 (.A1(N4961), .A2(N4962), .ZN(N15353));
    NOR2X1 U2482 (.A1(N4963), .A2(N4964), .ZN(N15354));
    NANDX1 U2483 (.A1(N4965), .A2(N4966), .ZN(n15355));
    NANDX1 U2484 (.A1(N4967), .A2(N4968), .ZN(n15356));
    NANDX1 U2485 (.A1(N4969), .A2(N4970), .ZN(n15357));
    NANDX1 U2486 (.A1(N4971), .A2(N4972), .ZN(n15358));
    NANDX1 U2487 (.A1(N4973), .A2(N4974), .ZN(n15359));
    NOR2X1 U2488 (.A1(N4975), .A2(N4976), .ZN(n15360));
    NOR2X1 U2489 (.A1(N4977), .A2(N4978), .ZN(n15361));
    NOR2X1 U2490 (.A1(N4979), .A2(N4980), .ZN(N15362));
    NOR2X1 U2491 (.A1(N4981), .A2(N4982), .ZN(n15363));
    NANDX1 U2492 (.A1(N4983), .A2(N4984), .ZN(n15364));
    NOR2X1 U2493 (.A1(N4985), .A2(N4986), .ZN(n15365));
    NOR2X1 U2494 (.A1(N4987), .A2(N4988), .ZN(N15366));
    NANDX1 U2495 (.A1(N4989), .A2(N4990), .ZN(n15367));
    NOR2X1 U2496 (.A1(N4991), .A2(N4992), .ZN(n15368));
    NANDX1 U2497 (.A1(N4993), .A2(N4994), .ZN(n15369));
    NANDX1 U2498 (.A1(N4995), .A2(N4996), .ZN(n15370));
    NOR2X1 U2499 (.A1(N4997), .A2(N4998), .ZN(n15371));
    NOR2X1 U2500 (.A1(N4999), .A2(N5000), .ZN(n15372));
    NANDX1 U2501 (.A1(N5001), .A2(N5002), .ZN(n15373));
    NANDX1 U2502 (.A1(N5003), .A2(N5004), .ZN(n15374));
    NANDX1 U2503 (.A1(N5005), .A2(N5006), .ZN(n15375));
    NOR2X1 U2504 (.A1(N5007), .A2(N5008), .ZN(n15376));
    NOR2X1 U2505 (.A1(N5009), .A2(N5010), .ZN(n15377));
    NANDX1 U2506 (.A1(N5011), .A2(N5012), .ZN(n15378));
    NANDX1 U2507 (.A1(N5013), .A2(N5014), .ZN(N15379));
    NOR2X1 U2508 (.A1(N5015), .A2(N5016), .ZN(n15380));
    NOR2X1 U2509 (.A1(N5017), .A2(N5018), .ZN(n15381));
    NOR2X1 U2510 (.A1(N5019), .A2(N5020), .ZN(n15382));
    NANDX1 U2511 (.A1(N5021), .A2(N5022), .ZN(n15383));
    NANDX1 U2512 (.A1(N5023), .A2(N5024), .ZN(n15384));
    NANDX1 U2513 (.A1(N5025), .A2(N5026), .ZN(n15385));
    NOR2X1 U2514 (.A1(N5027), .A2(N5028), .ZN(n15386));
    NOR2X1 U2515 (.A1(N5029), .A2(N5030), .ZN(n15387));
    NOR2X1 U2516 (.A1(N5031), .A2(N5032), .ZN(n15388));
    NOR2X1 U2517 (.A1(N5033), .A2(N5034), .ZN(n15389));
    NANDX1 U2518 (.A1(N5035), .A2(N5036), .ZN(N15390));
    NOR2X1 U2519 (.A1(N5037), .A2(N5038), .ZN(n15391));
    NOR2X1 U2520 (.A1(N5039), .A2(N5040), .ZN(n15392));
    NANDX1 U2521 (.A1(N5041), .A2(N5042), .ZN(n15393));
    NOR2X1 U2522 (.A1(N5043), .A2(N5044), .ZN(n15394));
    NANDX1 U2523 (.A1(N5045), .A2(N5046), .ZN(n15395));
    NOR2X1 U2524 (.A1(N5047), .A2(N5048), .ZN(n15396));
    NOR2X1 U2525 (.A1(N5049), .A2(N5050), .ZN(n15397));
    NOR2X1 U2526 (.A1(N5051), .A2(N5052), .ZN(n15398));
    NOR2X1 U2527 (.A1(N5053), .A2(N5054), .ZN(n15399));
    NOR2X1 U2528 (.A1(N5055), .A2(N5056), .ZN(n15400));
    NOR2X1 U2529 (.A1(N5057), .A2(N5058), .ZN(n15401));
    NOR2X1 U2530 (.A1(N5059), .A2(N5060), .ZN(N15402));
    NOR2X1 U2531 (.A1(N5061), .A2(N5062), .ZN(N15403));
    NANDX1 U2532 (.A1(N5063), .A2(N5064), .ZN(n15404));
    NOR2X1 U2533 (.A1(N5065), .A2(N5066), .ZN(n15405));
    NANDX1 U2534 (.A1(N5067), .A2(N5068), .ZN(n15406));
    NANDX1 U2535 (.A1(N5069), .A2(N5070), .ZN(n15407));
    NOR2X1 U2536 (.A1(N5071), .A2(N5072), .ZN(n15408));
    NOR2X1 U2537 (.A1(N5073), .A2(N5074), .ZN(n15409));
    NOR2X1 U2538 (.A1(N5075), .A2(N5076), .ZN(N15410));
    NOR2X1 U2539 (.A1(N5077), .A2(N5078), .ZN(n15411));
    NOR2X1 U2540 (.A1(N5079), .A2(N5080), .ZN(n15412));
    NANDX1 U2541 (.A1(N5081), .A2(N5082), .ZN(n15413));
    NANDX1 U2542 (.A1(N5083), .A2(N5084), .ZN(n15414));
    NANDX1 U2543 (.A1(N5085), .A2(N5086), .ZN(n15415));
    NOR2X1 U2544 (.A1(N5087), .A2(N5088), .ZN(n15416));
    NOR2X1 U2545 (.A1(N5089), .A2(N5090), .ZN(n15417));
    NOR2X1 U2546 (.A1(N5091), .A2(N5092), .ZN(n15418));
    NOR2X1 U2547 (.A1(N5093), .A2(N5094), .ZN(n15419));
    NOR2X1 U2548 (.A1(N5095), .A2(N5096), .ZN(n15420));
    NANDX1 U2549 (.A1(N5097), .A2(N5098), .ZN(n15421));
    NOR2X1 U2550 (.A1(N5099), .A2(N5100), .ZN(N15422));
    NOR2X1 U2551 (.A1(N5101), .A2(N5102), .ZN(n15423));
    NANDX1 U2552 (.A1(N5103), .A2(N5104), .ZN(n15424));
    NOR2X1 U2553 (.A1(N5105), .A2(N5106), .ZN(n15425));
    NANDX1 U2554 (.A1(N5107), .A2(N5108), .ZN(n15426));
    NANDX1 U2555 (.A1(N5109), .A2(N5110), .ZN(n15427));
    NOR2X1 U2556 (.A1(N5111), .A2(N5112), .ZN(n15428));
    NANDX1 U2557 (.A1(N5113), .A2(N5114), .ZN(n15429));
    NANDX1 U2558 (.A1(N5115), .A2(N5116), .ZN(n15430));
    NOR2X1 U2559 (.A1(N5117), .A2(N5118), .ZN(n15431));
    NANDX1 U2560 (.A1(N5119), .A2(N5120), .ZN(n15432));
    NOR2X1 U2561 (.A1(N5121), .A2(N5122), .ZN(n15433));
    NOR2X1 U2562 (.A1(N5123), .A2(N5124), .ZN(N15434));
    NOR2X1 U2563 (.A1(N5125), .A2(N5126), .ZN(n15435));
    NOR2X1 U2564 (.A1(N5127), .A2(N5128), .ZN(n15436));
    NANDX1 U2565 (.A1(N5129), .A2(N5130), .ZN(n15437));
    NOR2X1 U2566 (.A1(N5131), .A2(N5132), .ZN(n15438));
    NOR2X1 U2567 (.A1(N5133), .A2(N5134), .ZN(n15439));
    NANDX1 U2568 (.A1(N5135), .A2(N5136), .ZN(n15440));
    NOR2X1 U2569 (.A1(N5137), .A2(N5138), .ZN(n15441));
    NOR2X1 U2570 (.A1(N5139), .A2(N5140), .ZN(N15442));
    NOR2X1 U2571 (.A1(N5141), .A2(N5142), .ZN(n15443));
    NANDX1 U2572 (.A1(N5143), .A2(N5144), .ZN(N15444));
    NANDX1 U2573 (.A1(N5145), .A2(N5146), .ZN(n15445));
    NANDX1 U2574 (.A1(N5147), .A2(N5148), .ZN(n15446));
    NANDX1 U2575 (.A1(N5149), .A2(N5150), .ZN(n15447));
    NANDX1 U2576 (.A1(N5151), .A2(N5152), .ZN(n15448));
    NANDX1 U2577 (.A1(N5153), .A2(N5154), .ZN(n15449));
    NANDX1 U2578 (.A1(N5155), .A2(N5156), .ZN(n15450));
    NANDX1 U2579 (.A1(N5157), .A2(N5158), .ZN(n15451));
    NANDX1 U2580 (.A1(N5159), .A2(N5160), .ZN(n15452));
    NANDX1 U2581 (.A1(N5161), .A2(N5162), .ZN(N15453));
    NANDX1 U2582 (.A1(N5163), .A2(N5164), .ZN(n15454));
    NOR2X1 U2583 (.A1(N5165), .A2(N5166), .ZN(N15455));
    NANDX1 U2584 (.A1(N5167), .A2(N5168), .ZN(n15456));
    NOR2X1 U2585 (.A1(N5169), .A2(N5170), .ZN(n15457));
    NANDX1 U2586 (.A1(N5171), .A2(N5172), .ZN(n15458));
    NOR2X1 U2587 (.A1(N5173), .A2(N5174), .ZN(n15459));
    NOR2X1 U2588 (.A1(N5175), .A2(N5176), .ZN(n15460));
    NOR2X1 U2589 (.A1(N5177), .A2(N5178), .ZN(n15461));
    NOR2X1 U2590 (.A1(N5179), .A2(N5180), .ZN(n15462));
    NANDX1 U2591 (.A1(N5181), .A2(N5182), .ZN(n15463));
    NOR2X1 U2592 (.A1(N5183), .A2(N5184), .ZN(n15464));
    NANDX1 U2593 (.A1(N5185), .A2(N5186), .ZN(n15465));
    NOR2X1 U2594 (.A1(N5187), .A2(N5188), .ZN(n15466));
    NOR2X1 U2595 (.A1(N5189), .A2(N5190), .ZN(n15467));
    NOR2X1 U2596 (.A1(N5191), .A2(N5192), .ZN(n15468));
    NOR2X1 U2597 (.A1(N5193), .A2(N5194), .ZN(N15469));
    NOR2X1 U2598 (.A1(N5195), .A2(N5196), .ZN(n15470));
    NOR2X1 U2599 (.A1(N5197), .A2(N5198), .ZN(n15471));
    NOR2X1 U2600 (.A1(N5199), .A2(N5200), .ZN(n15472));
    NOR2X1 U2601 (.A1(N5201), .A2(N5202), .ZN(N15473));
    NOR2X1 U2602 (.A1(N5203), .A2(N5204), .ZN(n15474));
    NOR2X1 U2603 (.A1(N5205), .A2(N5206), .ZN(n15475));
    NOR2X1 U2604 (.A1(N5207), .A2(N5208), .ZN(n15476));
    NANDX1 U2605 (.A1(N5209), .A2(N5210), .ZN(n15477));
    NANDX1 U2606 (.A1(N5211), .A2(N5212), .ZN(n15478));
    NANDX1 U2607 (.A1(N5213), .A2(N5214), .ZN(n15479));
    NANDX1 U2608 (.A1(N5215), .A2(N5216), .ZN(n15480));
    NANDX1 U2609 (.A1(N5217), .A2(N5218), .ZN(n15481));
    NANDX1 U2610 (.A1(N5219), .A2(N5220), .ZN(n15482));
    NOR2X1 U2611 (.A1(N5221), .A2(N5222), .ZN(n15483));
    NOR2X1 U2612 (.A1(N5223), .A2(N5224), .ZN(n15484));
    NOR2X1 U2613 (.A1(N5225), .A2(N5226), .ZN(N15485));
    NOR2X1 U2614 (.A1(N5227), .A2(N5228), .ZN(n15486));
    NOR2X1 U2615 (.A1(N5229), .A2(N5230), .ZN(n15487));
    NANDX1 U2616 (.A1(N5231), .A2(N5232), .ZN(n15488));
    NANDX1 U2617 (.A1(N5233), .A2(N5234), .ZN(N15489));
    NOR2X1 U2618 (.A1(N5235), .A2(N5236), .ZN(n15490));
    NANDX1 U2619 (.A1(N5237), .A2(N5238), .ZN(n15491));
    NANDX1 U2620 (.A1(N5239), .A2(N5240), .ZN(n15492));
    NOR2X1 U2621 (.A1(N5241), .A2(N5242), .ZN(n15493));
    NOR2X1 U2622 (.A1(N5243), .A2(N5244), .ZN(N15494));
    NOR2X1 U2623 (.A1(N5245), .A2(N5246), .ZN(n15495));
    NANDX1 U2624 (.A1(N5247), .A2(N5248), .ZN(N15496));
    NOR2X1 U2625 (.A1(N5249), .A2(N5250), .ZN(N15497));
    NOR2X1 U2626 (.A1(N5251), .A2(N5252), .ZN(n15498));
    NOR2X1 U2627 (.A1(N5253), .A2(N5254), .ZN(n15499));
    NOR2X1 U2628 (.A1(N5255), .A2(N5256), .ZN(N15500));
    NANDX1 U2629 (.A1(N5257), .A2(N5258), .ZN(N15501));
    NOR2X1 U2630 (.A1(N5259), .A2(N5260), .ZN(n15502));
    NANDX1 U2631 (.A1(N5261), .A2(N5262), .ZN(n15503));
    NANDX1 U2632 (.A1(N5263), .A2(N5264), .ZN(N15504));
    NOR2X1 U2633 (.A1(N5265), .A2(N5266), .ZN(n15505));
    NANDX1 U2634 (.A1(N5267), .A2(N5268), .ZN(n15506));
    NANDX1 U2635 (.A1(N5269), .A2(N5270), .ZN(n15507));
    NANDX1 U2636 (.A1(N5271), .A2(N5272), .ZN(n15508));
    NOR2X1 U2637 (.A1(N5273), .A2(N5274), .ZN(n15509));
    NANDX1 U2638 (.A1(N5275), .A2(N5276), .ZN(n15510));
    NOR2X1 U2639 (.A1(N5277), .A2(N5278), .ZN(n15511));
    NANDX1 U2640 (.A1(N5279), .A2(N5280), .ZN(n15512));
    NOR2X1 U2641 (.A1(N5281), .A2(N5282), .ZN(N15513));
    NOR2X1 U2642 (.A1(N5283), .A2(N5284), .ZN(n15514));
    NOR2X1 U2643 (.A1(N5285), .A2(N5286), .ZN(n15515));
    NOR2X1 U2644 (.A1(N5287), .A2(N5288), .ZN(N15516));
    NOR2X1 U2645 (.A1(N5289), .A2(N5290), .ZN(n15517));
    NOR2X1 U2646 (.A1(N5291), .A2(N5292), .ZN(n15518));
    NANDX1 U2647 (.A1(N5293), .A2(N5294), .ZN(N15519));
    NANDX1 U2648 (.A1(N5295), .A2(N5296), .ZN(N15520));
    NOR2X1 U2649 (.A1(N5297), .A2(N5298), .ZN(n15521));
    NOR2X1 U2650 (.A1(N5299), .A2(N5300), .ZN(N15522));
    NANDX1 U2651 (.A1(N5301), .A2(N5302), .ZN(n15523));
    NOR2X1 U2652 (.A1(N5303), .A2(N5304), .ZN(n15524));
    NANDX1 U2653 (.A1(N5305), .A2(N5306), .ZN(n15525));
    NANDX1 U2654 (.A1(N5307), .A2(N5308), .ZN(n15526));
    NOR2X1 U2655 (.A1(N5309), .A2(N5310), .ZN(n15527));
    NANDX1 U2656 (.A1(N5311), .A2(N5312), .ZN(n15528));
    NANDX1 U2657 (.A1(N5313), .A2(N5314), .ZN(N15529));
    NOR2X1 U2658 (.A1(N5315), .A2(N5316), .ZN(n15530));
    NOR2X1 U2659 (.A1(N5317), .A2(N5318), .ZN(n15531));
    NOR2X1 U2660 (.A1(N5319), .A2(N5320), .ZN(N15532));
    NOR2X1 U2661 (.A1(N5321), .A2(N5322), .ZN(n15533));
    NANDX1 U2662 (.A1(N5323), .A2(N5324), .ZN(N15534));
    NOR2X1 U2663 (.A1(N5325), .A2(N5326), .ZN(n15535));
    NOR2X1 U2664 (.A1(N5327), .A2(N5328), .ZN(n15536));
    NOR2X1 U2665 (.A1(N5329), .A2(N5330), .ZN(N15537));
    NANDX1 U2666 (.A1(N5331), .A2(N5332), .ZN(n15538));
    NANDX1 U2667 (.A1(N5333), .A2(N5334), .ZN(n15539));
    NOR2X1 U2668 (.A1(N5335), .A2(N5336), .ZN(N15540));
    NOR2X1 U2669 (.A1(N5337), .A2(N5338), .ZN(N15541));
    NOR2X1 U2670 (.A1(N5339), .A2(N5340), .ZN(n15542));
    NOR2X1 U2671 (.A1(N5341), .A2(N5342), .ZN(N15543));
    NOR2X1 U2672 (.A1(N5343), .A2(N5344), .ZN(n15544));
    NOR2X1 U2673 (.A1(N5345), .A2(N5346), .ZN(N15545));
    NOR2X1 U2674 (.A1(N5347), .A2(N5348), .ZN(n15546));
    NANDX1 U2675 (.A1(N5349), .A2(N5350), .ZN(n15547));
    NANDX1 U2676 (.A1(N5351), .A2(N5352), .ZN(n15548));
    NOR2X1 U2677 (.A1(N5353), .A2(N5354), .ZN(n15549));
    NOR2X1 U2678 (.A1(N5355), .A2(N5356), .ZN(N15550));
    NOR2X1 U2679 (.A1(N5357), .A2(N5358), .ZN(n15551));
    NOR2X1 U2680 (.A1(N5359), .A2(N5360), .ZN(n15552));
    NANDX1 U2681 (.A1(N5361), .A2(N5362), .ZN(n15553));
    NANDX1 U2682 (.A1(N5363), .A2(N5364), .ZN(n15554));
    NOR2X1 U2683 (.A1(N5365), .A2(N5366), .ZN(n15555));
    NOR2X1 U2684 (.A1(N5367), .A2(N5368), .ZN(N15556));
    NOR2X1 U2685 (.A1(N5369), .A2(N5370), .ZN(n15557));
    NOR2X1 U2686 (.A1(N5371), .A2(N5372), .ZN(n15558));
    NANDX1 U2687 (.A1(N5373), .A2(N5374), .ZN(n15559));
    NOR2X1 U2688 (.A1(N5375), .A2(N5376), .ZN(n15560));
    NOR2X1 U2689 (.A1(N5377), .A2(N5378), .ZN(N15561));
    NANDX1 U2690 (.A1(N5379), .A2(N5380), .ZN(n15562));
    NOR2X1 U2691 (.A1(N5381), .A2(N5382), .ZN(n15563));
    NOR2X1 U2692 (.A1(N5383), .A2(N5384), .ZN(N15564));
    NOR2X1 U2693 (.A1(N5385), .A2(N5386), .ZN(n15565));
    NOR2X1 U2694 (.A1(N5387), .A2(N5388), .ZN(n15566));
    NOR2X1 U2695 (.A1(N5389), .A2(N5390), .ZN(n15567));
    NOR2X1 U2696 (.A1(N5391), .A2(N5392), .ZN(n15568));
    NOR2X1 U2697 (.A1(N5393), .A2(N5394), .ZN(n15569));
    NOR2X1 U2698 (.A1(N5395), .A2(N5396), .ZN(n15570));
    NANDX1 U2699 (.A1(N5397), .A2(N5398), .ZN(n15571));
    NOR2X1 U2700 (.A1(N5399), .A2(N5400), .ZN(N15572));
    NOR2X1 U2701 (.A1(N5401), .A2(N5402), .ZN(n15573));
    NANDX1 U2702 (.A1(N5403), .A2(N5404), .ZN(n15574));
    NANDX1 U2703 (.A1(N5405), .A2(N5406), .ZN(N15575));
    NOR2X1 U2704 (.A1(N5407), .A2(N5408), .ZN(n15576));
    NANDX1 U2705 (.A1(N5409), .A2(N5410), .ZN(n15577));
    NOR2X1 U2706 (.A1(N5411), .A2(N5412), .ZN(n15578));
    NANDX1 U2707 (.A1(N5413), .A2(N5414), .ZN(n15579));
    NANDX1 U2708 (.A1(N5415), .A2(N5416), .ZN(n15580));
    NOR2X1 U2709 (.A1(N5417), .A2(N5418), .ZN(n15581));
    NOR2X1 U2710 (.A1(N5419), .A2(N5420), .ZN(n15582));
    NANDX1 U2711 (.A1(N5421), .A2(N5422), .ZN(n15583));
    NANDX1 U2712 (.A1(N5423), .A2(N5424), .ZN(n15584));
    NANDX1 U2713 (.A1(N5425), .A2(N5426), .ZN(n15585));
    NANDX1 U2714 (.A1(N5427), .A2(N5428), .ZN(n15586));
    NANDX1 U2715 (.A1(N5429), .A2(N5430), .ZN(n15587));
    NOR2X1 U2716 (.A1(N5431), .A2(N5432), .ZN(n15588));
    NOR2X1 U2717 (.A1(N5433), .A2(N5434), .ZN(n15589));
    NANDX1 U2718 (.A1(N5435), .A2(N5436), .ZN(n15590));
    NOR2X1 U2719 (.A1(N5437), .A2(N5438), .ZN(N15591));
    NOR2X1 U2720 (.A1(N5439), .A2(N5440), .ZN(N15592));
    NOR2X1 U2721 (.A1(N5441), .A2(N5442), .ZN(n15593));
    NOR2X1 U2722 (.A1(N5443), .A2(N5444), .ZN(n15594));
    NANDX1 U2723 (.A1(N5445), .A2(N5446), .ZN(n15595));
    NANDX1 U2724 (.A1(N5447), .A2(N5448), .ZN(n15596));
    NANDX1 U2725 (.A1(N5449), .A2(N5450), .ZN(n15597));
    NANDX1 U2726 (.A1(N5451), .A2(N5452), .ZN(n15598));
    NANDX1 U2727 (.A1(N5453), .A2(N5454), .ZN(n15599));
    NANDX1 U2728 (.A1(N5455), .A2(N5456), .ZN(N15600));
    NANDX1 U2729 (.A1(N5457), .A2(N5458), .ZN(n15601));
    NOR2X1 U2730 (.A1(N5459), .A2(N5460), .ZN(n15602));
    NANDX1 U2731 (.A1(N5461), .A2(N5462), .ZN(n15603));
    NANDX1 U2732 (.A1(N5463), .A2(N5464), .ZN(n15604));
    NANDX1 U2733 (.A1(N5465), .A2(N5466), .ZN(n15605));
    NOR2X1 U2734 (.A1(N5467), .A2(N5468), .ZN(n15606));
    NOR2X1 U2735 (.A1(N5469), .A2(N5470), .ZN(n15607));
    NOR2X1 U2736 (.A1(N5471), .A2(N5472), .ZN(n15608));
    NOR2X1 U2737 (.A1(N5473), .A2(N5474), .ZN(n15609));
    NANDX1 U2738 (.A1(N5475), .A2(N5476), .ZN(n15610));
    NANDX1 U2739 (.A1(N5477), .A2(N5478), .ZN(n15611));
    NANDX1 U2740 (.A1(N5479), .A2(N5480), .ZN(n15612));
    NANDX1 U2741 (.A1(N5481), .A2(N5482), .ZN(n15613));
    NOR2X1 U2742 (.A1(N5483), .A2(N5484), .ZN(n15614));
    NOR2X1 U2743 (.A1(N5485), .A2(N5486), .ZN(n15615));
    NANDX1 U2744 (.A1(N5487), .A2(N5488), .ZN(n15616));
    NOR2X1 U2745 (.A1(N5489), .A2(N5490), .ZN(n15617));
    NOR2X1 U2746 (.A1(N5491), .A2(N5492), .ZN(n15618));
    NANDX1 U2747 (.A1(N5493), .A2(N5494), .ZN(n15619));
    NOR2X1 U2748 (.A1(N5495), .A2(N5496), .ZN(n15620));
    NANDX1 U2749 (.A1(N5497), .A2(N5498), .ZN(n15621));
    NANDX1 U2750 (.A1(N5499), .A2(N5500), .ZN(N15622));
    NOR2X1 U2751 (.A1(N5501), .A2(N5502), .ZN(n15623));
    NANDX1 U2752 (.A1(N5503), .A2(N5504), .ZN(n15624));
    NANDX1 U2753 (.A1(N5505), .A2(N5506), .ZN(n15625));
    NANDX1 U2754 (.A1(N5507), .A2(N5508), .ZN(n15626));
    NOR2X1 U2755 (.A1(N5509), .A2(N5510), .ZN(n15627));
    NOR2X1 U2756 (.A1(N5511), .A2(N5512), .ZN(n15628));
    NANDX1 U2757 (.A1(N5513), .A2(N5514), .ZN(n15629));
    NOR2X1 U2758 (.A1(N5515), .A2(N5516), .ZN(n15630));
    NANDX1 U2759 (.A1(N5517), .A2(N5518), .ZN(n15631));
    NOR2X1 U2760 (.A1(N5519), .A2(N5520), .ZN(n15632));
    NOR2X1 U2761 (.A1(N5521), .A2(N5522), .ZN(n15633));
    NANDX1 U2762 (.A1(N5523), .A2(N5524), .ZN(n15634));
    NOR2X1 U2763 (.A1(N5525), .A2(N5526), .ZN(n15635));
    NOR2X1 U2764 (.A1(N5527), .A2(N5528), .ZN(n15636));
    NANDX1 U2765 (.A1(N5529), .A2(N5530), .ZN(n15637));
    NOR2X1 U2766 (.A1(N5531), .A2(N5532), .ZN(N15638));
    NOR2X1 U2767 (.A1(N5533), .A2(N5534), .ZN(n15639));
    NOR2X1 U2768 (.A1(N5535), .A2(N5536), .ZN(n15640));
    NANDX1 U2769 (.A1(N5537), .A2(N5538), .ZN(n15641));
    NOR2X1 U2770 (.A1(N5539), .A2(N5540), .ZN(n15642));
    NANDX1 U2771 (.A1(N5541), .A2(N5542), .ZN(N15643));
    NANDX1 U2772 (.A1(N5543), .A2(N5544), .ZN(n15644));
    NOR2X1 U2773 (.A1(N5545), .A2(N5546), .ZN(n15645));
    NANDX1 U2774 (.A1(N5547), .A2(N5548), .ZN(N15646));
    NOR2X1 U2775 (.A1(N5549), .A2(N5550), .ZN(n15647));
    NOR2X1 U2776 (.A1(N5551), .A2(N5552), .ZN(n15648));
    NANDX1 U2777 (.A1(N5553), .A2(N5554), .ZN(n15649));
    NANDX1 U2778 (.A1(N5555), .A2(N5556), .ZN(n15650));
    NOR2X1 U2779 (.A1(N5557), .A2(N5558), .ZN(n15651));
    NOR2X1 U2780 (.A1(N5559), .A2(N5560), .ZN(n15652));
    NOR2X1 U2781 (.A1(N5561), .A2(N5562), .ZN(N15653));
    NANDX1 U2782 (.A1(N5563), .A2(N5564), .ZN(n15654));
    NOR2X1 U2783 (.A1(N5565), .A2(N5566), .ZN(n15655));
    NANDX1 U2784 (.A1(N5567), .A2(N5568), .ZN(n15656));
    NOR2X1 U2785 (.A1(N5569), .A2(N5570), .ZN(n15657));
    NOR2X1 U2786 (.A1(N5571), .A2(N5572), .ZN(n15658));
    NOR2X1 U2787 (.A1(N5573), .A2(N5574), .ZN(n15659));
    NANDX1 U2788 (.A1(N5575), .A2(N5576), .ZN(N15660));
    NOR2X1 U2789 (.A1(N5577), .A2(N5578), .ZN(n15661));
    NANDX1 U2790 (.A1(N5579), .A2(N5580), .ZN(n15662));
    NOR2X1 U2791 (.A1(N5581), .A2(N5582), .ZN(n15663));
    NANDX1 U2792 (.A1(N5583), .A2(N5584), .ZN(N15664));
    NOR2X1 U2793 (.A1(N5585), .A2(N5586), .ZN(n15665));
    NOR2X1 U2794 (.A1(N5587), .A2(N5588), .ZN(n15666));
    NANDX1 U2795 (.A1(N5589), .A2(N5590), .ZN(n15667));
    NOR2X1 U2796 (.A1(N5591), .A2(N5592), .ZN(n15668));
    NOR2X1 U2797 (.A1(N5593), .A2(N5594), .ZN(n15669));
    NANDX1 U2798 (.A1(N5595), .A2(N5596), .ZN(N15670));
    NOR2X1 U2799 (.A1(N5597), .A2(N5598), .ZN(n15671));
    NANDX1 U2800 (.A1(N5599), .A2(N5600), .ZN(n15672));
    NANDX1 U2801 (.A1(N5601), .A2(N5602), .ZN(N15673));
    NANDX1 U2802 (.A1(N5603), .A2(N5604), .ZN(n15674));
    NOR2X1 U2803 (.A1(N5605), .A2(N5606), .ZN(n15675));
    NOR2X1 U2804 (.A1(N5607), .A2(N5608), .ZN(n15676));
    NOR2X1 U2805 (.A1(N5609), .A2(N5610), .ZN(N15677));
    NOR2X1 U2806 (.A1(N5611), .A2(N5612), .ZN(N15678));
    NOR2X1 U2807 (.A1(N5613), .A2(N5614), .ZN(n15679));
    NOR2X1 U2808 (.A1(N5615), .A2(N5616), .ZN(N15680));
    NANDX1 U2809 (.A1(N5617), .A2(N5618), .ZN(n15681));
    NANDX1 U2810 (.A1(N5619), .A2(N5620), .ZN(n15682));
    NOR2X1 U2811 (.A1(N5621), .A2(N5622), .ZN(n15683));
    NANDX1 U2812 (.A1(N5623), .A2(N5624), .ZN(n15684));
    NOR2X1 U2813 (.A1(N5625), .A2(N5626), .ZN(n15685));
    NOR2X1 U2814 (.A1(N5627), .A2(N5628), .ZN(n15686));
    NANDX1 U2815 (.A1(N5629), .A2(N5630), .ZN(n15687));
    NOR2X1 U2816 (.A1(N5631), .A2(N5632), .ZN(n15688));
    NANDX1 U2817 (.A1(N5633), .A2(N5634), .ZN(n15689));
    NANDX1 U2818 (.A1(N5635), .A2(N5636), .ZN(n15690));
    NOR2X1 U2819 (.A1(N5637), .A2(N5638), .ZN(N15691));
    NANDX1 U2820 (.A1(N5639), .A2(N5640), .ZN(n15692));
    NOR2X1 U2821 (.A1(N5641), .A2(N5642), .ZN(N15693));
    NOR2X1 U2822 (.A1(N5643), .A2(N5644), .ZN(n15694));
    NOR2X1 U2823 (.A1(N5645), .A2(N5646), .ZN(n15695));
    NANDX1 U2824 (.A1(N5647), .A2(N5648), .ZN(n15696));
    NOR2X1 U2825 (.A1(N5649), .A2(N5650), .ZN(n15697));
    NANDX1 U2826 (.A1(N5651), .A2(N5652), .ZN(n15698));
    NANDX1 U2827 (.A1(N5653), .A2(N5654), .ZN(n15699));
    NOR2X1 U2828 (.A1(N5655), .A2(N5656), .ZN(n15700));
    NANDX1 U2829 (.A1(N5657), .A2(N5658), .ZN(n15701));
    NANDX1 U2830 (.A1(N5659), .A2(N5660), .ZN(n15702));
    NANDX1 U2831 (.A1(N5661), .A2(N5662), .ZN(n15703));
    NOR2X1 U2832 (.A1(N5663), .A2(N5664), .ZN(n15704));
    NOR2X1 U2833 (.A1(N5665), .A2(N5666), .ZN(N15705));
    NOR2X1 U2834 (.A1(N5667), .A2(N5668), .ZN(n15706));
    NOR2X1 U2835 (.A1(N5669), .A2(N5670), .ZN(n15707));
    NOR2X1 U2836 (.A1(N5671), .A2(N5672), .ZN(N15708));
    NOR2X1 U2837 (.A1(N5673), .A2(N5674), .ZN(N15709));
    NANDX1 U2838 (.A1(N5675), .A2(N5676), .ZN(n15710));
    NOR2X1 U2839 (.A1(N5677), .A2(N5678), .ZN(N15711));
    NOR2X1 U2840 (.A1(N5679), .A2(N5680), .ZN(n15712));
    NOR2X1 U2841 (.A1(N5681), .A2(N5682), .ZN(n15713));
    NANDX1 U2842 (.A1(N5683), .A2(N5684), .ZN(n15714));
    NANDX1 U2843 (.A1(N5685), .A2(N5686), .ZN(N15715));
    NOR2X1 U2844 (.A1(N5687), .A2(N5688), .ZN(n15716));
    NANDX1 U2845 (.A1(N5689), .A2(N5690), .ZN(n15717));
    NOR2X1 U2846 (.A1(N5691), .A2(N5692), .ZN(n15718));
    NOR2X1 U2847 (.A1(N5693), .A2(N5694), .ZN(N15719));
    NOR2X1 U2848 (.A1(N5695), .A2(N5696), .ZN(n15720));
    NANDX1 U2849 (.A1(N5697), .A2(N5698), .ZN(n15721));
    NOR2X1 U2850 (.A1(N5699), .A2(N5700), .ZN(N15722));
    NOR2X1 U2851 (.A1(N5701), .A2(N5702), .ZN(n15723));
    NOR2X1 U2852 (.A1(N5703), .A2(N5704), .ZN(N15724));
    NOR2X1 U2853 (.A1(N5705), .A2(N5706), .ZN(n15725));
    NOR2X1 U2854 (.A1(N5707), .A2(N5708), .ZN(n15726));
    NANDX1 U2855 (.A1(N5709), .A2(N5710), .ZN(n15727));
    NOR2X1 U2856 (.A1(N5711), .A2(N5712), .ZN(n15728));
    NOR2X1 U2857 (.A1(N5713), .A2(N5714), .ZN(n15729));
    NOR2X1 U2858 (.A1(N5715), .A2(N5716), .ZN(n15730));
    NOR2X1 U2859 (.A1(N5717), .A2(N5718), .ZN(n15731));
    NANDX1 U2860 (.A1(N5719), .A2(N5720), .ZN(n15732));
    NANDX1 U2861 (.A1(N5721), .A2(N5722), .ZN(n15733));
    NOR2X1 U2862 (.A1(N5723), .A2(N5724), .ZN(n15734));
    NANDX1 U2863 (.A1(N5725), .A2(N5726), .ZN(n15735));
    NANDX1 U2864 (.A1(N5727), .A2(N5728), .ZN(n15736));
    NOR2X1 U2865 (.A1(N5729), .A2(N5730), .ZN(n15737));
    NOR2X1 U2866 (.A1(N5731), .A2(N5732), .ZN(N15738));
    NANDX1 U2867 (.A1(N5733), .A2(N5734), .ZN(n15739));
    NOR2X1 U2868 (.A1(N5735), .A2(N5736), .ZN(N15740));
    NANDX1 U2869 (.A1(N5737), .A2(N5738), .ZN(N15741));
    NOR2X1 U2870 (.A1(N5739), .A2(N5740), .ZN(n15742));
    NOR2X1 U2871 (.A1(N5741), .A2(N5742), .ZN(n15743));
    NANDX1 U2872 (.A1(N5743), .A2(N5744), .ZN(n15744));
    NANDX1 U2873 (.A1(N5745), .A2(N5746), .ZN(n15745));
    NOR2X1 U2874 (.A1(N5747), .A2(N5748), .ZN(n15746));
    NANDX1 U2875 (.A1(N5749), .A2(N5750), .ZN(n15747));
    NOR2X1 U2876 (.A1(N5751), .A2(N5752), .ZN(N15748));
    NOR2X1 U2877 (.A1(N5753), .A2(N5754), .ZN(n15749));
    NANDX1 U2878 (.A1(N5755), .A2(N5756), .ZN(n15750));
    NANDX1 U2879 (.A1(N5757), .A2(N5758), .ZN(n15751));
    NOR2X1 U2880 (.A1(N5759), .A2(N5760), .ZN(n15752));
    NOR2X1 U2881 (.A1(N5761), .A2(N5762), .ZN(n15753));
    NANDX1 U2882 (.A1(N5763), .A2(N5764), .ZN(n15754));
    NOR2X1 U2883 (.A1(N5765), .A2(N5766), .ZN(n15755));
    NOR2X1 U2884 (.A1(N5767), .A2(N5768), .ZN(N15756));
    NANDX1 U2885 (.A1(N5769), .A2(N5770), .ZN(n15757));
    NANDX1 U2886 (.A1(N5771), .A2(N5772), .ZN(n15758));
    NANDX1 U2887 (.A1(N5773), .A2(N5774), .ZN(n15759));
    NANDX1 U2888 (.A1(N5775), .A2(N5776), .ZN(n15760));
    NANDX1 U2889 (.A1(N5777), .A2(N5778), .ZN(N15761));
    NANDX1 U2890 (.A1(N5779), .A2(N5780), .ZN(n15762));
    NOR2X1 U2891 (.A1(N5781), .A2(N5782), .ZN(n15763));
    NOR2X1 U2892 (.A1(N5783), .A2(N5784), .ZN(n15764));
    NANDX1 U2893 (.A1(N5785), .A2(N5786), .ZN(n15765));
    NOR2X1 U2894 (.A1(N5787), .A2(N5788), .ZN(N15766));
    NANDX1 U2895 (.A1(N5789), .A2(N5790), .ZN(n15767));
    NANDX1 U2896 (.A1(N5791), .A2(N5792), .ZN(n15768));
    NOR2X1 U2897 (.A1(N5793), .A2(N5794), .ZN(n15769));
    NOR2X1 U2898 (.A1(N5795), .A2(N5796), .ZN(n15770));
    NOR2X1 U2899 (.A1(N5797), .A2(N5798), .ZN(n15771));
    NANDX1 U2900 (.A1(N5799), .A2(N5800), .ZN(n15772));
    NOR2X1 U2901 (.A1(N5801), .A2(N5802), .ZN(n15773));
    NOR2X1 U2902 (.A1(N5803), .A2(N5804), .ZN(N15774));
    NOR2X1 U2903 (.A1(N5805), .A2(N5806), .ZN(n15775));
    NANDX1 U2904 (.A1(N5807), .A2(N5808), .ZN(n15776));
    NOR2X1 U2905 (.A1(N5809), .A2(N5810), .ZN(n15777));
    NANDX1 U2906 (.A1(N5811), .A2(N5812), .ZN(n15778));
    NOR2X1 U2907 (.A1(N5813), .A2(N5814), .ZN(n15779));
    NANDX1 U2908 (.A1(N5815), .A2(N5816), .ZN(n15780));
    NOR2X1 U2909 (.A1(N5817), .A2(N5818), .ZN(n15781));
    NANDX1 U2910 (.A1(N5819), .A2(N5820), .ZN(n15782));
    NANDX1 U2911 (.A1(N5821), .A2(N5822), .ZN(n15783));
    NOR2X1 U2912 (.A1(N5823), .A2(N5824), .ZN(n15784));
    NOR2X1 U2913 (.A1(N5825), .A2(N5826), .ZN(n15785));
    NANDX1 U2914 (.A1(N5827), .A2(N5828), .ZN(n15786));
    NANDX1 U2915 (.A1(N5829), .A2(N5830), .ZN(n15787));
    NANDX1 U2916 (.A1(N5831), .A2(N5832), .ZN(N15788));
    NOR2X1 U2917 (.A1(N5833), .A2(N5834), .ZN(n15789));
    NOR2X1 U2918 (.A1(N5835), .A2(N5836), .ZN(n15790));
    NANDX1 U2919 (.A1(N5837), .A2(N5838), .ZN(n15791));
    NANDX1 U2920 (.A1(N5839), .A2(N5840), .ZN(n15792));
    NANDX1 U2921 (.A1(N5841), .A2(N5842), .ZN(N15793));
    NANDX1 U2922 (.A1(N5843), .A2(N5844), .ZN(n15794));
    NANDX1 U2923 (.A1(N5845), .A2(N5846), .ZN(N15795));
    NANDX1 U2924 (.A1(N5847), .A2(N5848), .ZN(n15796));
    NANDX1 U2925 (.A1(N5849), .A2(N5850), .ZN(n15797));
    NOR2X1 U2926 (.A1(N5851), .A2(N5852), .ZN(N15798));
    NOR2X1 U2927 (.A1(N5853), .A2(N5854), .ZN(N15799));
    NANDX1 U2928 (.A1(N5855), .A2(N5856), .ZN(n15800));
    NOR2X1 U2929 (.A1(N5857), .A2(N5858), .ZN(n15801));
    NOR2X1 U2930 (.A1(N5859), .A2(N5860), .ZN(n15802));
    NOR2X1 U2931 (.A1(N5861), .A2(N5862), .ZN(n15803));
    NANDX1 U2932 (.A1(N5863), .A2(N5864), .ZN(n15804));
    NANDX1 U2933 (.A1(N5865), .A2(N5866), .ZN(n15805));
    NOR2X1 U2934 (.A1(N5867), .A2(N5868), .ZN(n15806));
    NOR2X1 U2935 (.A1(N5869), .A2(N5870), .ZN(n15807));
    NANDX1 U2936 (.A1(N5871), .A2(N5872), .ZN(n15808));
    NANDX1 U2937 (.A1(N5873), .A2(N5874), .ZN(n15809));
    NOR2X1 U2938 (.A1(N5875), .A2(N5876), .ZN(n15810));
    NOR2X1 U2939 (.A1(N5877), .A2(N5878), .ZN(n15811));
    NOR2X1 U2940 (.A1(N5879), .A2(N5880), .ZN(n15812));
    NANDX1 U2941 (.A1(N5881), .A2(N5882), .ZN(n15813));
    NANDX1 U2942 (.A1(N5883), .A2(N5884), .ZN(n15814));
    NOR2X1 U2943 (.A1(N5885), .A2(N5886), .ZN(n15815));
    NANDX1 U2944 (.A1(N5887), .A2(N5888), .ZN(n15816));
    NOR2X1 U2945 (.A1(N5889), .A2(N5890), .ZN(n15817));
    NANDX1 U2946 (.A1(N5891), .A2(N5892), .ZN(N15818));
    NANDX1 U2947 (.A1(N5893), .A2(N5894), .ZN(N15819));
    NOR2X1 U2948 (.A1(N5895), .A2(N5896), .ZN(n15820));
    NANDX1 U2949 (.A1(N5897), .A2(N5898), .ZN(n15821));
    NOR2X1 U2950 (.A1(N5899), .A2(N5900), .ZN(n15822));
    NANDX1 U2951 (.A1(N5901), .A2(N5902), .ZN(N15823));
    NANDX1 U2952 (.A1(N5903), .A2(N5904), .ZN(n15824));
    NANDX1 U2953 (.A1(N5905), .A2(N5906), .ZN(n15825));
    NOR2X1 U2954 (.A1(N5907), .A2(N5908), .ZN(n15826));
    NOR2X1 U2955 (.A1(N5909), .A2(N5910), .ZN(n15827));
    NANDX1 U2956 (.A1(N5911), .A2(N5912), .ZN(N15828));
    NOR2X1 U2957 (.A1(N5913), .A2(N5914), .ZN(n15829));
    NOR2X1 U2958 (.A1(N5915), .A2(N5916), .ZN(n15830));
    NOR2X1 U2959 (.A1(N5917), .A2(N5918), .ZN(N15831));
    NANDX1 U2960 (.A1(N5919), .A2(N5920), .ZN(n15832));
    NANDX1 U2961 (.A1(N5921), .A2(N5922), .ZN(n15833));
    NANDX1 U2962 (.A1(N5923), .A2(N5924), .ZN(n15834));
    NOR2X1 U2963 (.A1(N5925), .A2(N5926), .ZN(N15835));
    NOR2X1 U2964 (.A1(N5927), .A2(N5928), .ZN(N15836));
    NANDX1 U2965 (.A1(N5929), .A2(N5930), .ZN(N15837));
    NOR2X1 U2966 (.A1(N5931), .A2(N5932), .ZN(n15838));
    NANDX1 U2967 (.A1(N5933), .A2(N5934), .ZN(n15839));
    NANDX1 U2968 (.A1(N5935), .A2(N5936), .ZN(n15840));
    NANDX1 U2969 (.A1(N5937), .A2(N5938), .ZN(n15841));
    NOR2X1 U2970 (.A1(N5939), .A2(N5940), .ZN(n15842));
    NANDX1 U2971 (.A1(N5941), .A2(N5942), .ZN(n15843));
    NOR2X1 U2972 (.A1(N5943), .A2(N5944), .ZN(N15844));
    NANDX1 U2973 (.A1(N5945), .A2(N5946), .ZN(n15845));
    NANDX1 U2974 (.A1(N5947), .A2(N5948), .ZN(n15846));
    NOR2X1 U2975 (.A1(N5949), .A2(N5950), .ZN(N15847));
    NOR2X1 U2976 (.A1(N5951), .A2(N5952), .ZN(n15848));
    NANDX1 U2977 (.A1(N5953), .A2(N5954), .ZN(n15849));
    NANDX1 U2978 (.A1(N5955), .A2(N5956), .ZN(n15850));
    NOR2X1 U2979 (.A1(N5957), .A2(N5958), .ZN(n15851));
    NOR2X1 U2980 (.A1(N5959), .A2(N5960), .ZN(N15852));
    NANDX1 U2981 (.A1(N5961), .A2(N5962), .ZN(n15853));
    NOR2X1 U2982 (.A1(N5963), .A2(N5964), .ZN(N15854));
    NANDX1 U2983 (.A1(N5965), .A2(N5966), .ZN(n15855));
    NOR2X1 U2984 (.A1(N5967), .A2(N5968), .ZN(n15856));
    NOR2X1 U2985 (.A1(N5969), .A2(N5970), .ZN(n15857));
    NANDX1 U2986 (.A1(N5971), .A2(N5972), .ZN(n15858));
    NANDX1 U2987 (.A1(N5973), .A2(N5974), .ZN(n15859));
    NANDX1 U2988 (.A1(N5975), .A2(N5976), .ZN(n15860));
    NOR2X1 U2989 (.A1(N5977), .A2(N5978), .ZN(n15861));
    NOR2X1 U2990 (.A1(N5979), .A2(N5980), .ZN(n15862));
    NOR2X1 U2991 (.A1(N5981), .A2(N5982), .ZN(n15863));
    NANDX1 U2992 (.A1(N5983), .A2(N5984), .ZN(n15864));
    NANDX1 U2993 (.A1(N5985), .A2(N5986), .ZN(n15865));
    NOR2X1 U2994 (.A1(N5987), .A2(N5988), .ZN(n15866));
    NANDX1 U2995 (.A1(N5989), .A2(N5990), .ZN(n15867));
    NOR2X1 U2996 (.A1(N5991), .A2(N5992), .ZN(n15868));
    NOR2X1 U2997 (.A1(N5993), .A2(N5994), .ZN(n15869));
    NOR2X1 U2998 (.A1(N5995), .A2(N5996), .ZN(n15870));
    NANDX1 U2999 (.A1(N5997), .A2(N5998), .ZN(n15871));
    NANDX1 U3000 (.A1(N5999), .A2(N6000), .ZN(n15872));
    NOR2X1 U3001 (.A1(N6001), .A2(N6002), .ZN(n15873));
    NOR2X1 U3002 (.A1(N6003), .A2(N6004), .ZN(n15874));
    NOR2X1 U3003 (.A1(N6005), .A2(N6006), .ZN(n15875));
    NOR2X1 U3004 (.A1(N6007), .A2(N6008), .ZN(n15876));
    NOR2X1 U3005 (.A1(N6009), .A2(N6010), .ZN(n15877));
    NOR2X1 U3006 (.A1(N6011), .A2(N6012), .ZN(N15878));
    NOR2X1 U3007 (.A1(N6013), .A2(N6014), .ZN(n15879));
    NANDX1 U3008 (.A1(N6015), .A2(N6016), .ZN(n15880));
    NANDX1 U3009 (.A1(N6017), .A2(N6018), .ZN(n15881));
    NOR2X1 U3010 (.A1(N6019), .A2(N6020), .ZN(n15882));
    NANDX1 U3011 (.A1(N6021), .A2(N6022), .ZN(n15883));
    NOR2X1 U3012 (.A1(N6023), .A2(N6024), .ZN(n15884));
    NOR2X1 U3013 (.A1(N6025), .A2(N6026), .ZN(n15885));
    NANDX1 U3014 (.A1(N6027), .A2(N6028), .ZN(n15886));
    NOR2X1 U3015 (.A1(N6029), .A2(N6030), .ZN(n15887));
    NANDX1 U3016 (.A1(N6031), .A2(N6032), .ZN(n15888));
    NOR2X1 U3017 (.A1(N6033), .A2(N6034), .ZN(N15889));
    NOR2X1 U3018 (.A1(N6035), .A2(N6036), .ZN(N15890));
    NOR2X1 U3019 (.A1(N6037), .A2(N6038), .ZN(n15891));
    NOR2X1 U3020 (.A1(N6039), .A2(N6040), .ZN(n15892));
    NOR2X1 U3021 (.A1(N6041), .A2(N6042), .ZN(N15893));
    NOR2X1 U3022 (.A1(N6043), .A2(N6044), .ZN(n15894));
    NANDX1 U3023 (.A1(N6045), .A2(N6046), .ZN(n15895));
    NANDX1 U3024 (.A1(N6047), .A2(N6048), .ZN(n15896));
    NOR2X1 U3025 (.A1(N6049), .A2(N6050), .ZN(n15897));
    NOR2X1 U3026 (.A1(N6051), .A2(N6052), .ZN(n15898));
    NANDX1 U3027 (.A1(N6053), .A2(N6054), .ZN(n15899));
    NOR2X1 U3028 (.A1(N6055), .A2(N6056), .ZN(n15900));
    NANDX1 U3029 (.A1(N6057), .A2(N6058), .ZN(n15901));
    NANDX1 U3030 (.A1(N6059), .A2(N6060), .ZN(n15902));
    NOR2X1 U3031 (.A1(N6061), .A2(N6062), .ZN(n15903));
    NANDX1 U3032 (.A1(N6063), .A2(N6064), .ZN(n15904));
    NANDX1 U3033 (.A1(N6065), .A2(N6066), .ZN(n15905));
    NOR2X1 U3034 (.A1(N6067), .A2(N6068), .ZN(n15906));
    NANDX1 U3035 (.A1(N6069), .A2(N6070), .ZN(n15907));
    NANDX1 U3036 (.A1(N6071), .A2(N6072), .ZN(N15908));
    NOR2X1 U3037 (.A1(N6073), .A2(N6074), .ZN(n15909));
    NANDX1 U3038 (.A1(N6075), .A2(N6076), .ZN(N15910));
    NOR2X1 U3039 (.A1(N6077), .A2(N6078), .ZN(n15911));
    NANDX1 U3040 (.A1(N6079), .A2(N6080), .ZN(n15912));
    NOR2X1 U3041 (.A1(N6081), .A2(N6082), .ZN(n15913));
    NOR2X1 U3042 (.A1(N6083), .A2(N6084), .ZN(n15914));
    NANDX1 U3043 (.A1(N6085), .A2(N6086), .ZN(n15915));
    NOR2X1 U3044 (.A1(N6087), .A2(N6088), .ZN(N15916));
    NANDX1 U3045 (.A1(N6089), .A2(N6090), .ZN(n15917));
    NANDX1 U3046 (.A1(N6091), .A2(N6092), .ZN(n15918));
    NANDX1 U3047 (.A1(N6093), .A2(N6094), .ZN(n15919));
    NANDX1 U3048 (.A1(N6095), .A2(N6096), .ZN(n15920));
    NANDX1 U3049 (.A1(N6097), .A2(N6098), .ZN(n15921));
    NANDX1 U3050 (.A1(N6099), .A2(N6100), .ZN(n15922));
    NOR2X1 U3051 (.A1(N6101), .A2(N6102), .ZN(n15923));
    NANDX1 U3052 (.A1(N6103), .A2(N6104), .ZN(n15924));
    NANDX1 U3053 (.A1(N6105), .A2(N6106), .ZN(n15925));
    NANDX1 U3054 (.A1(N6107), .A2(N6108), .ZN(n15926));
    NOR2X1 U3055 (.A1(N6109), .A2(N6110), .ZN(n15927));
    NANDX1 U3056 (.A1(N6111), .A2(N6112), .ZN(n15928));
    NOR2X1 U3057 (.A1(N6113), .A2(N6114), .ZN(N15929));
    NOR2X1 U3058 (.A1(N6115), .A2(N6116), .ZN(n15930));
    NOR2X1 U3059 (.A1(N6117), .A2(N6118), .ZN(n15931));
    NANDX1 U3060 (.A1(N6119), .A2(N6120), .ZN(n15932));
    NANDX1 U3061 (.A1(N6121), .A2(N6122), .ZN(n15933));
    NOR2X1 U3062 (.A1(N6123), .A2(N6124), .ZN(N15934));
    NOR2X1 U3063 (.A1(N6125), .A2(N6126), .ZN(n15935));
    NOR2X1 U3064 (.A1(N6127), .A2(N6128), .ZN(n15936));
    NOR2X1 U3065 (.A1(N6129), .A2(N6130), .ZN(n15937));
    NOR2X1 U3066 (.A1(N6131), .A2(N6132), .ZN(n15938));
    NOR2X1 U3067 (.A1(N6133), .A2(N6134), .ZN(n15939));
    NOR2X1 U3068 (.A1(N6135), .A2(N6136), .ZN(n15940));
    NANDX1 U3069 (.A1(N6137), .A2(N6138), .ZN(n15941));
    NOR2X1 U3070 (.A1(N6139), .A2(N6140), .ZN(n15942));
    NANDX1 U3071 (.A1(N6141), .A2(N6142), .ZN(n15943));
    NANDX1 U3072 (.A1(N6143), .A2(N6144), .ZN(n15944));
    NOR2X1 U3073 (.A1(N6145), .A2(N6146), .ZN(n15945));
    NOR2X1 U3074 (.A1(N6147), .A2(N6148), .ZN(n15946));
    NOR2X1 U3075 (.A1(N6149), .A2(N6150), .ZN(n15947));
    NANDX1 U3076 (.A1(N6151), .A2(N6152), .ZN(N15948));
    NANDX1 U3077 (.A1(N6153), .A2(N6154), .ZN(n15949));
    NANDX1 U3078 (.A1(N6155), .A2(N6156), .ZN(n15950));
    NANDX1 U3079 (.A1(N6157), .A2(N6158), .ZN(N15951));
    NANDX1 U3080 (.A1(N6159), .A2(N6160), .ZN(n15952));
    NANDX1 U3081 (.A1(N6161), .A2(N6162), .ZN(n15953));
    NANDX1 U3082 (.A1(N6163), .A2(N6164), .ZN(n15954));
    NOR2X1 U3083 (.A1(N6165), .A2(N6166), .ZN(n15955));
    NOR2X1 U3084 (.A1(N6167), .A2(N6168), .ZN(n15956));
    NOR2X1 U3085 (.A1(N6169), .A2(N6170), .ZN(n15957));
    NANDX1 U3086 (.A1(N6171), .A2(N6172), .ZN(n15958));
    NOR2X1 U3087 (.A1(N6173), .A2(N6174), .ZN(n15959));
    NOR2X1 U3088 (.A1(N6175), .A2(N6176), .ZN(n15960));
    NANDX1 U3089 (.A1(N6177), .A2(N6178), .ZN(n15961));
    NOR2X1 U3090 (.A1(N6179), .A2(N6180), .ZN(n15962));
    NANDX1 U3091 (.A1(N6181), .A2(N6182), .ZN(N15963));
    NOR2X1 U3092 (.A1(N6183), .A2(N6184), .ZN(n15964));
    NOR2X1 U3093 (.A1(N6185), .A2(N6186), .ZN(n15965));
    NOR2X1 U3094 (.A1(N6187), .A2(N6188), .ZN(n15966));
    NOR2X1 U3095 (.A1(N6189), .A2(N6190), .ZN(n15967));
    NOR2X1 U3096 (.A1(N6191), .A2(N6192), .ZN(n15968));
    NOR2X1 U3097 (.A1(N6193), .A2(N6194), .ZN(N15969));
    NOR2X1 U3098 (.A1(N6195), .A2(N6196), .ZN(N15970));
    NOR2X1 U3099 (.A1(N6197), .A2(N6198), .ZN(n15971));
    NANDX1 U3100 (.A1(N6199), .A2(N6200), .ZN(n15972));
    NANDX1 U3101 (.A1(N6201), .A2(N6202), .ZN(n15973));
    NANDX1 U3102 (.A1(N6203), .A2(N6204), .ZN(n15974));
    NANDX1 U3103 (.A1(N6205), .A2(N6206), .ZN(N15975));
    NANDX1 U3104 (.A1(N6207), .A2(N6208), .ZN(n15976));
    NANDX1 U3105 (.A1(N6209), .A2(N6210), .ZN(n15977));
    NANDX1 U3106 (.A1(N6211), .A2(N6212), .ZN(n15978));
    NANDX1 U3107 (.A1(N6213), .A2(N6214), .ZN(n15979));
    NOR2X1 U3108 (.A1(N6215), .A2(N6216), .ZN(n15980));
    NOR2X1 U3109 (.A1(N6217), .A2(N6218), .ZN(n15981));
    NOR2X1 U3110 (.A1(N6219), .A2(N6220), .ZN(n15982));
    NANDX1 U3111 (.A1(N6221), .A2(N6222), .ZN(n15983));
    NANDX1 U3112 (.A1(N6223), .A2(N6224), .ZN(N15984));
    NANDX1 U3113 (.A1(N6225), .A2(N6226), .ZN(n15985));
    NOR2X1 U3114 (.A1(N6227), .A2(N6228), .ZN(n15986));
    NOR2X1 U3115 (.A1(N6229), .A2(N6230), .ZN(n15987));
    NANDX1 U3116 (.A1(N6231), .A2(N6232), .ZN(n15988));
    NANDX1 U3117 (.A1(N6233), .A2(N6234), .ZN(n15989));
    NOR2X1 U3118 (.A1(N6235), .A2(N6236), .ZN(n15990));
    NOR2X1 U3119 (.A1(N6237), .A2(N6238), .ZN(N15991));
    NOR2X1 U3120 (.A1(N6239), .A2(N6240), .ZN(n15992));
    NOR2X1 U3121 (.A1(N6241), .A2(N6242), .ZN(n15993));
    NANDX1 U3122 (.A1(N6243), .A2(N6244), .ZN(n15994));
    NOR2X1 U3123 (.A1(N6245), .A2(N6246), .ZN(n15995));
    NOR2X1 U3124 (.A1(N6247), .A2(N6248), .ZN(n15996));
    NANDX1 U3125 (.A1(N6249), .A2(N6250), .ZN(n15997));
    NOR2X1 U3126 (.A1(N6251), .A2(N6252), .ZN(n15998));
    NOR2X1 U3127 (.A1(N6253), .A2(N6254), .ZN(n15999));
    NANDX1 U3128 (.A1(N6255), .A2(N6256), .ZN(n16000));
    NANDX1 U3129 (.A1(N6257), .A2(N6258), .ZN(n16001));
    NOR2X1 U3130 (.A1(N6259), .A2(N6260), .ZN(n16002));
    NANDX1 U3131 (.A1(N6261), .A2(N6262), .ZN(n16003));
    NOR2X1 U3132 (.A1(N6263), .A2(N6264), .ZN(n16004));
    NANDX1 U3133 (.A1(N6265), .A2(N6266), .ZN(n16005));
    NOR2X1 U3134 (.A1(N6267), .A2(N6268), .ZN(n16006));
    NANDX1 U3135 (.A1(N6269), .A2(N6270), .ZN(n16007));
    NOR2X1 U3136 (.A1(N6271), .A2(N6272), .ZN(N16008));
    NANDX1 U3137 (.A1(N6273), .A2(N6274), .ZN(N16009));
    NOR2X1 U3138 (.A1(N6275), .A2(N6276), .ZN(N16010));
    NOR2X1 U3139 (.A1(N6277), .A2(N6278), .ZN(n16011));
    NANDX1 U3140 (.A1(N6279), .A2(N6280), .ZN(N16012));
    NOR2X1 U3141 (.A1(N6281), .A2(N6282), .ZN(n16013));
    NOR2X1 U3142 (.A1(N6283), .A2(N6284), .ZN(N16014));
    NANDX1 U3143 (.A1(N6285), .A2(N6286), .ZN(n16015));
    NANDX1 U3144 (.A1(N6287), .A2(N6288), .ZN(n16016));
    NOR2X1 U3145 (.A1(N6289), .A2(N6290), .ZN(n16017));
    NANDX1 U3146 (.A1(N6291), .A2(N6292), .ZN(n16018));
    NANDX1 U3147 (.A1(N6293), .A2(N6294), .ZN(n16019));
    NANDX1 U3148 (.A1(N6295), .A2(N6296), .ZN(N16020));
    NANDX1 U3149 (.A1(N6297), .A2(N6298), .ZN(n16021));
    NANDX1 U3150 (.A1(N6299), .A2(N6300), .ZN(N16022));
    NANDX1 U3151 (.A1(N6301), .A2(N6302), .ZN(n16023));
    NANDX1 U3152 (.A1(N6303), .A2(N6304), .ZN(n16024));
    NOR2X1 U3153 (.A1(N6305), .A2(N6306), .ZN(n16025));
    NANDX1 U3154 (.A1(N6307), .A2(N6308), .ZN(N16026));
    NANDX1 U3155 (.A1(N6309), .A2(N6310), .ZN(n16027));
    NOR2X1 U3156 (.A1(N6311), .A2(N6312), .ZN(n16028));
    NANDX1 U3157 (.A1(N6313), .A2(N6314), .ZN(N16029));
    NANDX1 U3158 (.A1(N6315), .A2(N6316), .ZN(n16030));
    NANDX1 U3159 (.A1(N6317), .A2(N6318), .ZN(n16031));
    NOR2X1 U3160 (.A1(N6319), .A2(N6320), .ZN(n16032));
    NANDX1 U3161 (.A1(N6321), .A2(N6322), .ZN(n16033));
    NOR2X1 U3162 (.A1(N6323), .A2(N6324), .ZN(n16034));
    NOR2X1 U3163 (.A1(N6325), .A2(N6326), .ZN(N16035));
    NOR2X1 U3164 (.A1(N6327), .A2(N6328), .ZN(N16036));
    NOR2X1 U3165 (.A1(N6329), .A2(N6330), .ZN(n16037));
    NOR2X1 U3166 (.A1(N6331), .A2(N6332), .ZN(n16038));
    NOR2X1 U3167 (.A1(N6333), .A2(N6334), .ZN(n16039));
    NANDX1 U3168 (.A1(N6335), .A2(N6336), .ZN(n16040));
    NOR2X1 U3169 (.A1(N6337), .A2(N6338), .ZN(n16041));
    NOR2X1 U3170 (.A1(N6339), .A2(N6340), .ZN(N16042));
    NANDX1 U3171 (.A1(N6341), .A2(N6342), .ZN(n16043));
    NANDX1 U3172 (.A1(N6343), .A2(N6344), .ZN(n16044));
    NOR2X1 U3173 (.A1(N6345), .A2(N6346), .ZN(n16045));
    NOR2X1 U3174 (.A1(N6347), .A2(N6348), .ZN(N16046));
    NOR2X1 U3175 (.A1(N6349), .A2(N6350), .ZN(n16047));
    NOR2X1 U3176 (.A1(N6351), .A2(N6352), .ZN(n16048));
    NANDX1 U3177 (.A1(N6353), .A2(N6354), .ZN(n16049));
    NANDX1 U3178 (.A1(N6355), .A2(N6356), .ZN(N16050));
    NANDX1 U3179 (.A1(N6357), .A2(N6358), .ZN(n16051));
    NOR2X1 U3180 (.A1(N6359), .A2(N6360), .ZN(n16052));
    NOR2X1 U3181 (.A1(N6361), .A2(N6362), .ZN(n16053));
    NOR2X1 U3182 (.A1(N6363), .A2(N6364), .ZN(n16054));
    NANDX1 U3183 (.A1(N6365), .A2(N6366), .ZN(n16055));
    NANDX1 U3184 (.A1(N6367), .A2(N6368), .ZN(n16056));
    NANDX1 U3185 (.A1(N6369), .A2(N6370), .ZN(N16057));
    NOR2X1 U3186 (.A1(N6371), .A2(N6372), .ZN(N16058));
    NANDX1 U3187 (.A1(N6373), .A2(N6374), .ZN(n16059));
    NANDX1 U3188 (.A1(N6375), .A2(N6376), .ZN(N16060));
    NANDX1 U3189 (.A1(N6377), .A2(N6378), .ZN(n16061));
    NOR2X1 U3190 (.A1(N6379), .A2(N6380), .ZN(n16062));
    NANDX1 U3191 (.A1(N6381), .A2(N6382), .ZN(n16063));
    NOR2X1 U3192 (.A1(N6383), .A2(N6384), .ZN(n16064));
    NANDX1 U3193 (.A1(N6385), .A2(N6386), .ZN(n16065));
    NOR2X1 U3194 (.A1(N6387), .A2(N6388), .ZN(n16066));
    NOR2X1 U3195 (.A1(N6389), .A2(N6390), .ZN(n16067));
    NANDX1 U3196 (.A1(N6391), .A2(N6392), .ZN(N16068));
    NOR2X1 U3197 (.A1(N6393), .A2(N6394), .ZN(n16069));
    NOR2X1 U3198 (.A1(N6395), .A2(N6396), .ZN(n16070));
    NANDX1 U3199 (.A1(N6397), .A2(N6398), .ZN(n16071));
    NOR2X1 U3200 (.A1(N6399), .A2(N6400), .ZN(n16072));
    NOR2X1 U3201 (.A1(N6401), .A2(N6402), .ZN(n16073));
    NOR2X1 U3202 (.A1(N6403), .A2(N6404), .ZN(n16074));
    NANDX1 U3203 (.A1(N6405), .A2(N6406), .ZN(n16075));
    NANDX1 U3204 (.A1(N6407), .A2(N6408), .ZN(n16076));
    NOR2X1 U3205 (.A1(N6409), .A2(N6410), .ZN(n16077));
    NOR2X1 U3206 (.A1(N6411), .A2(N6412), .ZN(n16078));
    NANDX1 U3207 (.A1(N6413), .A2(N6414), .ZN(N16079));
    NANDX1 U3208 (.A1(N6415), .A2(N6416), .ZN(n16080));
    NANDX1 U3209 (.A1(N6417), .A2(N6418), .ZN(N16081));
    NANDX1 U3210 (.A1(N6419), .A2(N6420), .ZN(n16082));
    NANDX1 U3211 (.A1(N6421), .A2(N6422), .ZN(n16083));
    NOR2X1 U3212 (.A1(N6423), .A2(N6424), .ZN(n16084));
    NANDX1 U3213 (.A1(N6425), .A2(N6426), .ZN(n16085));
    NOR2X1 U3214 (.A1(N6427), .A2(N6428), .ZN(n16086));
    NANDX1 U3215 (.A1(N6429), .A2(N6430), .ZN(n16087));
    NANDX1 U3216 (.A1(N6431), .A2(N6432), .ZN(n16088));
    NOR2X1 U3217 (.A1(N6433), .A2(N6434), .ZN(n16089));
    NOR2X1 U3218 (.A1(N6435), .A2(N6436), .ZN(n16090));
    NOR2X1 U3219 (.A1(N6437), .A2(N6438), .ZN(n16091));
    NANDX1 U3220 (.A1(N6439), .A2(N6440), .ZN(n16092));
    NOR2X1 U3221 (.A1(N6441), .A2(N6442), .ZN(n16093));
    NANDX1 U3222 (.A1(N6443), .A2(N6444), .ZN(n16094));
    NANDX1 U3223 (.A1(N6445), .A2(N6446), .ZN(N16095));
    NANDX1 U3224 (.A1(N6447), .A2(N6448), .ZN(n16096));
    NANDX1 U3225 (.A1(N6449), .A2(N6450), .ZN(n16097));
    NANDX1 U3226 (.A1(N6451), .A2(N6452), .ZN(n16098));
    NANDX1 U3227 (.A1(N6453), .A2(N6454), .ZN(n16099));
    NANDX1 U3228 (.A1(N6455), .A2(N6456), .ZN(n16100));
    NANDX1 U3229 (.A1(N6457), .A2(N6458), .ZN(n16101));
    NOR2X1 U3230 (.A1(N6459), .A2(N6460), .ZN(n16102));
    NOR2X1 U3231 (.A1(N6461), .A2(N6462), .ZN(n16103));
    NANDX1 U3232 (.A1(N6463), .A2(N6464), .ZN(n16104));
    NOR2X1 U3233 (.A1(N6465), .A2(N6466), .ZN(n16105));
    NANDX1 U3234 (.A1(N6467), .A2(N6468), .ZN(n16106));
    NOR2X1 U3235 (.A1(N6469), .A2(N6470), .ZN(n16107));
    NOR2X1 U3236 (.A1(N6471), .A2(N6472), .ZN(n16108));
    NANDX1 U3237 (.A1(N6473), .A2(N6474), .ZN(n16109));
    NOR2X1 U3238 (.A1(N6475), .A2(N6476), .ZN(N16110));
    NANDX1 U3239 (.A1(N6477), .A2(N6478), .ZN(N16111));
    NANDX1 U3240 (.A1(N6479), .A2(N6480), .ZN(N16112));
    NANDX1 U3241 (.A1(N6481), .A2(N6482), .ZN(N16113));
    NOR2X1 U3242 (.A1(N6483), .A2(N6484), .ZN(n16114));
    NANDX1 U3243 (.A1(N6485), .A2(N6486), .ZN(n16115));
    NOR2X1 U3244 (.A1(N6487), .A2(N6488), .ZN(N16116));
    NOR2X1 U3245 (.A1(N6489), .A2(N6490), .ZN(n16117));
    NOR2X1 U3246 (.A1(N6491), .A2(N6492), .ZN(N16118));
    NANDX1 U3247 (.A1(N6493), .A2(N6494), .ZN(n16119));
    NOR2X1 U3248 (.A1(N6495), .A2(N6496), .ZN(n16120));
    NOR2X1 U3249 (.A1(N6497), .A2(N6498), .ZN(N16121));
    NANDX1 U3250 (.A1(N6499), .A2(N6500), .ZN(n16122));
    NANDX1 U3251 (.A1(N6501), .A2(N6502), .ZN(N16123));
    NOR2X1 U3252 (.A1(N6503), .A2(N6504), .ZN(n16124));
    NANDX1 U3253 (.A1(N6505), .A2(N6506), .ZN(n16125));
    NOR2X1 U3254 (.A1(N6507), .A2(N6508), .ZN(n16126));
    NOR2X1 U3255 (.A1(N6509), .A2(N6510), .ZN(n16127));
    NOR2X1 U3256 (.A1(N6511), .A2(N6512), .ZN(n16128));
    NANDX1 U3257 (.A1(N6513), .A2(N6514), .ZN(n16129));
    NANDX1 U3258 (.A1(N6515), .A2(N6516), .ZN(n16130));
    NOR2X1 U3259 (.A1(N6517), .A2(N6518), .ZN(n16131));
    NOR2X1 U3260 (.A1(N6519), .A2(N6520), .ZN(n16132));
    NANDX1 U3261 (.A1(N6521), .A2(N6522), .ZN(N16133));
    NOR2X1 U3262 (.A1(N6523), .A2(N6524), .ZN(n16134));
    NANDX1 U3263 (.A1(N6525), .A2(N6526), .ZN(n16135));
    NANDX1 U3264 (.A1(N6527), .A2(N6528), .ZN(n16136));
    NANDX1 U3265 (.A1(N6529), .A2(N6530), .ZN(n16137));
    NOR2X1 U3266 (.A1(N6531), .A2(N6532), .ZN(N16138));
    NANDX1 U3267 (.A1(N6533), .A2(N6534), .ZN(n16139));
    NANDX1 U3268 (.A1(N6535), .A2(N6536), .ZN(n16140));
    NOR2X1 U3269 (.A1(N6537), .A2(N6538), .ZN(n16141));
    NOR2X1 U3270 (.A1(N6539), .A2(N6540), .ZN(N16142));
    NOR2X1 U3271 (.A1(N6541), .A2(N6542), .ZN(n16143));
    NANDX1 U3272 (.A1(N6543), .A2(N6544), .ZN(n16144));
    NOR2X1 U3273 (.A1(N6545), .A2(N6546), .ZN(n16145));
    NANDX1 U3274 (.A1(N6547), .A2(N6548), .ZN(n16146));
    NANDX1 U3275 (.A1(N6549), .A2(N6550), .ZN(n16147));
    NOR2X1 U3276 (.A1(N6551), .A2(N6552), .ZN(n16148));
    NANDX1 U3277 (.A1(N6553), .A2(N6554), .ZN(n16149));
    NANDX1 U3278 (.A1(N6555), .A2(N6556), .ZN(n16150));
    NOR2X1 U3279 (.A1(N6557), .A2(N6558), .ZN(n16151));
    NANDX1 U3280 (.A1(N6559), .A2(N6560), .ZN(n16152));
    NOR2X1 U3281 (.A1(N6561), .A2(N6562), .ZN(n16153));
    NANDX1 U3282 (.A1(N6563), .A2(N6564), .ZN(N16154));
    NANDX1 U3283 (.A1(N6565), .A2(N6566), .ZN(n16155));
    NANDX1 U3284 (.A1(N6567), .A2(N6568), .ZN(n16156));
    NANDX1 U3285 (.A1(N6569), .A2(N6570), .ZN(n16157));
    NANDX1 U3286 (.A1(N6571), .A2(N6572), .ZN(n16158));
    NOR2X1 U3287 (.A1(N6573), .A2(N6574), .ZN(n16159));
    NOR2X1 U3288 (.A1(N6575), .A2(N6576), .ZN(N16160));
    NOR2X1 U3289 (.A1(N6577), .A2(N6578), .ZN(n16161));
    NOR2X1 U3290 (.A1(N6579), .A2(N6580), .ZN(n16162));
    NOR2X1 U3291 (.A1(N6581), .A2(N6582), .ZN(n16163));
    NANDX1 U3292 (.A1(N6583), .A2(N6584), .ZN(n16164));
    NOR2X1 U3293 (.A1(N6585), .A2(N6586), .ZN(n16165));
    NANDX1 U3294 (.A1(N6587), .A2(N6588), .ZN(n16166));
    NOR2X1 U3295 (.A1(N6589), .A2(N6590), .ZN(n16167));
    NANDX1 U3296 (.A1(N6591), .A2(N6592), .ZN(n16168));
    NANDX1 U3297 (.A1(N6593), .A2(N6594), .ZN(n16169));
    NANDX1 U3298 (.A1(N6595), .A2(N6596), .ZN(N16170));
    NOR2X1 U3299 (.A1(N6597), .A2(N6598), .ZN(n16171));
    NANDX1 U3300 (.A1(N6599), .A2(N6600), .ZN(n16172));
    NANDX1 U3301 (.A1(N6601), .A2(N6602), .ZN(n16173));
    NOR2X1 U3302 (.A1(N6603), .A2(N6604), .ZN(n16174));
    NOR2X1 U3303 (.A1(N6605), .A2(N6606), .ZN(n16175));
    NANDX1 U3304 (.A1(N6607), .A2(N6608), .ZN(n16176));
    NANDX1 U3305 (.A1(N6609), .A2(N6610), .ZN(N16177));
    NOR2X1 U3306 (.A1(N6611), .A2(N6612), .ZN(n16178));
    NANDX1 U3307 (.A1(N6613), .A2(N6614), .ZN(n16179));
    NOR2X1 U3308 (.A1(N6615), .A2(N6616), .ZN(n16180));
    NANDX1 U3309 (.A1(N6617), .A2(N6618), .ZN(n16181));
    NANDX1 U3310 (.A1(N6619), .A2(N6620), .ZN(n16182));
    NANDX1 U3311 (.A1(N6621), .A2(N6622), .ZN(N16183));
    NANDX1 U3312 (.A1(N6623), .A2(N6624), .ZN(n16184));
    NOR2X1 U3313 (.A1(N6625), .A2(N6626), .ZN(n16185));
    NANDX1 U3314 (.A1(N6627), .A2(N6628), .ZN(n16186));
    NANDX1 U3315 (.A1(N6629), .A2(N6630), .ZN(n16187));
    NANDX1 U3316 (.A1(N6631), .A2(N6632), .ZN(n16188));
    NOR2X1 U3317 (.A1(N6633), .A2(N6634), .ZN(n16189));
    NANDX1 U3318 (.A1(N6635), .A2(N6636), .ZN(n16190));
    NANDX1 U3319 (.A1(N6637), .A2(N6638), .ZN(N16191));
    NANDX1 U3320 (.A1(N6639), .A2(N6640), .ZN(n16192));
    NANDX1 U3321 (.A1(N6641), .A2(N6642), .ZN(N16193));
    NANDX1 U3322 (.A1(N6643), .A2(N6644), .ZN(n16194));
    NOR2X1 U3323 (.A1(N6645), .A2(N6646), .ZN(n16195));
    NANDX1 U3324 (.A1(N6647), .A2(N6648), .ZN(n16196));
    NANDX1 U3325 (.A1(N6649), .A2(N6650), .ZN(N16197));
    NANDX1 U3326 (.A1(N6651), .A2(N6652), .ZN(N16198));
    NOR2X1 U3327 (.A1(N6653), .A2(N6654), .ZN(n16199));
    NOR2X1 U3328 (.A1(N6655), .A2(N6656), .ZN(n16200));
    NOR2X1 U3329 (.A1(N6657), .A2(N6658), .ZN(N16201));
    NANDX1 U3330 (.A1(N6659), .A2(N6660), .ZN(N16202));
    NOR2X1 U3331 (.A1(N6661), .A2(N6662), .ZN(n16203));
    NOR2X1 U3332 (.A1(N6663), .A2(N6664), .ZN(n16204));
    NANDX1 U3333 (.A1(N6665), .A2(N6666), .ZN(n16205));
    NOR2X1 U3334 (.A1(N6667), .A2(N6668), .ZN(n16206));
    NANDX1 U3335 (.A1(N6669), .A2(N6670), .ZN(n16207));
    NANDX1 U3336 (.A1(N6671), .A2(N6672), .ZN(n16208));
    NOR2X1 U3337 (.A1(N6673), .A2(N6674), .ZN(n16209));
    NANDX1 U3338 (.A1(N6675), .A2(N6676), .ZN(N16210));
    NANDX1 U3339 (.A1(N6677), .A2(N6678), .ZN(n16211));
    NANDX1 U3340 (.A1(N6679), .A2(N6680), .ZN(n16212));
    NOR2X1 U3341 (.A1(N6681), .A2(N6682), .ZN(n16213));
    NANDX1 U3342 (.A1(N6683), .A2(N6684), .ZN(n16214));
    NANDX1 U3343 (.A1(N6685), .A2(N6686), .ZN(N16215));
    NANDX1 U3344 (.A1(N6687), .A2(N6688), .ZN(n16216));
    NOR2X1 U3345 (.A1(N6689), .A2(N6690), .ZN(n16217));
    NOR2X1 U3346 (.A1(N6691), .A2(N6692), .ZN(n16218));
    NOR2X1 U3347 (.A1(N6693), .A2(N6694), .ZN(n16219));
    NOR2X1 U3348 (.A1(N6695), .A2(N6696), .ZN(n16220));
    NANDX1 U3349 (.A1(N6697), .A2(N6698), .ZN(n16221));
    NOR2X1 U3350 (.A1(N6699), .A2(N6700), .ZN(n16222));
    NANDX1 U3351 (.A1(N6701), .A2(N6702), .ZN(n16223));
    NOR2X1 U3352 (.A1(N6703), .A2(N6704), .ZN(n16224));
    NANDX1 U3353 (.A1(N6705), .A2(N6706), .ZN(n16225));
    NOR2X1 U3354 (.A1(N6707), .A2(N6708), .ZN(n16226));
    NANDX1 U3355 (.A1(N6709), .A2(N6710), .ZN(n16227));
    NOR2X1 U3356 (.A1(N6711), .A2(N6712), .ZN(n16228));
    NANDX1 U3357 (.A1(N6713), .A2(N6714), .ZN(n16229));
    NANDX1 U3358 (.A1(N6715), .A2(N6716), .ZN(n16230));
    NANDX1 U3359 (.A1(N6717), .A2(N6718), .ZN(N16231));
    NANDX1 U3360 (.A1(N6719), .A2(N6720), .ZN(n16232));
    NOR2X1 U3361 (.A1(N6721), .A2(N6722), .ZN(N16233));
    NANDX1 U3362 (.A1(N6723), .A2(N6724), .ZN(n16234));
    NANDX1 U3363 (.A1(N6725), .A2(N6726), .ZN(n16235));
    NOR2X1 U3364 (.A1(N6727), .A2(N6728), .ZN(n16236));
    NANDX1 U3365 (.A1(N6729), .A2(N6730), .ZN(n16237));
    NANDX1 U3366 (.A1(N6731), .A2(N6732), .ZN(n16238));
    NANDX1 U3367 (.A1(N6733), .A2(N6734), .ZN(n16239));
    NOR2X1 U3368 (.A1(N6735), .A2(N6736), .ZN(n16240));
    NOR2X1 U3369 (.A1(N6737), .A2(N6738), .ZN(n16241));
    NOR2X1 U3370 (.A1(N6739), .A2(N6740), .ZN(n16242));
    NANDX1 U3371 (.A1(N6741), .A2(N6742), .ZN(n16243));
    NOR2X1 U3372 (.A1(N6743), .A2(N6744), .ZN(n16244));
    NANDX1 U3373 (.A1(N6745), .A2(N6746), .ZN(n16245));
    NOR2X1 U3374 (.A1(N6747), .A2(N6748), .ZN(n16246));
    NANDX1 U3375 (.A1(N6749), .A2(N6750), .ZN(n16247));
    NANDX1 U3376 (.A1(N6751), .A2(N6752), .ZN(n16248));
    NOR2X1 U3377 (.A1(N6753), .A2(N6754), .ZN(n16249));
    NOR2X1 U3378 (.A1(N6755), .A2(N6756), .ZN(n16250));
    NOR2X1 U3379 (.A1(N6757), .A2(N6758), .ZN(n16251));
    NANDX1 U3380 (.A1(N6759), .A2(N6760), .ZN(n16252));
    NOR2X1 U3381 (.A1(N6761), .A2(N6762), .ZN(n16253));
    NANDX1 U3382 (.A1(N6763), .A2(N6764), .ZN(n16254));
    NANDX1 U3383 (.A1(N6765), .A2(N6766), .ZN(N16255));
    NANDX1 U3384 (.A1(N6767), .A2(N6768), .ZN(N16256));
    NANDX1 U3385 (.A1(N6769), .A2(N6770), .ZN(n16257));
    NOR2X1 U3386 (.A1(N6771), .A2(N6772), .ZN(n16258));
    NOR2X1 U3387 (.A1(N6773), .A2(N6774), .ZN(n16259));
    NOR2X1 U3388 (.A1(N6775), .A2(N6776), .ZN(n16260));
    NOR2X1 U3389 (.A1(N6777), .A2(N6778), .ZN(n16261));
    NANDX1 U3390 (.A1(N6779), .A2(N6780), .ZN(n16262));
    NOR2X1 U3391 (.A1(N6781), .A2(N6782), .ZN(n16263));
    NOR2X1 U3392 (.A1(N6783), .A2(N6784), .ZN(n16264));
    NOR2X1 U3393 (.A1(N6785), .A2(N6786), .ZN(n16265));
    NANDX1 U3394 (.A1(N6787), .A2(N6788), .ZN(N16266));
    NOR2X1 U3395 (.A1(N6789), .A2(N6790), .ZN(n16267));
    NANDX1 U3396 (.A1(N6791), .A2(N6792), .ZN(n16268));
    NOR2X1 U3397 (.A1(N6793), .A2(N6794), .ZN(n16269));
    NANDX1 U3398 (.A1(N6795), .A2(N6796), .ZN(n16270));
    NANDX1 U3399 (.A1(N6797), .A2(N6798), .ZN(n16271));
    NOR2X1 U3400 (.A1(N6799), .A2(N6800), .ZN(n16272));
    NOR2X1 U3401 (.A1(N6801), .A2(N6802), .ZN(n16273));
    NANDX1 U3402 (.A1(N6803), .A2(N6804), .ZN(N16274));
    NANDX1 U3403 (.A1(N6805), .A2(N6806), .ZN(n16275));
    NANDX1 U3404 (.A1(N6807), .A2(N6808), .ZN(n16276));
    NANDX1 U3405 (.A1(N6809), .A2(N6810), .ZN(n16277));
    NOR2X1 U3406 (.A1(N6811), .A2(N6812), .ZN(N16278));
    NANDX1 U3407 (.A1(N6813), .A2(N6814), .ZN(n16279));
    NOR2X1 U3408 (.A1(N6815), .A2(N6816), .ZN(n16280));
    NOR2X1 U3409 (.A1(N6817), .A2(N6818), .ZN(n16281));
    NANDX1 U3410 (.A1(N6819), .A2(N6820), .ZN(N16282));
    NANDX1 U3411 (.A1(N6821), .A2(N6822), .ZN(N16283));
    NOR2X1 U3412 (.A1(N6823), .A2(N6824), .ZN(n16284));
    NOR2X1 U3413 (.A1(N6825), .A2(N6826), .ZN(n16285));
    NANDX1 U3414 (.A1(N6827), .A2(N6828), .ZN(n16286));
    NOR2X1 U3415 (.A1(N6829), .A2(N6830), .ZN(n16287));
    NOR2X1 U3416 (.A1(N6831), .A2(N6832), .ZN(n16288));
    NANDX1 U3417 (.A1(N6833), .A2(N6834), .ZN(N16289));
    NOR2X1 U3418 (.A1(N6835), .A2(N6836), .ZN(N16290));
    NOR2X1 U3419 (.A1(N6837), .A2(N6838), .ZN(n16291));
    NANDX1 U3420 (.A1(N6839), .A2(N6840), .ZN(n16292));
    NANDX1 U3421 (.A1(N6841), .A2(N6842), .ZN(n16293));
    NOR2X1 U3422 (.A1(N6843), .A2(N6844), .ZN(n16294));
    NOR2X1 U3423 (.A1(N6845), .A2(N6846), .ZN(n16295));
    NANDX1 U3424 (.A1(N6847), .A2(N6848), .ZN(n16296));
    NOR2X1 U3425 (.A1(N6849), .A2(N6850), .ZN(n16297));
    NOR2X1 U3426 (.A1(N6851), .A2(N6852), .ZN(n16298));
    NOR2X1 U3427 (.A1(N6853), .A2(N6854), .ZN(n16299));
    NOR2X1 U3428 (.A1(N6855), .A2(N6856), .ZN(n16300));
    NOR2X1 U3429 (.A1(N6857), .A2(N6858), .ZN(N16301));
    NOR2X1 U3430 (.A1(N6859), .A2(N6860), .ZN(n16302));
    NANDX1 U3431 (.A1(N6861), .A2(N6862), .ZN(N16303));
    NOR2X1 U3432 (.A1(N6863), .A2(N6864), .ZN(n16304));
    NANDX1 U3433 (.A1(N6865), .A2(N6866), .ZN(n16305));
    NOR2X1 U3434 (.A1(N6867), .A2(N6868), .ZN(n16306));
    NANDX1 U3435 (.A1(N6869), .A2(N6870), .ZN(n16307));
    NOR2X1 U3436 (.A1(N6871), .A2(N6872), .ZN(n16308));
    NOR2X1 U3437 (.A1(N6873), .A2(N6874), .ZN(n16309));
    NOR2X1 U3438 (.A1(N6875), .A2(N6876), .ZN(n16310));
    NOR2X1 U3439 (.A1(N6877), .A2(N6878), .ZN(n16311));
    NANDX1 U3440 (.A1(N6879), .A2(N6880), .ZN(n16312));
    NANDX1 U3441 (.A1(N6881), .A2(N6882), .ZN(n16313));
    NOR2X1 U3442 (.A1(N6883), .A2(N6884), .ZN(n16314));
    NANDX1 U3443 (.A1(N6885), .A2(N6886), .ZN(n16315));
    NOR2X1 U3444 (.A1(N6887), .A2(N6888), .ZN(n16316));
    NANDX1 U3445 (.A1(N6889), .A2(N6890), .ZN(n16317));
    NANDX1 U3446 (.A1(N6891), .A2(N6892), .ZN(n16318));
    NOR2X1 U3447 (.A1(N6893), .A2(N6894), .ZN(n16319));
    NOR2X1 U3448 (.A1(N6895), .A2(N6896), .ZN(n16320));
    NANDX1 U3449 (.A1(N6897), .A2(N6898), .ZN(n16321));
    NOR2X1 U3450 (.A1(N6899), .A2(N6900), .ZN(n16322));
    NOR2X1 U3451 (.A1(N6901), .A2(N6902), .ZN(N16323));
    NOR2X1 U3452 (.A1(N6903), .A2(N6904), .ZN(n16324));
    NANDX1 U3453 (.A1(N6905), .A2(N6906), .ZN(n16325));
    NOR2X1 U3454 (.A1(N6907), .A2(N6908), .ZN(N16326));
    NANDX1 U3455 (.A1(N6909), .A2(N6910), .ZN(n16327));
    NANDX1 U3456 (.A1(N6911), .A2(N6912), .ZN(N16328));
    NOR2X1 U3457 (.A1(N6913), .A2(N6914), .ZN(n16329));
    NOR2X1 U3458 (.A1(N6915), .A2(N6916), .ZN(N16330));
    NANDX1 U3459 (.A1(N6917), .A2(N6918), .ZN(n16331));
    NOR2X1 U3460 (.A1(N6919), .A2(N6920), .ZN(N16332));
    NOR2X1 U3461 (.A1(N6921), .A2(N6922), .ZN(n16333));
    NOR2X1 U3462 (.A1(N6923), .A2(N6924), .ZN(N16334));
    NOR2X1 U3463 (.A1(N6925), .A2(N6926), .ZN(n16335));
    NANDX1 U3464 (.A1(N6927), .A2(N6928), .ZN(n16336));
    NOR2X1 U3465 (.A1(N6929), .A2(N6930), .ZN(n16337));
    NOR2X1 U3466 (.A1(N6931), .A2(N6932), .ZN(n16338));
    NANDX1 U3467 (.A1(N6933), .A2(N6934), .ZN(n16339));
    NANDX1 U3468 (.A1(N6935), .A2(N6936), .ZN(n16340));
    NOR2X1 U3469 (.A1(N6937), .A2(N6938), .ZN(N16341));
    NOR2X1 U3470 (.A1(N6939), .A2(N6940), .ZN(n16342));
    NOR2X1 U3471 (.A1(N6941), .A2(N6942), .ZN(n16343));
    NOR2X1 U3472 (.A1(N6943), .A2(N6944), .ZN(n16344));
    NOR2X1 U3473 (.A1(N6945), .A2(N6946), .ZN(n16345));
    NANDX1 U3474 (.A1(N6947), .A2(N6948), .ZN(n16346));
    NOR2X1 U3475 (.A1(N6949), .A2(N6950), .ZN(n16347));
    NANDX1 U3476 (.A1(N6951), .A2(N6952), .ZN(n16348));
    NANDX1 U3477 (.A1(N6953), .A2(N6954), .ZN(n16349));
    NOR2X1 U3478 (.A1(N6955), .A2(N6956), .ZN(n16350));
    NANDX1 U3479 (.A1(N6957), .A2(N6958), .ZN(n16351));
    NOR2X1 U3480 (.A1(N6959), .A2(N6960), .ZN(n16352));
    NOR2X1 U3481 (.A1(N6961), .A2(N6962), .ZN(N16353));
    NANDX1 U3482 (.A1(N6963), .A2(N6964), .ZN(n16354));
    NANDX1 U3483 (.A1(N6965), .A2(N6966), .ZN(n16355));
    NANDX1 U3484 (.A1(N6967), .A2(N6968), .ZN(n16356));
    NANDX1 U3485 (.A1(N6969), .A2(N6970), .ZN(n16357));
    NOR2X1 U3486 (.A1(N6971), .A2(N6972), .ZN(n16358));
    NOR2X1 U3487 (.A1(N6973), .A2(N6974), .ZN(n16359));
    NOR2X1 U3488 (.A1(N6975), .A2(N6976), .ZN(n16360));
    NOR2X1 U3489 (.A1(N6977), .A2(N6978), .ZN(n16361));
    NOR2X1 U3490 (.A1(N6979), .A2(N6980), .ZN(n16362));
    NOR2X1 U3491 (.A1(N6981), .A2(N6982), .ZN(n16363));
    NOR2X1 U3492 (.A1(N6983), .A2(N6984), .ZN(N16364));
    NOR2X1 U3493 (.A1(N6985), .A2(N6986), .ZN(n16365));
    NANDX1 U3494 (.A1(N6987), .A2(N6988), .ZN(n16366));
    NANDX1 U3495 (.A1(N6989), .A2(N6990), .ZN(N16367));
    NANDX1 U3496 (.A1(N6991), .A2(N6992), .ZN(n16368));
    NANDX1 U3497 (.A1(N6993), .A2(N6994), .ZN(n16369));
    NANDX1 U3498 (.A1(N6995), .A2(N6996), .ZN(n16370));
    NOR2X1 U3499 (.A1(N6997), .A2(N6998), .ZN(n16371));
    NANDX1 U3500 (.A1(N6999), .A2(N7000), .ZN(n16372));
    NANDX1 U3501 (.A1(N7001), .A2(N7002), .ZN(n16373));
    NOR2X1 U3502 (.A1(N7003), .A2(N7004), .ZN(n16374));
    NANDX1 U3503 (.A1(N7005), .A2(N7006), .ZN(n16375));
    NANDX1 U3504 (.A1(N7007), .A2(N7008), .ZN(n16376));
    NANDX1 U3505 (.A1(N7009), .A2(N7010), .ZN(n16377));
    NANDX1 U3506 (.A1(N7011), .A2(N7012), .ZN(n16378));
    NOR2X1 U3507 (.A1(N7013), .A2(N7014), .ZN(N16379));
    NOR2X1 U3508 (.A1(N7015), .A2(N7016), .ZN(n16380));
    NANDX1 U3509 (.A1(N7017), .A2(N7018), .ZN(n16381));
    NANDX1 U3510 (.A1(N7019), .A2(N7020), .ZN(n16382));
    NANDX1 U3511 (.A1(N7021), .A2(N7022), .ZN(n16383));
    NOR2X1 U3512 (.A1(N7023), .A2(N7024), .ZN(n16384));
    NANDX1 U3513 (.A1(N7025), .A2(N7026), .ZN(N16385));
    NOR2X1 U3514 (.A1(N7027), .A2(N7028), .ZN(n16386));
    NANDX1 U3515 (.A1(N7029), .A2(N7030), .ZN(n16387));
    NOR2X1 U3516 (.A1(N7031), .A2(N7032), .ZN(n16388));
    NOR2X1 U3517 (.A1(N7033), .A2(N7034), .ZN(n16389));
    NOR2X1 U3518 (.A1(N7035), .A2(N7036), .ZN(n16390));
    NOR2X1 U3519 (.A1(N7037), .A2(N7038), .ZN(n16391));
    NANDX1 U3520 (.A1(N7039), .A2(N7040), .ZN(n16392));
    NOR2X1 U3521 (.A1(N7041), .A2(N7042), .ZN(n16393));
    NANDX1 U3522 (.A1(N7043), .A2(N7044), .ZN(N16394));
    NANDX1 U3523 (.A1(N7045), .A2(N7046), .ZN(n16395));
    NOR2X1 U3524 (.A1(N7047), .A2(N7048), .ZN(n16396));
    NOR2X1 U3525 (.A1(N7049), .A2(N7050), .ZN(n16397));
    NANDX1 U3526 (.A1(N7051), .A2(N7052), .ZN(N16398));
    NANDX1 U3527 (.A1(N7053), .A2(N7054), .ZN(n16399));
    NANDX1 U3528 (.A1(N7055), .A2(N7056), .ZN(N16400));
    NOR2X1 U3529 (.A1(N7057), .A2(N7058), .ZN(n16401));
    NANDX1 U3530 (.A1(N7059), .A2(N7060), .ZN(N16402));
    NOR2X1 U3531 (.A1(N7061), .A2(N7062), .ZN(N16403));
    NANDX1 U3532 (.A1(N7063), .A2(N7064), .ZN(n16404));
    NANDX1 U3533 (.A1(N7065), .A2(N7066), .ZN(n16405));
    NOR2X1 U3534 (.A1(N7067), .A2(N7068), .ZN(n16406));
    NOR2X1 U3535 (.A1(N7069), .A2(N7070), .ZN(n16407));
    NANDX1 U3536 (.A1(N7071), .A2(N7072), .ZN(n16408));
    NANDX1 U3537 (.A1(N7073), .A2(N7074), .ZN(N16409));
    NOR2X1 U3538 (.A1(N7075), .A2(N7076), .ZN(n16410));
    NANDX1 U3539 (.A1(N7077), .A2(N7078), .ZN(n16411));
    NANDX1 U3540 (.A1(N7079), .A2(N7080), .ZN(n16412));
    NANDX1 U3541 (.A1(N7081), .A2(N7082), .ZN(n16413));
    NOR2X1 U3542 (.A1(N7083), .A2(N7084), .ZN(n16414));
    NANDX1 U3543 (.A1(N7085), .A2(N7086), .ZN(n16415));
    NOR2X1 U3544 (.A1(N7087), .A2(N7088), .ZN(N16416));
    NOR2X1 U3545 (.A1(N7089), .A2(N7090), .ZN(N16417));
    NOR2X1 U3546 (.A1(N7091), .A2(N7092), .ZN(n16418));
    NANDX1 U3547 (.A1(N7093), .A2(N7094), .ZN(n16419));
    NANDX1 U3548 (.A1(N7095), .A2(N7096), .ZN(n16420));
    NOR2X1 U3549 (.A1(N7097), .A2(N7098), .ZN(N16421));
    NANDX1 U3550 (.A1(N7099), .A2(N7100), .ZN(n16422));
    NOR2X1 U3551 (.A1(N7101), .A2(N7102), .ZN(n16423));
    NOR2X1 U3552 (.A1(N7103), .A2(N7104), .ZN(n16424));
    NOR2X1 U3553 (.A1(N7105), .A2(N7106), .ZN(n16425));
    NANDX1 U3554 (.A1(N7107), .A2(N7108), .ZN(n16426));
    NANDX1 U3555 (.A1(N7109), .A2(N7110), .ZN(n16427));
    NOR2X1 U3556 (.A1(N7111), .A2(N7112), .ZN(N16428));
    NOR2X1 U3557 (.A1(N7113), .A2(N7114), .ZN(n16429));
    NOR2X1 U3558 (.A1(N7115), .A2(N7116), .ZN(n16430));
    NANDX1 U3559 (.A1(N7117), .A2(N7118), .ZN(n16431));
    NOR2X1 U3560 (.A1(N7119), .A2(N7120), .ZN(n16432));
    NOR2X1 U3561 (.A1(N7121), .A2(N7122), .ZN(n16433));
    NOR2X1 U3562 (.A1(N7123), .A2(N7124), .ZN(n16434));
    NANDX1 U3563 (.A1(N7125), .A2(N7126), .ZN(n16435));
    NANDX1 U3564 (.A1(N7127), .A2(N7128), .ZN(n16436));
    NOR2X1 U3565 (.A1(N7129), .A2(N7130), .ZN(n16437));
    NANDX1 U3566 (.A1(N7131), .A2(N7132), .ZN(n16438));
    NOR2X1 U3567 (.A1(N7133), .A2(N7134), .ZN(n16439));
    NANDX1 U3568 (.A1(N7135), .A2(N7136), .ZN(n16440));
    NANDX1 U3569 (.A1(N7137), .A2(N7138), .ZN(n16441));
    NOR2X1 U3570 (.A1(N7139), .A2(N7140), .ZN(N16442));
    NOR2X1 U3571 (.A1(N7141), .A2(N7142), .ZN(n16443));
    NANDX1 U3572 (.A1(N7143), .A2(N7144), .ZN(n16444));
    NOR2X1 U3573 (.A1(N7145), .A2(N7146), .ZN(n16445));
    NANDX1 U3574 (.A1(N7147), .A2(N7148), .ZN(n16446));
    NANDX1 U3575 (.A1(N7149), .A2(N7150), .ZN(n16447));
    NANDX1 U3576 (.A1(N7151), .A2(N7152), .ZN(n16448));
    NOR2X1 U3577 (.A1(N7153), .A2(N7154), .ZN(n16449));
    NOR2X1 U3578 (.A1(N7155), .A2(N7156), .ZN(N16450));
    NOR2X1 U3579 (.A1(N7157), .A2(N7158), .ZN(n16451));
    NOR2X1 U3580 (.A1(N7159), .A2(N7160), .ZN(n16452));
    NOR2X1 U3581 (.A1(N7161), .A2(N7162), .ZN(N16453));
    NOR2X1 U3582 (.A1(N7163), .A2(N7164), .ZN(n16454));
    NANDX1 U3583 (.A1(N7165), .A2(N7166), .ZN(n16455));
    NOR2X1 U3584 (.A1(N7167), .A2(N7168), .ZN(n16456));
    NANDX1 U3585 (.A1(N7169), .A2(N7170), .ZN(N16457));
    NOR2X1 U3586 (.A1(N7171), .A2(N7172), .ZN(N16458));
    NANDX1 U3587 (.A1(N7173), .A2(N7174), .ZN(n16459));
    NOR2X1 U3588 (.A1(N7175), .A2(N7176), .ZN(n16460));
    NOR2X1 U3589 (.A1(N7177), .A2(N7178), .ZN(n16461));
    NOR2X1 U3590 (.A1(N7179), .A2(N7180), .ZN(N16462));
    NOR2X1 U3591 (.A1(N7181), .A2(N7182), .ZN(n16463));
    NOR2X1 U3592 (.A1(N7183), .A2(N7184), .ZN(n16464));
    NOR2X1 U3593 (.A1(N7185), .A2(N7186), .ZN(n16465));
    NOR2X1 U3594 (.A1(N7187), .A2(N7188), .ZN(N16466));
    NOR2X1 U3595 (.A1(N7189), .A2(N7190), .ZN(n16467));
    NOR2X1 U3596 (.A1(N7191), .A2(N7192), .ZN(n16468));
    NANDX1 U3597 (.A1(N7193), .A2(N7194), .ZN(n16469));
    NOR2X1 U3598 (.A1(N7195), .A2(N7196), .ZN(n16470));
    NOR2X1 U3599 (.A1(N7197), .A2(N7198), .ZN(n16471));
    NANDX1 U3600 (.A1(N7199), .A2(N7200), .ZN(n16472));
    NOR2X1 U3601 (.A1(N7201), .A2(N7202), .ZN(n16473));
    NOR2X1 U3602 (.A1(N7203), .A2(N7204), .ZN(N16474));
    NOR2X1 U3603 (.A1(N7205), .A2(N7206), .ZN(n16475));
    NANDX1 U3604 (.A1(N7207), .A2(N7208), .ZN(n16476));
    NOR2X1 U3605 (.A1(N7209), .A2(N7210), .ZN(n16477));
    NANDX1 U3606 (.A1(N7211), .A2(N7212), .ZN(n16478));
    NOR2X1 U3607 (.A1(N7213), .A2(N7214), .ZN(n16479));
    NOR2X1 U3608 (.A1(N7215), .A2(N7216), .ZN(N16480));
    NOR2X1 U3609 (.A1(N7217), .A2(N7218), .ZN(n16481));
    NOR2X1 U3610 (.A1(N7219), .A2(N7220), .ZN(n16482));
    NOR2X1 U3611 (.A1(N7221), .A2(N7222), .ZN(n16483));
    NOR2X1 U3612 (.A1(N7223), .A2(N7224), .ZN(n16484));
    NOR2X1 U3613 (.A1(N7225), .A2(N7226), .ZN(n16485));
    NANDX1 U3614 (.A1(N7227), .A2(N7228), .ZN(n16486));
    NOR2X1 U3615 (.A1(N7229), .A2(N7230), .ZN(N16487));
    NANDX1 U3616 (.A1(N7231), .A2(N7232), .ZN(n16488));
    NANDX1 U3617 (.A1(N7233), .A2(N7234), .ZN(n16489));
    NANDX1 U3618 (.A1(N7235), .A2(N7236), .ZN(n16490));
    NANDX1 U3619 (.A1(N7237), .A2(N7238), .ZN(n16491));
    NOR2X1 U3620 (.A1(N7239), .A2(N7240), .ZN(n16492));
    NOR2X1 U3621 (.A1(N7241), .A2(N7242), .ZN(n16493));
    NOR2X1 U3622 (.A1(N7243), .A2(N7244), .ZN(N16494));
    NOR2X1 U3623 (.A1(N7245), .A2(N7246), .ZN(n16495));
    NOR2X1 U3624 (.A1(N7247), .A2(N7248), .ZN(n16496));
    NOR2X1 U3625 (.A1(N7249), .A2(N7250), .ZN(n16497));
    NOR2X1 U3626 (.A1(N7251), .A2(N7252), .ZN(n16498));
    NANDX1 U3627 (.A1(N7253), .A2(N7254), .ZN(N16499));
    NANDX1 U3628 (.A1(N7255), .A2(N7256), .ZN(n16500));
    NANDX1 U3629 (.A1(N7257), .A2(N7258), .ZN(n16501));
    NANDX1 U3630 (.A1(N7259), .A2(N7260), .ZN(n16502));
    NOR2X1 U3631 (.A1(N7261), .A2(N7262), .ZN(n16503));
    NANDX1 U3632 (.A1(N7263), .A2(N7264), .ZN(n16504));
    NANDX1 U3633 (.A1(N7265), .A2(N7266), .ZN(n16505));
    NOR2X1 U3634 (.A1(N7267), .A2(N7268), .ZN(n16506));
    NOR2X1 U3635 (.A1(N7269), .A2(N7270), .ZN(n16507));
    NANDX1 U3636 (.A1(N7271), .A2(N7272), .ZN(n16508));
    NOR2X1 U3637 (.A1(N7273), .A2(N7274), .ZN(n16509));
    NOR2X1 U3638 (.A1(N7275), .A2(N7276), .ZN(n16510));
    NANDX1 U3639 (.A1(N7277), .A2(N7278), .ZN(n16511));
    NOR2X1 U3640 (.A1(N7279), .A2(N7280), .ZN(n16512));
    NOR2X1 U3641 (.A1(N7281), .A2(N7282), .ZN(n16513));
    NOR2X1 U3642 (.A1(N7283), .A2(N7284), .ZN(n16514));
    NOR2X1 U3643 (.A1(N7285), .A2(N7286), .ZN(n16515));
    NOR2X1 U3644 (.A1(N7287), .A2(N7288), .ZN(N16516));
    NANDX1 U3645 (.A1(N7289), .A2(N7290), .ZN(n16517));
    NOR2X1 U3646 (.A1(N7291), .A2(N7292), .ZN(n16518));
    NOR2X1 U3647 (.A1(N7293), .A2(N7294), .ZN(N16519));
    NANDX1 U3648 (.A1(N7295), .A2(N7296), .ZN(n16520));
    NOR2X1 U3649 (.A1(N7297), .A2(N7298), .ZN(n16521));
    NANDX1 U3650 (.A1(N7299), .A2(N7300), .ZN(n16522));
    NANDX1 U3651 (.A1(N7301), .A2(N7302), .ZN(n16523));
    NOR2X1 U3652 (.A1(N7303), .A2(N7304), .ZN(n16524));
    NANDX1 U3653 (.A1(N7305), .A2(N7306), .ZN(n16525));
    NANDX1 U3654 (.A1(N7307), .A2(N7308), .ZN(n16526));
    NOR2X1 U3655 (.A1(N7309), .A2(N7310), .ZN(N16527));
    NANDX1 U3656 (.A1(N7311), .A2(N7312), .ZN(n16528));
    NOR2X1 U3657 (.A1(N7313), .A2(N7314), .ZN(N16529));
    NANDX1 U3658 (.A1(N7315), .A2(N7316), .ZN(n16530));
    NANDX1 U3659 (.A1(N7317), .A2(N7318), .ZN(n16531));
    NANDX1 U3660 (.A1(N7319), .A2(N7320), .ZN(n16532));
    NOR2X1 U3661 (.A1(N7321), .A2(N7322), .ZN(N16533));
    NANDX1 U3662 (.A1(N7323), .A2(N7324), .ZN(n16534));
    NOR2X1 U3663 (.A1(N7325), .A2(N7326), .ZN(n16535));
    NOR2X1 U3664 (.A1(N7327), .A2(N7328), .ZN(n16536));
    NOR2X1 U3665 (.A1(N7329), .A2(N7330), .ZN(N16537));
    NANDX1 U3666 (.A1(N7331), .A2(N7332), .ZN(n16538));
    NANDX1 U3667 (.A1(N7333), .A2(N7334), .ZN(n16539));
    NOR2X1 U3668 (.A1(N7335), .A2(N7336), .ZN(n16540));
    NANDX1 U3669 (.A1(N7337), .A2(N7338), .ZN(n16541));
    NANDX1 U3670 (.A1(N7339), .A2(N7340), .ZN(n16542));
    NOR2X1 U3671 (.A1(N7341), .A2(N7342), .ZN(n16543));
    NOR2X1 U3672 (.A1(N7343), .A2(N7344), .ZN(n16544));
    NANDX1 U3673 (.A1(N7345), .A2(N7346), .ZN(n16545));
    NOR2X1 U3674 (.A1(N7347), .A2(N7348), .ZN(n16546));
    NOR2X1 U3675 (.A1(N7349), .A2(N7350), .ZN(n16547));
    NOR2X1 U3676 (.A1(N7351), .A2(N7352), .ZN(n16548));
    NOR2X1 U3677 (.A1(N7353), .A2(N7354), .ZN(n16549));
    NOR2X1 U3678 (.A1(N7355), .A2(N7356), .ZN(n16550));
    NANDX1 U3679 (.A1(N7357), .A2(N7358), .ZN(N16551));
    NOR2X1 U3680 (.A1(N7359), .A2(N7360), .ZN(n16552));
    NOR2X1 U3681 (.A1(N7361), .A2(N7362), .ZN(n16553));
    NOR2X1 U3682 (.A1(N7363), .A2(N7364), .ZN(n16554));
    NOR2X1 U3683 (.A1(N7365), .A2(N7366), .ZN(n16555));
    NANDX1 U3684 (.A1(N7367), .A2(N7368), .ZN(N16556));
    NOR2X1 U3685 (.A1(N7369), .A2(N7370), .ZN(n16557));
    NANDX1 U3686 (.A1(N7371), .A2(N7372), .ZN(n16558));
    NANDX1 U3687 (.A1(N7373), .A2(N7374), .ZN(n16559));
    NOR2X1 U3688 (.A1(N7375), .A2(N7376), .ZN(N16560));
    NOR2X1 U3689 (.A1(N7377), .A2(N7378), .ZN(n16561));
    NOR2X1 U3690 (.A1(N7379), .A2(N7380), .ZN(n16562));
    NANDX1 U3691 (.A1(N7381), .A2(N7382), .ZN(n16563));
    NANDX1 U3692 (.A1(N7383), .A2(N7384), .ZN(n16564));
    NANDX1 U3693 (.A1(N7385), .A2(N7386), .ZN(N16565));
    NANDX1 U3694 (.A1(N7387), .A2(N7388), .ZN(n16566));
    NANDX1 U3695 (.A1(N7389), .A2(N7390), .ZN(n16567));
    NANDX1 U3696 (.A1(N7391), .A2(N7392), .ZN(n16568));
    NOR2X1 U3697 (.A1(N7393), .A2(N7394), .ZN(n16569));
    NOR2X1 U3698 (.A1(N7395), .A2(N7396), .ZN(n16570));
    NANDX1 U3699 (.A1(N7397), .A2(N7398), .ZN(N16571));
    NOR2X1 U3700 (.A1(N7399), .A2(N7400), .ZN(n16572));
    NANDX1 U3701 (.A1(N7401), .A2(N7402), .ZN(n16573));
    NANDX1 U3702 (.A1(N7403), .A2(N7404), .ZN(n16574));
    NOR2X1 U3703 (.A1(N7405), .A2(N7406), .ZN(n16575));
    NOR2X1 U3704 (.A1(N7407), .A2(N7408), .ZN(N16576));
    NANDX1 U3705 (.A1(N7409), .A2(N7410), .ZN(n16577));
    NOR2X1 U3706 (.A1(N7411), .A2(N7412), .ZN(N16578));
    NANDX1 U3707 (.A1(N7413), .A2(N7414), .ZN(n16579));
    NOR2X1 U3708 (.A1(N7415), .A2(N7416), .ZN(n16580));
    NANDX1 U3709 (.A1(N7417), .A2(N7418), .ZN(n16581));
    NOR2X1 U3710 (.A1(N7419), .A2(N7420), .ZN(N16582));
    NOR2X1 U3711 (.A1(N7421), .A2(N7422), .ZN(n16583));
    NANDX1 U3712 (.A1(N7423), .A2(N7424), .ZN(n16584));
    NANDX1 U3713 (.A1(N7425), .A2(N7426), .ZN(n16585));
    NANDX1 U3714 (.A1(N7427), .A2(N7428), .ZN(N16586));
    NOR2X1 U3715 (.A1(N7429), .A2(N7430), .ZN(n16587));
    NANDX1 U3716 (.A1(N7431), .A2(N7432), .ZN(n16588));
    NOR2X1 U3717 (.A1(N7433), .A2(N7434), .ZN(n16589));
    NANDX1 U3718 (.A1(N7435), .A2(N7436), .ZN(n16590));
    NANDX1 U3719 (.A1(N7437), .A2(N7438), .ZN(N16591));
    NOR2X1 U3720 (.A1(N7439), .A2(N7440), .ZN(N16592));
    NANDX1 U3721 (.A1(N7441), .A2(N7442), .ZN(n16593));
    NOR2X1 U3722 (.A1(N7443), .A2(N7444), .ZN(n16594));
    NANDX1 U3723 (.A1(N7445), .A2(N7446), .ZN(n16595));
    NANDX1 U3724 (.A1(N7447), .A2(N7448), .ZN(n16596));
    NANDX1 U3725 (.A1(N7449), .A2(N7450), .ZN(n16597));
    NOR2X1 U3726 (.A1(N7451), .A2(N7452), .ZN(N16598));
    NOR2X1 U3727 (.A1(N7453), .A2(N7454), .ZN(n16599));
    NOR2X1 U3728 (.A1(N7455), .A2(N7456), .ZN(n16600));
    NANDX1 U3729 (.A1(N7457), .A2(N7458), .ZN(N16601));
    NOR2X1 U3730 (.A1(N7459), .A2(N7460), .ZN(N16602));
    NOR2X1 U3731 (.A1(N7461), .A2(N7462), .ZN(n16603));
    NOR2X1 U3732 (.A1(N7463), .A2(N7464), .ZN(n16604));
    NANDX1 U3733 (.A1(N7465), .A2(N7466), .ZN(n16605));
    NOR2X1 U3734 (.A1(N7467), .A2(N7468), .ZN(n16606));
    NANDX1 U3735 (.A1(N7469), .A2(N7470), .ZN(n16607));
    NANDX1 U3736 (.A1(N7471), .A2(N7472), .ZN(n16608));
    NOR2X1 U3737 (.A1(N7473), .A2(N7474), .ZN(n16609));
    NOR2X1 U3738 (.A1(N7475), .A2(N7476), .ZN(n16610));
    NANDX1 U3739 (.A1(N7477), .A2(N7478), .ZN(n16611));
    NANDX1 U3740 (.A1(N7479), .A2(N7480), .ZN(n16612));
    NOR2X1 U3741 (.A1(N7481), .A2(N7482), .ZN(n16613));
    NANDX1 U3742 (.A1(N7483), .A2(N7484), .ZN(n16614));
    NOR2X1 U3743 (.A1(N7485), .A2(N7486), .ZN(n16615));
    NANDX1 U3744 (.A1(N7487), .A2(N7488), .ZN(N16616));
    NOR2X1 U3745 (.A1(N7489), .A2(N7490), .ZN(n16617));
    NANDX1 U3746 (.A1(N7491), .A2(N7492), .ZN(n16618));
    NOR2X1 U3747 (.A1(N7493), .A2(N7494), .ZN(n16619));
    NOR2X1 U3748 (.A1(N7495), .A2(N7496), .ZN(n16620));
    NOR2X1 U3749 (.A1(N7497), .A2(N7498), .ZN(n16621));
    NANDX1 U3750 (.A1(N7499), .A2(N7500), .ZN(n16622));
    NANDX1 U3751 (.A1(N7501), .A2(N7502), .ZN(n16623));
    NOR2X1 U3752 (.A1(N7503), .A2(N7504), .ZN(n16624));
    NANDX1 U3753 (.A1(N7505), .A2(N7506), .ZN(n16625));
    NOR2X1 U3754 (.A1(N7507), .A2(N7508), .ZN(n16626));
    NANDX1 U3755 (.A1(N7509), .A2(N7510), .ZN(n16627));
    NANDX1 U3756 (.A1(N7511), .A2(N7512), .ZN(n16628));
    NANDX1 U3757 (.A1(N7513), .A2(N7514), .ZN(N16629));
    NANDX1 U3758 (.A1(N7515), .A2(N7516), .ZN(n16630));
    NANDX1 U3759 (.A1(N7517), .A2(N7518), .ZN(N16631));
    NOR2X1 U3760 (.A1(N7519), .A2(N7520), .ZN(N16632));
    NANDX1 U3761 (.A1(N7521), .A2(N7522), .ZN(n16633));
    NANDX1 U3762 (.A1(N7523), .A2(N7524), .ZN(N16634));
    NOR2X1 U3763 (.A1(N7525), .A2(N7526), .ZN(n16635));
    NANDX1 U3764 (.A1(N7527), .A2(N7528), .ZN(n16636));
    NANDX1 U3765 (.A1(N7529), .A2(N7530), .ZN(n16637));
    NANDX1 U3766 (.A1(N7531), .A2(N7532), .ZN(n16638));
    NOR2X1 U3767 (.A1(N7533), .A2(N7534), .ZN(n16639));
    NANDX1 U3768 (.A1(N7535), .A2(N7536), .ZN(n16640));
    NANDX1 U3769 (.A1(N7537), .A2(N7538), .ZN(n16641));
    NANDX1 U3770 (.A1(N7539), .A2(N7540), .ZN(N16642));
    NANDX1 U3771 (.A1(N7541), .A2(N7542), .ZN(n16643));
    NOR2X1 U3772 (.A1(N7543), .A2(N7544), .ZN(n16644));
    NOR2X1 U3773 (.A1(N7545), .A2(N7546), .ZN(N16645));
    NANDX1 U3774 (.A1(N7547), .A2(N7548), .ZN(n16646));
    NANDX1 U3775 (.A1(N7549), .A2(N7550), .ZN(n16647));
    NANDX1 U3776 (.A1(N7551), .A2(N7552), .ZN(n16648));
    NOR2X1 U3777 (.A1(N7553), .A2(N7554), .ZN(N16649));
    NOR2X1 U3778 (.A1(N7555), .A2(N7556), .ZN(n16650));
    NANDX1 U3779 (.A1(N7557), .A2(N7558), .ZN(n16651));
    NANDX1 U3780 (.A1(N7559), .A2(N7560), .ZN(n16652));
    NANDX1 U3781 (.A1(N7561), .A2(N7562), .ZN(n16653));
    NOR2X1 U3782 (.A1(N7563), .A2(N7564), .ZN(n16654));
    NANDX1 U3783 (.A1(N7565), .A2(N7566), .ZN(n16655));
    NANDX1 U3784 (.A1(N7567), .A2(N7568), .ZN(n16656));
    NANDX1 U3785 (.A1(N7569), .A2(N7570), .ZN(n16657));
    NOR2X1 U3786 (.A1(N7571), .A2(N7572), .ZN(n16658));
    NOR2X1 U3787 (.A1(N7573), .A2(N7574), .ZN(n16659));
    NOR2X1 U3788 (.A1(N7575), .A2(N7576), .ZN(n16660));
    NANDX1 U3789 (.A1(N7577), .A2(N7578), .ZN(n16661));
    NANDX1 U3790 (.A1(N7579), .A2(N7580), .ZN(n16662));
    NOR2X1 U3791 (.A1(N7581), .A2(N7582), .ZN(n16663));
    NANDX1 U3792 (.A1(N7583), .A2(N7584), .ZN(n16664));
    NOR2X1 U3793 (.A1(N7585), .A2(N7586), .ZN(n16665));
    NOR2X1 U3794 (.A1(N7587), .A2(N7588), .ZN(N16666));
    NOR2X1 U3795 (.A1(N7589), .A2(N7590), .ZN(N16667));
    NANDX1 U3796 (.A1(N7591), .A2(N7592), .ZN(n16668));
    NOR2X1 U3797 (.A1(N7593), .A2(N7594), .ZN(n16669));
    NOR2X1 U3798 (.A1(N7595), .A2(N7596), .ZN(n16670));
    NOR2X1 U3799 (.A1(N7597), .A2(N7598), .ZN(n16671));
    NANDX1 U3800 (.A1(N7599), .A2(N7600), .ZN(n16672));
    NANDX1 U3801 (.A1(N7601), .A2(N7602), .ZN(n16673));
    NANDX1 U3802 (.A1(N7603), .A2(N7604), .ZN(N16674));
    NANDX1 U3803 (.A1(N7605), .A2(N7606), .ZN(n16675));
    NANDX1 U3804 (.A1(N7607), .A2(N7608), .ZN(n16676));
    NANDX1 U3805 (.A1(N7609), .A2(N7610), .ZN(N16677));
    NANDX1 U3806 (.A1(N7611), .A2(N7612), .ZN(n16678));
    NOR2X1 U3807 (.A1(N7613), .A2(N7614), .ZN(n16679));
    NANDX1 U3808 (.A1(N7615), .A2(N7616), .ZN(n16680));
    NANDX1 U3809 (.A1(N7617), .A2(N7618), .ZN(n16681));
    NOR2X1 U3810 (.A1(N7619), .A2(N7620), .ZN(N16682));
    NOR2X1 U3811 (.A1(N7621), .A2(N7622), .ZN(n16683));
    NOR2X1 U3812 (.A1(N7623), .A2(N7624), .ZN(N16684));
    NOR2X1 U3813 (.A1(N7625), .A2(N7626), .ZN(n16685));
    NANDX1 U3814 (.A1(N7627), .A2(N7628), .ZN(n16686));
    NANDX1 U3815 (.A1(N7629), .A2(N7630), .ZN(N16687));
    NANDX1 U3816 (.A1(N7631), .A2(N7632), .ZN(n16688));
    NANDX1 U3817 (.A1(N7633), .A2(N7634), .ZN(n16689));
    NANDX1 U3818 (.A1(N7635), .A2(N7636), .ZN(n16690));
    NANDX1 U3819 (.A1(N7637), .A2(N7638), .ZN(n16691));
    NANDX1 U3820 (.A1(N7639), .A2(N7640), .ZN(n16692));
    NOR2X1 U3821 (.A1(N7641), .A2(N7642), .ZN(n16693));
    NANDX1 U3822 (.A1(N7643), .A2(N7644), .ZN(n16694));
    NOR2X1 U3823 (.A1(N7645), .A2(N7646), .ZN(N16695));
    NOR2X1 U3824 (.A1(N7647), .A2(N7648), .ZN(n16696));
    NOR2X1 U3825 (.A1(N7649), .A2(N7650), .ZN(n16697));
    NOR2X1 U3826 (.A1(N7651), .A2(N7652), .ZN(n16698));
    NANDX1 U3827 (.A1(N7653), .A2(N7654), .ZN(n16699));
    NOR2X1 U3828 (.A1(N7655), .A2(N7656), .ZN(n16700));
    NOR2X1 U3829 (.A1(N7657), .A2(N7658), .ZN(n16701));
    NOR2X1 U3830 (.A1(N7659), .A2(N7660), .ZN(n16702));
    NANDX1 U3831 (.A1(N7661), .A2(N7662), .ZN(n16703));
    NANDX1 U3832 (.A1(N7663), .A2(N7664), .ZN(n16704));
    NANDX1 U3833 (.A1(N7665), .A2(N7666), .ZN(n16705));
    NANDX1 U3834 (.A1(N7667), .A2(N7668), .ZN(n16706));
    NOR2X1 U3835 (.A1(N7669), .A2(N7670), .ZN(n16707));
    NOR2X1 U3836 (.A1(N7671), .A2(N7672), .ZN(n16708));
    NOR2X1 U3837 (.A1(N7673), .A2(N7674), .ZN(N16709));
    NANDX1 U3838 (.A1(N7675), .A2(N7676), .ZN(n16710));
    NOR2X1 U3839 (.A1(N7677), .A2(N7678), .ZN(n16711));
    NANDX1 U3840 (.A1(N7679), .A2(N7680), .ZN(n16712));
    NANDX1 U3841 (.A1(N7681), .A2(N7682), .ZN(n16713));
    NOR2X1 U3842 (.A1(N7683), .A2(N7684), .ZN(n16714));
    NANDX1 U3843 (.A1(N7685), .A2(N7686), .ZN(n16715));
    NANDX1 U3844 (.A1(N7687), .A2(N7688), .ZN(n16716));
    NOR2X1 U3845 (.A1(N7689), .A2(N7690), .ZN(N16717));
    NANDX1 U3846 (.A1(N7691), .A2(N7692), .ZN(n16718));
    NANDX1 U3847 (.A1(N7693), .A2(N7694), .ZN(n16719));
    NANDX1 U3848 (.A1(N7695), .A2(N7696), .ZN(n16720));
    NOR2X1 U3849 (.A1(N7697), .A2(N7698), .ZN(n16721));
    NOR2X1 U3850 (.A1(N7699), .A2(N7700), .ZN(n16722));
    NOR2X1 U3851 (.A1(N7701), .A2(N7702), .ZN(n16723));
    NANDX1 U3852 (.A1(N7703), .A2(N7704), .ZN(n16724));
    NOR2X1 U3853 (.A1(N7705), .A2(N7706), .ZN(N16725));
    NOR2X1 U3854 (.A1(N7707), .A2(N7708), .ZN(n16726));
    NANDX1 U3855 (.A1(N7709), .A2(N7710), .ZN(n16727));
    NOR2X1 U3856 (.A1(N7711), .A2(N7712), .ZN(n16728));
    NOR2X1 U3857 (.A1(N7713), .A2(N7714), .ZN(n16729));
    NANDX1 U3858 (.A1(N7715), .A2(N7716), .ZN(N16730));
    NOR2X1 U3859 (.A1(N7717), .A2(N7718), .ZN(n16731));
    NOR2X1 U3860 (.A1(N7719), .A2(N7720), .ZN(n16732));
    NANDX1 U3861 (.A1(N7721), .A2(N7722), .ZN(n16733));
    NANDX1 U3862 (.A1(N7723), .A2(N7724), .ZN(n16734));
    NANDX1 U3863 (.A1(N7725), .A2(N7726), .ZN(n16735));
    NOR2X1 U3864 (.A1(N7727), .A2(N7728), .ZN(n16736));
    NOR2X1 U3865 (.A1(N7729), .A2(N7730), .ZN(n16737));
    NOR2X1 U3866 (.A1(N7731), .A2(N7732), .ZN(N16738));
    NANDX1 U3867 (.A1(N7733), .A2(N7734), .ZN(n16739));
    NOR2X1 U3868 (.A1(N7735), .A2(N7736), .ZN(n16740));
    NANDX1 U3869 (.A1(N7737), .A2(N7738), .ZN(n16741));
    NANDX1 U3870 (.A1(N7739), .A2(N7740), .ZN(N16742));
    NANDX1 U3871 (.A1(N7741), .A2(N7742), .ZN(n16743));
    NOR2X1 U3872 (.A1(N7743), .A2(N7744), .ZN(n16744));
    NANDX1 U3873 (.A1(N7745), .A2(N7746), .ZN(n16745));
    NANDX1 U3874 (.A1(N7747), .A2(N7748), .ZN(n16746));
    NANDX1 U3875 (.A1(N7749), .A2(N7750), .ZN(N16747));
    NANDX1 U3876 (.A1(N7751), .A2(N7752), .ZN(n16748));
    NOR2X1 U3877 (.A1(N7753), .A2(N7754), .ZN(n16749));
    NOR2X1 U3878 (.A1(N7755), .A2(N7756), .ZN(n16750));
    NANDX1 U3879 (.A1(N7757), .A2(N7758), .ZN(n16751));
    NOR2X1 U3880 (.A1(N7759), .A2(N7760), .ZN(n16752));
    NANDX1 U3881 (.A1(N7761), .A2(N7762), .ZN(n16753));
    NANDX1 U3882 (.A1(N7763), .A2(N7764), .ZN(n16754));
    NANDX1 U3883 (.A1(N7765), .A2(N7766), .ZN(n16755));
    NANDX1 U3884 (.A1(N7767), .A2(N7768), .ZN(n16756));
    NOR2X1 U3885 (.A1(N7769), .A2(N7770), .ZN(n16757));
    NANDX1 U3886 (.A1(N7771), .A2(N7772), .ZN(n16758));
    NANDX1 U3887 (.A1(N7773), .A2(N7774), .ZN(n16759));
    NOR2X1 U3888 (.A1(N7775), .A2(N7776), .ZN(N16760));
    NOR2X1 U3889 (.A1(N7777), .A2(N7778), .ZN(n16761));
    NANDX1 U3890 (.A1(N7779), .A2(N7780), .ZN(n16762));
    NANDX1 U3891 (.A1(N7781), .A2(N7782), .ZN(n16763));
    NANDX1 U3892 (.A1(N7783), .A2(N7784), .ZN(n16764));
    NOR2X1 U3893 (.A1(N7785), .A2(N7786), .ZN(N16765));
    NOR2X1 U3894 (.A1(N7787), .A2(N7788), .ZN(n16766));
    NANDX1 U3895 (.A1(N7789), .A2(N7790), .ZN(n16767));
    NANDX1 U3896 (.A1(N7791), .A2(N7792), .ZN(n16768));
    NOR2X1 U3897 (.A1(N7793), .A2(N7794), .ZN(n16769));
    NOR2X1 U3898 (.A1(N7795), .A2(N7796), .ZN(n16770));
    NANDX1 U3899 (.A1(N7797), .A2(N7798), .ZN(n16771));
    NANDX1 U3900 (.A1(N7799), .A2(N7800), .ZN(n16772));
    NANDX1 U3901 (.A1(N7801), .A2(N7802), .ZN(n16773));
    NANDX1 U3902 (.A1(N7803), .A2(N7804), .ZN(n16774));
    NANDX1 U3903 (.A1(N7805), .A2(N7806), .ZN(n16775));
    NANDX1 U3904 (.A1(N7807), .A2(N7808), .ZN(n16776));
    NOR2X1 U3905 (.A1(N7809), .A2(N7810), .ZN(n16777));
    NANDX1 U3906 (.A1(N7811), .A2(N7812), .ZN(n16778));
    NOR2X1 U3907 (.A1(N7813), .A2(N7814), .ZN(n16779));
    NOR2X1 U3908 (.A1(N7815), .A2(N7816), .ZN(n16780));
    NANDX1 U3909 (.A1(N7817), .A2(N7818), .ZN(n16781));
    NANDX1 U3910 (.A1(N7819), .A2(N7820), .ZN(N16782));
    NOR2X1 U3911 (.A1(N7821), .A2(N7822), .ZN(n16783));
    NOR2X1 U3912 (.A1(N7823), .A2(N7824), .ZN(n16784));
    NANDX1 U3913 (.A1(N7825), .A2(N7826), .ZN(n16785));
    NOR2X1 U3914 (.A1(N7827), .A2(N7828), .ZN(n16786));
    NANDX1 U3915 (.A1(N7829), .A2(N7830), .ZN(n16787));
    NANDX1 U3916 (.A1(N7831), .A2(N7832), .ZN(n16788));
    NANDX1 U3917 (.A1(N7833), .A2(N7834), .ZN(n16789));
    NOR2X1 U3918 (.A1(N7835), .A2(N7836), .ZN(n16790));
    NANDX1 U3919 (.A1(N7837), .A2(N7838), .ZN(n16791));
    NANDX1 U3920 (.A1(N7839), .A2(N7840), .ZN(n16792));
    NANDX1 U3921 (.A1(N7841), .A2(N7842), .ZN(n16793));
    NOR2X1 U3922 (.A1(N7843), .A2(N7844), .ZN(n16794));
    NOR2X1 U3923 (.A1(N7845), .A2(N7846), .ZN(n16795));
    NOR2X1 U3924 (.A1(N7847), .A2(N7848), .ZN(N16796));
    NANDX1 U3925 (.A1(N7849), .A2(N7850), .ZN(N16797));
    NANDX1 U3926 (.A1(N7851), .A2(N7852), .ZN(n16798));
    NANDX1 U3927 (.A1(N7853), .A2(N7854), .ZN(n16799));
    NANDX1 U3928 (.A1(N7855), .A2(N7856), .ZN(n16800));
    NOR2X1 U3929 (.A1(N7857), .A2(N7858), .ZN(N16801));
    NOR2X1 U3930 (.A1(N7859), .A2(N7860), .ZN(n16802));
    NANDX1 U3931 (.A1(N7861), .A2(N7862), .ZN(N16803));
    NANDX1 U3932 (.A1(N7863), .A2(N7864), .ZN(n16804));
    NANDX1 U3933 (.A1(N7865), .A2(N7866), .ZN(n16805));
    NOR2X1 U3934 (.A1(N7867), .A2(N7868), .ZN(N16806));
    NOR2X1 U3935 (.A1(N7869), .A2(N7870), .ZN(n16807));
    NANDX1 U3936 (.A1(N7871), .A2(N7872), .ZN(n16808));
    NANDX1 U3937 (.A1(N7873), .A2(N7874), .ZN(N16809));
    NANDX1 U3938 (.A1(N7875), .A2(N7876), .ZN(n16810));
    NANDX1 U3939 (.A1(N7877), .A2(N7878), .ZN(n16811));
    NANDX1 U3940 (.A1(N7879), .A2(N7880), .ZN(n16812));
    NOR2X1 U3941 (.A1(N7881), .A2(N7882), .ZN(n16813));
    NOR2X1 U3942 (.A1(N7883), .A2(N7884), .ZN(N16814));
    NANDX1 U3943 (.A1(N7885), .A2(N7886), .ZN(n16815));
    NANDX1 U3944 (.A1(N7887), .A2(N7888), .ZN(n16816));
    NOR2X1 U3945 (.A1(N7889), .A2(N7890), .ZN(n16817));
    NANDX1 U3946 (.A1(N7891), .A2(N7892), .ZN(N16818));
    NOR2X1 U3947 (.A1(N7893), .A2(N7894), .ZN(n16819));
    NANDX1 U3948 (.A1(N7895), .A2(N7896), .ZN(n16820));
    NANDX1 U3949 (.A1(N7897), .A2(N7898), .ZN(n16821));
    NOR2X1 U3950 (.A1(N7899), .A2(N7900), .ZN(n16822));
    NOR2X1 U3951 (.A1(N7901), .A2(N7902), .ZN(n16823));
    NANDX1 U3952 (.A1(N7903), .A2(N7904), .ZN(n16824));
    NOR2X1 U3953 (.A1(N7905), .A2(N7906), .ZN(n16825));
    NOR2X1 U3954 (.A1(N7907), .A2(N7908), .ZN(n16826));
    NANDX1 U3955 (.A1(N7909), .A2(N7910), .ZN(n16827));
    NANDX1 U3956 (.A1(N7911), .A2(N7912), .ZN(N16828));
    NANDX1 U3957 (.A1(N7913), .A2(N7914), .ZN(n16829));
    NOR2X1 U3958 (.A1(N7915), .A2(N7916), .ZN(N16830));
    NANDX1 U3959 (.A1(N7917), .A2(N7918), .ZN(n16831));
    NANDX1 U3960 (.A1(N7919), .A2(N7920), .ZN(n16832));
    NOR2X1 U3961 (.A1(N7921), .A2(N7922), .ZN(n16833));
    NOR2X1 U3962 (.A1(N7923), .A2(N7924), .ZN(n16834));
    NANDX1 U3963 (.A1(N7925), .A2(N7926), .ZN(n16835));
    NOR2X1 U3964 (.A1(N7927), .A2(N7928), .ZN(n16836));
    NOR2X1 U3965 (.A1(N7929), .A2(N7930), .ZN(n16837));
    NANDX1 U3966 (.A1(N7931), .A2(N7932), .ZN(n16838));
    NANDX1 U3967 (.A1(N7933), .A2(N7934), .ZN(N16839));
    NOR2X1 U3968 (.A1(N7935), .A2(N7936), .ZN(n16840));
    NOR2X1 U3969 (.A1(N7937), .A2(N7938), .ZN(N16841));
    NANDX1 U3970 (.A1(N7939), .A2(N7940), .ZN(n16842));
    NANDX1 U3971 (.A1(N7941), .A2(N7942), .ZN(n16843));
    NANDX1 U3972 (.A1(N7943), .A2(N7944), .ZN(n16844));
    NANDX1 U3973 (.A1(N7945), .A2(N7946), .ZN(n16845));
    NOR2X1 U3974 (.A1(N7947), .A2(N7948), .ZN(N16846));
    NOR2X1 U3975 (.A1(N7949), .A2(N7950), .ZN(N16847));
    NANDX1 U3976 (.A1(N7951), .A2(N7952), .ZN(N16848));
    NANDX1 U3977 (.A1(N7953), .A2(N7954), .ZN(n16849));
    NANDX1 U3978 (.A1(N7955), .A2(N7956), .ZN(n16850));
    NOR2X1 U3979 (.A1(N7957), .A2(N7958), .ZN(n16851));
    NANDX1 U3980 (.A1(N7959), .A2(N7960), .ZN(n16852));
    NANDX1 U3981 (.A1(N7961), .A2(N7962), .ZN(n16853));
    NOR2X1 U3982 (.A1(N7963), .A2(N7964), .ZN(N16854));
    NOR2X1 U3983 (.A1(N7965), .A2(N7966), .ZN(n16855));
    NANDX1 U3984 (.A1(N7967), .A2(N7968), .ZN(n16856));
    NOR2X1 U3985 (.A1(N7969), .A2(N7970), .ZN(n16857));
    NANDX1 U3986 (.A1(N7971), .A2(N7972), .ZN(n16858));
    NANDX1 U3987 (.A1(N7973), .A2(N7974), .ZN(n16859));
    NANDX1 U3988 (.A1(N7975), .A2(N7976), .ZN(n16860));
    NANDX1 U3989 (.A1(N7977), .A2(N7978), .ZN(n16861));
    NOR2X1 U3990 (.A1(N7979), .A2(N7980), .ZN(n16862));
    NANDX1 U3991 (.A1(N7981), .A2(N7982), .ZN(n16863));
    NANDX1 U3992 (.A1(N7983), .A2(N7984), .ZN(n16864));
    NOR2X1 U3993 (.A1(N7985), .A2(N7986), .ZN(n16865));
    NOR2X1 U3994 (.A1(N7987), .A2(N7988), .ZN(n16866));
    NANDX1 U3995 (.A1(N7989), .A2(N7990), .ZN(N16867));
    NOR2X1 U3996 (.A1(N7991), .A2(N7992), .ZN(n16868));
    NANDX1 U3997 (.A1(N7993), .A2(N7994), .ZN(n16869));
    NANDX1 U3998 (.A1(N7995), .A2(N7996), .ZN(n16870));
    NOR2X1 U3999 (.A1(N7997), .A2(N7998), .ZN(N16871));
    NOR2X1 U4000 (.A1(N7999), .A2(N8000), .ZN(n16872));
    NOR2X1 U4001 (.A1(N8001), .A2(N8002), .ZN(n16873));
    NANDX1 U4002 (.A1(N8003), .A2(N8004), .ZN(n16874));
    NANDX1 U4003 (.A1(N8005), .A2(N8006), .ZN(n16875));
    NANDX1 U4004 (.A1(N8007), .A2(N8008), .ZN(n16876));
    NOR2X1 U4005 (.A1(N8009), .A2(N8010), .ZN(n16877));
    NANDX1 U4006 (.A1(N8011), .A2(N8012), .ZN(n16878));
    NOR2X1 U4007 (.A1(N8013), .A2(N8014), .ZN(N16879));
    NANDX1 U4008 (.A1(N8015), .A2(N8016), .ZN(n16880));
    NOR2X1 U4009 (.A1(N8017), .A2(N8018), .ZN(n16881));
    NOR2X1 U4010 (.A1(N8019), .A2(N8020), .ZN(n16882));
    NOR2X1 U4011 (.A1(N8021), .A2(N8022), .ZN(N16883));
    NANDX1 U4012 (.A1(N8023), .A2(N8024), .ZN(n16884));
    NOR2X1 U4013 (.A1(N8025), .A2(N8026), .ZN(n16885));
    NOR2X1 U4014 (.A1(N8027), .A2(N8028), .ZN(n16886));
    NANDX1 U4015 (.A1(N8029), .A2(N8030), .ZN(n16887));
    NOR2X1 U4016 (.A1(N8031), .A2(N8032), .ZN(n16888));
    NANDX1 U4017 (.A1(N8033), .A2(N8034), .ZN(n16889));
    NOR2X1 U4018 (.A1(N8035), .A2(N8036), .ZN(n16890));
    NANDX1 U4019 (.A1(N8037), .A2(N8038), .ZN(N16891));
    NOR2X1 U4020 (.A1(N8039), .A2(N8040), .ZN(n16892));
    NOR2X1 U4021 (.A1(N8041), .A2(N8042), .ZN(n16893));
    NOR2X1 U4022 (.A1(N8043), .A2(N8044), .ZN(n16894));
    NOR2X1 U4023 (.A1(N8045), .A2(N8046), .ZN(n16895));
    NOR2X1 U4024 (.A1(N8047), .A2(N8048), .ZN(n16896));
    NOR2X1 U4025 (.A1(N8049), .A2(N8050), .ZN(n16897));
    NANDX1 U4026 (.A1(N8051), .A2(N8052), .ZN(n16898));
    NOR2X1 U4027 (.A1(N8053), .A2(N8054), .ZN(n16899));
    NOR2X1 U4028 (.A1(N8055), .A2(N8056), .ZN(n16900));
    NOR2X1 U4029 (.A1(N8057), .A2(N8058), .ZN(n16901));
    NANDX1 U4030 (.A1(N8059), .A2(N8060), .ZN(n16902));
    NOR2X1 U4031 (.A1(N8061), .A2(N8062), .ZN(n16903));
    NOR2X1 U4032 (.A1(N8063), .A2(N8064), .ZN(n16904));
    NOR2X1 U4033 (.A1(N8065), .A2(N8066), .ZN(n16905));
    NANDX1 U4034 (.A1(N8067), .A2(N8068), .ZN(N16906));
    NANDX1 U4035 (.A1(N8069), .A2(N8070), .ZN(n16907));
    NOR2X1 U4036 (.A1(N8071), .A2(N8072), .ZN(n16908));
    NOR2X1 U4037 (.A1(N8073), .A2(N8074), .ZN(n16909));
    NANDX1 U4038 (.A1(N8075), .A2(N8076), .ZN(n16910));
    NOR2X1 U4039 (.A1(N8077), .A2(N8078), .ZN(N16911));
    NANDX1 U4040 (.A1(N8079), .A2(N8080), .ZN(n16912));
    NANDX1 U4041 (.A1(N8081), .A2(N8082), .ZN(n16913));
    NOR2X1 U4042 (.A1(N8083), .A2(N8084), .ZN(n16914));
    NOR2X1 U4043 (.A1(N8085), .A2(N8086), .ZN(n16915));
    NANDX1 U4044 (.A1(N8087), .A2(N8088), .ZN(n16916));
    NANDX1 U4045 (.A1(N8089), .A2(N8090), .ZN(n16917));
    NANDX1 U4046 (.A1(N8091), .A2(N8092), .ZN(n16918));
    NANDX1 U4047 (.A1(N8093), .A2(N8094), .ZN(n16919));
    NOR2X1 U4048 (.A1(N8095), .A2(N8096), .ZN(N16920));
    NANDX1 U4049 (.A1(N8097), .A2(N8098), .ZN(n16921));
    NANDX1 U4050 (.A1(N8099), .A2(N8100), .ZN(n16922));
    NANDX1 U4051 (.A1(N8101), .A2(N8102), .ZN(n16923));
    NANDX1 U4052 (.A1(N8103), .A2(N8104), .ZN(n16924));
    NANDX1 U4053 (.A1(N8105), .A2(N8106), .ZN(N16925));
    NANDX1 U4054 (.A1(N8107), .A2(N8108), .ZN(n16926));
    NANDX1 U4055 (.A1(N8109), .A2(N8110), .ZN(n16927));
    NOR2X1 U4056 (.A1(N8111), .A2(N8112), .ZN(n16928));
    NOR2X1 U4057 (.A1(N8113), .A2(N8114), .ZN(n16929));
    NOR2X1 U4058 (.A1(N8115), .A2(N8116), .ZN(n16930));
    NOR2X1 U4059 (.A1(N8117), .A2(N8118), .ZN(n16931));
    NANDX1 U4060 (.A1(N8119), .A2(N8120), .ZN(n16932));
    NANDX1 U4061 (.A1(N8121), .A2(N8122), .ZN(n16933));
    NOR2X1 U4062 (.A1(N8123), .A2(N8124), .ZN(n16934));
    NANDX1 U4063 (.A1(N8125), .A2(N8126), .ZN(n16935));
    NANDX1 U4064 (.A1(N8127), .A2(N8128), .ZN(n16936));
    NANDX1 U4065 (.A1(N8129), .A2(N8130), .ZN(n16937));
    NANDX1 U4066 (.A1(N8131), .A2(N8132), .ZN(n16938));
    NOR2X1 U4067 (.A1(N8133), .A2(N8134), .ZN(N16939));
    NANDX1 U4068 (.A1(N8135), .A2(N8136), .ZN(N16940));
    NOR2X1 U4069 (.A1(N8137), .A2(N8138), .ZN(n16941));
    NOR2X1 U4070 (.A1(N8139), .A2(N8140), .ZN(N16942));
    NOR2X1 U4071 (.A1(N8141), .A2(N8142), .ZN(n16943));
    NOR2X1 U4072 (.A1(N8143), .A2(N8144), .ZN(n16944));
    NOR2X1 U4073 (.A1(N8145), .A2(N8146), .ZN(n16945));
    NANDX1 U4074 (.A1(N8147), .A2(N8148), .ZN(n16946));
    NANDX1 U4075 (.A1(N8149), .A2(N8150), .ZN(n16947));
    NANDX1 U4076 (.A1(N8151), .A2(N8152), .ZN(n16948));
    NOR2X1 U4077 (.A1(N8153), .A2(N8154), .ZN(N16949));
    NANDX1 U4078 (.A1(N8155), .A2(N8156), .ZN(n16950));
    NOR2X1 U4079 (.A1(N8157), .A2(N8158), .ZN(n16951));
    NOR2X1 U4080 (.A1(N8159), .A2(N8160), .ZN(n16952));
    NOR2X1 U4081 (.A1(N8161), .A2(N8162), .ZN(n16953));
    NANDX1 U4082 (.A1(N8163), .A2(N8164), .ZN(N16954));
    NANDX1 U4083 (.A1(N8165), .A2(N8166), .ZN(n16955));
    NANDX1 U4084 (.A1(N8167), .A2(N8168), .ZN(N16956));
    NOR2X1 U4085 (.A1(N8169), .A2(N8170), .ZN(n16957));
    NANDX1 U4086 (.A1(N8171), .A2(N8172), .ZN(n16958));
    NANDX1 U4087 (.A1(N8173), .A2(N8174), .ZN(n16959));
    NOR2X1 U4088 (.A1(N8175), .A2(N8176), .ZN(n16960));
    NANDX1 U4089 (.A1(N8177), .A2(N8178), .ZN(n16961));
    NANDX1 U4090 (.A1(N8179), .A2(N8180), .ZN(n16962));
    NANDX1 U4091 (.A1(N8181), .A2(N8182), .ZN(n16963));
    NOR2X1 U4092 (.A1(N8183), .A2(N8184), .ZN(n16964));
    NANDX1 U4093 (.A1(N8185), .A2(N8186), .ZN(n16965));
    NANDX1 U4094 (.A1(N8187), .A2(N8188), .ZN(n16966));
    NANDX1 U4095 (.A1(N8189), .A2(N8190), .ZN(n16967));
    NOR2X1 U4096 (.A1(N8191), .A2(N8192), .ZN(n16968));
    NOR2X1 U4097 (.A1(N8193), .A2(N8194), .ZN(n16969));
    NANDX1 U4098 (.A1(N8195), .A2(N8196), .ZN(n16970));
    NOR2X1 U4099 (.A1(N8197), .A2(N8198), .ZN(N16971));
    NOR2X1 U4100 (.A1(N8199), .A2(N8200), .ZN(n16972));
    NANDX1 U4101 (.A1(N8201), .A2(N8202), .ZN(n16973));
    NOR2X1 U4102 (.A1(N8203), .A2(N8204), .ZN(n16974));
    NOR2X1 U4103 (.A1(N8205), .A2(N8206), .ZN(n16975));
    NOR2X1 U4104 (.A1(N8207), .A2(N8208), .ZN(n16976));
    NANDX1 U4105 (.A1(N8209), .A2(N8210), .ZN(n16977));
    NOR2X1 U4106 (.A1(N8211), .A2(N8212), .ZN(n16978));
    NANDX1 U4107 (.A1(N8213), .A2(N8214), .ZN(n16979));
    NOR2X1 U4108 (.A1(N8215), .A2(N8216), .ZN(n16980));
    NANDX1 U4109 (.A1(N8217), .A2(N8218), .ZN(N16981));
    NANDX1 U4110 (.A1(N8219), .A2(N8220), .ZN(n16982));
    NOR2X1 U4111 (.A1(N8221), .A2(N8222), .ZN(n16983));
    NANDX1 U4112 (.A1(N8223), .A2(N8224), .ZN(N16984));
    NOR2X1 U4113 (.A1(N8225), .A2(N8226), .ZN(n16985));
    NANDX1 U4114 (.A1(N8227), .A2(N8228), .ZN(n16986));
    NOR2X1 U4115 (.A1(N8229), .A2(N8230), .ZN(n16987));
    NOR2X1 U4116 (.A1(N8231), .A2(N8232), .ZN(n16988));
    NOR2X1 U4117 (.A1(N8233), .A2(N8234), .ZN(n16989));
    NOR2X1 U4118 (.A1(N8235), .A2(N8236), .ZN(N16990));
    NANDX1 U4119 (.A1(N8237), .A2(N8238), .ZN(n16991));
    NANDX1 U4120 (.A1(N8239), .A2(N8240), .ZN(n16992));
    NANDX1 U4121 (.A1(N8241), .A2(N8242), .ZN(n16993));
    NOR2X1 U4122 (.A1(N8243), .A2(N8244), .ZN(n16994));
    NANDX1 U4123 (.A1(N8245), .A2(N8246), .ZN(n16995));
    NANDX1 U4124 (.A1(N8247), .A2(N8248), .ZN(N16996));
    NANDX1 U4125 (.A1(N8249), .A2(N8250), .ZN(n16997));
    NANDX1 U4126 (.A1(N8251), .A2(N8252), .ZN(n16998));
    NANDX1 U4127 (.A1(N8253), .A2(N8254), .ZN(N16999));
    NANDX1 U4128 (.A1(N8255), .A2(N8256), .ZN(n17000));
    NOR2X1 U4129 (.A1(N8257), .A2(N8258), .ZN(n17001));
    NANDX1 U4130 (.A1(N8259), .A2(N8260), .ZN(N17002));
    NOR2X1 U4131 (.A1(N8261), .A2(N8262), .ZN(n17003));
    NOR2X1 U4132 (.A1(N8263), .A2(N8264), .ZN(N17004));
    NOR2X1 U4133 (.A1(N8265), .A2(N8266), .ZN(n17005));
    NOR2X1 U4134 (.A1(N8267), .A2(N8268), .ZN(n17006));
    NOR2X1 U4135 (.A1(N8269), .A2(N8270), .ZN(n17007));
    NANDX1 U4136 (.A1(N8271), .A2(N8272), .ZN(n17008));
    NOR2X1 U4137 (.A1(N8273), .A2(N8274), .ZN(n17009));
    NANDX1 U4138 (.A1(N8275), .A2(N8276), .ZN(n17010));
    NANDX1 U4139 (.A1(N8277), .A2(N8278), .ZN(n17011));
    NANDX1 U4140 (.A1(N8279), .A2(N8280), .ZN(n17012));
    NANDX1 U4141 (.A1(N8281), .A2(N8282), .ZN(n17013));
    NANDX1 U4142 (.A1(N8283), .A2(N8284), .ZN(n17014));
    NOR2X1 U4143 (.A1(N8285), .A2(N8286), .ZN(n17015));
    NANDX1 U4144 (.A1(N8287), .A2(N8288), .ZN(n17016));
    NANDX1 U4145 (.A1(N8289), .A2(N8290), .ZN(N17017));
    NANDX1 U4146 (.A1(N8291), .A2(N8292), .ZN(N17018));
    NOR2X1 U4147 (.A1(N8293), .A2(N8294), .ZN(N17019));
    NANDX1 U4148 (.A1(N8295), .A2(N8296), .ZN(n17020));
    NANDX1 U4149 (.A1(N8297), .A2(N8298), .ZN(n17021));
    NANDX1 U4150 (.A1(N8299), .A2(N8300), .ZN(n17022));
    NANDX1 U4151 (.A1(N8301), .A2(N8302), .ZN(n17023));
    NOR2X1 U4152 (.A1(N8303), .A2(N8304), .ZN(N17024));
    NANDX1 U4153 (.A1(N8305), .A2(N8306), .ZN(n17025));
    NOR2X1 U4154 (.A1(N8307), .A2(N8308), .ZN(n17026));
    NANDX1 U4155 (.A1(N8309), .A2(N8310), .ZN(n17027));
    NANDX1 U4156 (.A1(N8311), .A2(N8312), .ZN(n17028));
    NANDX1 U4157 (.A1(N8313), .A2(N8314), .ZN(n17029));
    NANDX1 U4158 (.A1(N8315), .A2(N8316), .ZN(n17030));
    NOR2X1 U4159 (.A1(N8317), .A2(N8318), .ZN(n17031));
    NOR2X1 U4160 (.A1(N8319), .A2(N8320), .ZN(n17032));
    NOR2X1 U4161 (.A1(N8321), .A2(N8322), .ZN(n17033));
    NOR2X1 U4162 (.A1(N8323), .A2(N8324), .ZN(n17034));
    NOR2X1 U4163 (.A1(N8325), .A2(N8326), .ZN(n17035));
    NOR2X1 U4164 (.A1(N8327), .A2(N8328), .ZN(n17036));
    NANDX1 U4165 (.A1(N8329), .A2(N8330), .ZN(n17037));
    NOR2X1 U4166 (.A1(N8331), .A2(N8332), .ZN(n17038));
    NOR2X1 U4167 (.A1(N8333), .A2(N8334), .ZN(n17039));
    NANDX1 U4168 (.A1(N8335), .A2(N8336), .ZN(n17040));
    NANDX1 U4169 (.A1(N8337), .A2(N8338), .ZN(N17041));
    NANDX1 U4170 (.A1(N8339), .A2(N8340), .ZN(n17042));
    NANDX1 U4171 (.A1(N8341), .A2(N8342), .ZN(N17043));
    NOR2X1 U4172 (.A1(N8343), .A2(N8344), .ZN(n17044));
    NANDX1 U4173 (.A1(N8345), .A2(N8346), .ZN(n17045));
    NANDX1 U4174 (.A1(N8347), .A2(N8348), .ZN(n17046));
    NOR2X1 U4175 (.A1(N8349), .A2(N8350), .ZN(n17047));
    NOR2X1 U4176 (.A1(N8351), .A2(N8352), .ZN(n17048));
    NOR2X1 U4177 (.A1(N8353), .A2(N8354), .ZN(n17049));
    NOR2X1 U4178 (.A1(N8355), .A2(N8356), .ZN(n17050));
    NANDX1 U4179 (.A1(N8357), .A2(N8358), .ZN(n17051));
    NANDX1 U4180 (.A1(N8359), .A2(N8360), .ZN(N17052));
    NANDX1 U4181 (.A1(N8361), .A2(N8362), .ZN(N17053));
    NOR2X1 U4182 (.A1(N8363), .A2(N8364), .ZN(n17054));
    NOR2X1 U4183 (.A1(N8365), .A2(N8366), .ZN(n17055));
    NOR2X1 U4184 (.A1(N8367), .A2(N8368), .ZN(n17056));
    NANDX1 U4185 (.A1(N8369), .A2(N8370), .ZN(n17057));
    NANDX1 U4186 (.A1(N8371), .A2(N8372), .ZN(n17058));
    NANDX1 U4187 (.A1(N8373), .A2(N8374), .ZN(n17059));
    NOR2X1 U4188 (.A1(N8375), .A2(N8376), .ZN(n17060));
    NOR2X1 U4189 (.A1(N8377), .A2(N8378), .ZN(n17061));
    NOR2X1 U4190 (.A1(N8379), .A2(N8380), .ZN(n17062));
    NOR2X1 U4191 (.A1(N8381), .A2(N8382), .ZN(N17063));
    NANDX1 U4192 (.A1(N8383), .A2(N8384), .ZN(n17064));
    NOR2X1 U4193 (.A1(N8385), .A2(N8386), .ZN(n17065));
    NOR2X1 U4194 (.A1(N8387), .A2(N8388), .ZN(N17066));
    NANDX1 U4195 (.A1(N8389), .A2(N8390), .ZN(n17067));
    NANDX1 U4196 (.A1(N8391), .A2(N8392), .ZN(n17068));
    NOR2X1 U4197 (.A1(N8393), .A2(N8394), .ZN(n17069));
    NANDX1 U4198 (.A1(N8395), .A2(N8396), .ZN(n17070));
    NANDX1 U4199 (.A1(N8397), .A2(N8398), .ZN(n17071));
    NOR2X1 U4200 (.A1(N8399), .A2(N8400), .ZN(n17072));
    NANDX1 U4201 (.A1(N8401), .A2(N8402), .ZN(n17073));
    NOR2X1 U4202 (.A1(N8403), .A2(N8404), .ZN(n17074));
    NOR2X1 U4203 (.A1(N8405), .A2(N8406), .ZN(n17075));
    NOR2X1 U4204 (.A1(N8407), .A2(N8408), .ZN(N17076));
    NANDX1 U4205 (.A1(N8409), .A2(N8410), .ZN(n17077));
    NOR2X1 U4206 (.A1(N8411), .A2(N8412), .ZN(n17078));
    NOR2X1 U4207 (.A1(N8413), .A2(N8414), .ZN(n17079));
    NOR2X1 U4208 (.A1(N8415), .A2(N8416), .ZN(n17080));
    NOR2X1 U4209 (.A1(N8417), .A2(N8418), .ZN(n17081));
    NANDX1 U4210 (.A1(N8419), .A2(N8420), .ZN(N17082));
    NANDX1 U4211 (.A1(N8421), .A2(N8422), .ZN(N17083));
    NANDX1 U4212 (.A1(N8423), .A2(N8424), .ZN(n17084));
    NOR2X1 U4213 (.A1(N8425), .A2(N8426), .ZN(n17085));
    NANDX1 U4214 (.A1(N8427), .A2(N8428), .ZN(n17086));
    NOR2X1 U4215 (.A1(N8429), .A2(N8430), .ZN(n17087));
    NANDX1 U4216 (.A1(N8431), .A2(N8432), .ZN(n17088));
    NANDX1 U4217 (.A1(N8433), .A2(N8434), .ZN(n17089));
    NANDX1 U4218 (.A1(N8435), .A2(N8436), .ZN(n17090));
    NANDX1 U4219 (.A1(N8437), .A2(N8438), .ZN(N17091));
    NANDX1 U4220 (.A1(N8439), .A2(N8440), .ZN(n17092));
    NANDX1 U4221 (.A1(N8441), .A2(N8442), .ZN(n17093));
    NOR2X1 U4222 (.A1(N8443), .A2(N8444), .ZN(n17094));
    NOR2X1 U4223 (.A1(N8445), .A2(N8446), .ZN(N17095));
    NOR2X1 U4224 (.A1(N8447), .A2(N8448), .ZN(n17096));
    NOR2X1 U4225 (.A1(N8449), .A2(N8450), .ZN(n17097));
    NOR2X1 U4226 (.A1(N8451), .A2(N8452), .ZN(N17098));
    NANDX1 U4227 (.A1(N8453), .A2(N8454), .ZN(n17099));
    NANDX1 U4228 (.A1(N8455), .A2(N8456), .ZN(n17100));
    NANDX1 U4229 (.A1(N8457), .A2(N8458), .ZN(n17101));
    NOR2X1 U4230 (.A1(N8459), .A2(N8460), .ZN(N17102));
    NANDX1 U4231 (.A1(N8461), .A2(N8462), .ZN(n17103));
    NOR2X1 U4232 (.A1(N8463), .A2(N8464), .ZN(n17104));
    NOR2X1 U4233 (.A1(N8465), .A2(N8466), .ZN(n17105));
    NANDX1 U4234 (.A1(N8467), .A2(N8468), .ZN(N17106));
    NOR2X1 U4235 (.A1(N8469), .A2(N8470), .ZN(N17107));
    NOR2X1 U4236 (.A1(N8471), .A2(N8472), .ZN(n17108));
    NOR2X1 U4237 (.A1(N8473), .A2(N8474), .ZN(n17109));
    NOR2X1 U4238 (.A1(N8475), .A2(N8476), .ZN(N17110));
    NOR2X1 U4239 (.A1(N8477), .A2(N8478), .ZN(n17111));
    NOR2X1 U4240 (.A1(N8479), .A2(N8480), .ZN(n17112));
    NOR2X1 U4241 (.A1(N8481), .A2(N8482), .ZN(n17113));
    NANDX1 U4242 (.A1(N8483), .A2(N8484), .ZN(n17114));
    NOR2X1 U4243 (.A1(N8485), .A2(N8486), .ZN(N17115));
    NOR2X1 U4244 (.A1(N8487), .A2(N8488), .ZN(n17116));
    NANDX1 U4245 (.A1(N8489), .A2(N8490), .ZN(n17117));
    NOR2X1 U4246 (.A1(N8491), .A2(N8492), .ZN(n17118));
    NANDX1 U4247 (.A1(N8493), .A2(N8494), .ZN(n17119));
    NOR2X1 U4248 (.A1(N8495), .A2(N8496), .ZN(n17120));
    NANDX1 U4249 (.A1(N8497), .A2(N8498), .ZN(n17121));
    NOR2X1 U4250 (.A1(N8499), .A2(N8500), .ZN(n17122));
    NANDX1 U4251 (.A1(N8501), .A2(N8502), .ZN(n17123));
    NANDX1 U4252 (.A1(N8503), .A2(N8504), .ZN(N17124));
    NOR2X1 U4253 (.A1(N8505), .A2(N8506), .ZN(n17125));
    NOR2X1 U4254 (.A1(N8507), .A2(N8508), .ZN(n17126));
    NANDX1 U4255 (.A1(N8509), .A2(N8510), .ZN(N17127));
    NANDX1 U4256 (.A1(N8511), .A2(N8512), .ZN(n17128));
    NOR2X1 U4257 (.A1(N8513), .A2(N8514), .ZN(n17129));
    NOR2X1 U4258 (.A1(N8515), .A2(N8516), .ZN(n17130));
    NOR2X1 U4259 (.A1(N8517), .A2(N8518), .ZN(n17131));
    NANDX1 U4260 (.A1(N8519), .A2(N8520), .ZN(n17132));
    NANDX1 U4261 (.A1(N8521), .A2(N8522), .ZN(n17133));
    NANDX1 U4262 (.A1(N8523), .A2(N8524), .ZN(n17134));
    NOR2X1 U4263 (.A1(N8525), .A2(N8526), .ZN(n17135));
    NANDX1 U4264 (.A1(N8527), .A2(N8528), .ZN(n17136));
    NOR2X1 U4265 (.A1(N8529), .A2(N8530), .ZN(n17137));
    NOR2X1 U4266 (.A1(N8531), .A2(N8532), .ZN(n17138));
    NANDX1 U4267 (.A1(N8533), .A2(N8534), .ZN(n17139));
    NOR2X1 U4268 (.A1(N8535), .A2(N8536), .ZN(n17140));
    NANDX1 U4269 (.A1(N8537), .A2(N8538), .ZN(N17141));
    NANDX1 U4270 (.A1(N8539), .A2(N8540), .ZN(n17142));
    NANDX1 U4271 (.A1(N8541), .A2(N8542), .ZN(n17143));
    NANDX1 U4272 (.A1(N8543), .A2(N8544), .ZN(n17144));
    NANDX1 U4273 (.A1(N8545), .A2(N8546), .ZN(n17145));
    NANDX1 U4274 (.A1(N8547), .A2(N8548), .ZN(n17146));
    NANDX1 U4275 (.A1(N8549), .A2(N8550), .ZN(n17147));
    NOR2X1 U4276 (.A1(N8551), .A2(N8552), .ZN(N17148));
    NANDX1 U4277 (.A1(N8553), .A2(N8554), .ZN(n17149));
    NOR2X1 U4278 (.A1(N8555), .A2(N8556), .ZN(n17150));
    NOR2X1 U4279 (.A1(N8557), .A2(N8558), .ZN(n17151));
    NOR2X1 U4280 (.A1(N8559), .A2(N8560), .ZN(n17152));
    NOR2X1 U4281 (.A1(N8561), .A2(N8562), .ZN(n17153));
    NANDX1 U4282 (.A1(N8563), .A2(N8564), .ZN(n17154));
    NANDX1 U4283 (.A1(N8565), .A2(N8566), .ZN(n17155));
    NANDX1 U4284 (.A1(N8567), .A2(N8568), .ZN(N17156));
    NANDX1 U4285 (.A1(N8569), .A2(N8570), .ZN(n17157));
    NOR2X1 U4286 (.A1(N8571), .A2(N8572), .ZN(n17158));
    NOR2X1 U4287 (.A1(N8573), .A2(N8574), .ZN(n17159));
    NANDX1 U4288 (.A1(N8575), .A2(N8576), .ZN(n17160));
    NANDX1 U4289 (.A1(N8577), .A2(N8578), .ZN(n17161));
    NOR2X1 U4290 (.A1(N8579), .A2(N8580), .ZN(n17162));
    NANDX1 U4291 (.A1(N8581), .A2(N8582), .ZN(n17163));
    NOR2X1 U4292 (.A1(N8583), .A2(N8584), .ZN(n17164));
    NANDX1 U4293 (.A1(N8585), .A2(N8586), .ZN(n17165));
    NANDX1 U4294 (.A1(N8587), .A2(N8588), .ZN(n17166));
    NANDX1 U4295 (.A1(N8589), .A2(N8590), .ZN(n17167));
    NANDX1 U4296 (.A1(N8591), .A2(N8592), .ZN(n17168));
    NANDX1 U4297 (.A1(N8593), .A2(N8594), .ZN(N17169));
    NANDX1 U4298 (.A1(N8595), .A2(N8596), .ZN(n17170));
    NOR2X1 U4299 (.A1(N8597), .A2(N8598), .ZN(n17171));
    NOR2X1 U4300 (.A1(N8599), .A2(N8600), .ZN(n17172));
    NOR2X1 U4301 (.A1(N8601), .A2(N8602), .ZN(n17173));
    NANDX1 U4302 (.A1(N8603), .A2(N8604), .ZN(n17174));
    NANDX1 U4303 (.A1(N8605), .A2(N8606), .ZN(n17175));
    NANDX1 U4304 (.A1(N8607), .A2(N8608), .ZN(n17176));
    NOR2X1 U4305 (.A1(N8609), .A2(N8610), .ZN(n17177));
    NOR2X1 U4306 (.A1(N8611), .A2(N8612), .ZN(n17178));
    NANDX1 U4307 (.A1(N8613), .A2(N8614), .ZN(n17179));
    NANDX1 U4308 (.A1(N8615), .A2(N8616), .ZN(n17180));
    NOR2X1 U4309 (.A1(N8617), .A2(N8618), .ZN(N17181));
    NANDX1 U4310 (.A1(N8619), .A2(N8620), .ZN(N17182));
    NANDX1 U4311 (.A1(N8621), .A2(N8622), .ZN(N17183));
    NANDX1 U4312 (.A1(N8623), .A2(N8624), .ZN(n17184));
    NANDX1 U4313 (.A1(N8625), .A2(N8626), .ZN(n17185));
    NANDX1 U4314 (.A1(N8627), .A2(N8628), .ZN(n17186));
    NOR2X1 U4315 (.A1(N8629), .A2(N8630), .ZN(n17187));
    NOR2X1 U4316 (.A1(N8631), .A2(N8632), .ZN(N17188));
    NANDX1 U4317 (.A1(N8633), .A2(N8634), .ZN(n17189));
    NOR2X1 U4318 (.A1(N8635), .A2(N8636), .ZN(n17190));
    NOR2X1 U4319 (.A1(N8637), .A2(N8638), .ZN(N17191));
    NOR2X1 U4320 (.A1(N8639), .A2(N8640), .ZN(n17192));
    NOR2X1 U4321 (.A1(N8641), .A2(N8642), .ZN(N17193));
    NANDX1 U4322 (.A1(N8643), .A2(N8644), .ZN(n17194));
    NOR2X1 U4323 (.A1(N8645), .A2(N8646), .ZN(n17195));
    NANDX1 U4324 (.A1(N8647), .A2(N8648), .ZN(n17196));
    NOR2X1 U4325 (.A1(N8649), .A2(N8650), .ZN(n17197));
    NOR2X1 U4326 (.A1(N8651), .A2(N8652), .ZN(n17198));
    NOR2X1 U4327 (.A1(N8653), .A2(N8654), .ZN(n17199));
    NANDX1 U4328 (.A1(N8655), .A2(N8656), .ZN(n17200));
    NANDX1 U4329 (.A1(N8657), .A2(N8658), .ZN(n17201));
    NOR2X1 U4330 (.A1(N8659), .A2(N8660), .ZN(n17202));
    NOR2X1 U4331 (.A1(N8661), .A2(N8662), .ZN(N17203));
    NANDX1 U4332 (.A1(N8663), .A2(N8664), .ZN(n17204));
    NANDX1 U4333 (.A1(N8665), .A2(N8666), .ZN(n17205));
    NANDX1 U4334 (.A1(N8667), .A2(N8668), .ZN(n17206));
    NANDX1 U4335 (.A1(N8669), .A2(N8670), .ZN(n17207));
    NANDX1 U4336 (.A1(N8671), .A2(N8672), .ZN(n17208));
    NOR2X1 U4337 (.A1(N8673), .A2(N8674), .ZN(N17209));
    NOR2X1 U4338 (.A1(N8675), .A2(N8676), .ZN(N17210));
    NOR2X1 U4339 (.A1(N8677), .A2(N8678), .ZN(n17211));
    NOR2X1 U4340 (.A1(N8679), .A2(N8680), .ZN(n17212));
    NOR2X1 U4341 (.A1(N8681), .A2(N8682), .ZN(n17213));
    NOR2X1 U4342 (.A1(N8683), .A2(N8684), .ZN(N17214));
    NANDX1 U4343 (.A1(N8685), .A2(N8686), .ZN(n17215));
    NANDX1 U4344 (.A1(N8687), .A2(N8688), .ZN(N17216));
    NANDX1 U4345 (.A1(N8689), .A2(N8690), .ZN(n17217));
    NANDX1 U4346 (.A1(N8691), .A2(N8692), .ZN(n17218));
    NANDX1 U4347 (.A1(N8693), .A2(N8694), .ZN(N17219));
    NOR2X1 U4348 (.A1(N8695), .A2(N8696), .ZN(n17220));
    NANDX1 U4349 (.A1(N8697), .A2(N8698), .ZN(N17221));
    NANDX1 U4350 (.A1(N8699), .A2(N8700), .ZN(n17222));
    NANDX1 U4351 (.A1(N8701), .A2(N8702), .ZN(N17223));
    NANDX1 U4352 (.A1(N8703), .A2(N8704), .ZN(n17224));
    NOR2X1 U4353 (.A1(N8705), .A2(N8706), .ZN(n17225));
    NANDX1 U4354 (.A1(N8707), .A2(N8708), .ZN(n17226));
    NOR2X1 U4355 (.A1(N8709), .A2(N8710), .ZN(n17227));
    NOR2X1 U4356 (.A1(N8711), .A2(N8712), .ZN(n17228));
    NANDX1 U4357 (.A1(N8713), .A2(N8714), .ZN(n17229));
    NANDX1 U4358 (.A1(N8715), .A2(N8716), .ZN(n17230));
    NOR2X1 U4359 (.A1(N8717), .A2(N8718), .ZN(n17231));
    NOR2X1 U4360 (.A1(N8719), .A2(N8720), .ZN(n17232));
    NANDX1 U4361 (.A1(N8721), .A2(N8722), .ZN(n17233));
    NOR2X1 U4362 (.A1(N8723), .A2(N8724), .ZN(n17234));
    NOR2X1 U4363 (.A1(N8725), .A2(N8726), .ZN(n17235));
    NANDX1 U4364 (.A1(N8727), .A2(N8728), .ZN(N17236));
    NANDX1 U4365 (.A1(N8729), .A2(N8730), .ZN(n17237));
    NANDX1 U4366 (.A1(N8731), .A2(N8732), .ZN(n17238));
    NOR2X1 U4367 (.A1(N8733), .A2(N8734), .ZN(n17239));
    NANDX1 U4368 (.A1(N8735), .A2(N8736), .ZN(n17240));
    NANDX1 U4369 (.A1(N8737), .A2(N8738), .ZN(n17241));
    NANDX1 U4370 (.A1(N8739), .A2(N8740), .ZN(n17242));
    NOR2X1 U4371 (.A1(N8741), .A2(N8742), .ZN(N17243));
    NANDX1 U4372 (.A1(N8743), .A2(N8744), .ZN(n17244));
    NANDX1 U4373 (.A1(N8745), .A2(N8746), .ZN(n17245));
    NANDX1 U4374 (.A1(N8747), .A2(N8748), .ZN(n17246));
    NOR2X1 U4375 (.A1(N8749), .A2(N8750), .ZN(n17247));
    NOR2X1 U4376 (.A1(N8751), .A2(N8752), .ZN(n17248));
    NANDX1 U4377 (.A1(N8753), .A2(N8754), .ZN(n17249));
    NOR2X1 U4378 (.A1(N8755), .A2(N8756), .ZN(N17250));
    NOR2X1 U4379 (.A1(N8757), .A2(N8758), .ZN(N17251));
    NOR2X1 U4380 (.A1(N8759), .A2(N8760), .ZN(N17252));
    NANDX1 U4381 (.A1(N8761), .A2(N8762), .ZN(n17253));
    NANDX1 U4382 (.A1(N8763), .A2(N8764), .ZN(n17254));
    NOR2X1 U4383 (.A1(N8765), .A2(N8766), .ZN(N17255));
    NOR2X1 U4384 (.A1(N8767), .A2(N8768), .ZN(n17256));
    NANDX1 U4385 (.A1(N8769), .A2(N8770), .ZN(n17257));
    NOR2X1 U4386 (.A1(N8771), .A2(N8772), .ZN(n17258));
    NOR2X1 U4387 (.A1(N8773), .A2(N8774), .ZN(n17259));
    NOR2X1 U4388 (.A1(N8775), .A2(N8776), .ZN(N17260));
    NANDX1 U4389 (.A1(N8777), .A2(N8778), .ZN(n17261));
    NOR2X1 U4390 (.A1(N8779), .A2(N8780), .ZN(n17262));
    NANDX1 U4391 (.A1(N8781), .A2(N8782), .ZN(n17263));
    NANDX1 U4392 (.A1(N8783), .A2(N8784), .ZN(N17264));
    NOR2X1 U4393 (.A1(N8785), .A2(N8786), .ZN(n17265));
    NANDX1 U4394 (.A1(N8787), .A2(N8788), .ZN(n17266));
    NOR2X1 U4395 (.A1(N8789), .A2(N8790), .ZN(n17267));
    NOR2X1 U4396 (.A1(N8791), .A2(N8792), .ZN(n17268));
    NOR2X1 U4397 (.A1(N8793), .A2(N8794), .ZN(n17269));
    NOR2X1 U4398 (.A1(N8795), .A2(N8796), .ZN(n17270));
    NANDX1 U4399 (.A1(N8797), .A2(N8798), .ZN(n17271));
    NANDX1 U4400 (.A1(N8799), .A2(N8800), .ZN(n17272));
    NANDX1 U4401 (.A1(N8801), .A2(N8802), .ZN(n17273));
    NANDX1 U4402 (.A1(N8803), .A2(N8804), .ZN(N17274));
    NANDX1 U4403 (.A1(N8805), .A2(N8806), .ZN(n17275));
    NOR2X1 U4404 (.A1(N8807), .A2(N8808), .ZN(n17276));
    NANDX1 U4405 (.A1(N8809), .A2(N8810), .ZN(n17277));
    NANDX1 U4406 (.A1(N8811), .A2(N8812), .ZN(N17278));
    NOR2X1 U4407 (.A1(N8813), .A2(N8814), .ZN(n17279));
    NOR2X1 U4408 (.A1(N8815), .A2(N8816), .ZN(n17280));
    NANDX1 U4409 (.A1(N8817), .A2(N8818), .ZN(n17281));
    NANDX1 U4410 (.A1(N8819), .A2(N8820), .ZN(n17282));
    NOR2X1 U4411 (.A1(N8821), .A2(N8822), .ZN(n17283));
    NANDX1 U4412 (.A1(N8823), .A2(N8824), .ZN(n17284));
    NOR2X1 U4413 (.A1(N8825), .A2(N8826), .ZN(N17285));
    NOR2X1 U4414 (.A1(N8827), .A2(N8828), .ZN(n17286));
    NANDX1 U4415 (.A1(N8829), .A2(N8830), .ZN(n17287));
    NANDX1 U4416 (.A1(N8831), .A2(N8832), .ZN(n17288));
    NANDX1 U4417 (.A1(N8833), .A2(N8834), .ZN(n17289));
    NANDX1 U4418 (.A1(N8835), .A2(N8836), .ZN(n17290));
    NOR2X1 U4419 (.A1(N8837), .A2(N8838), .ZN(N17291));
    NOR2X1 U4420 (.A1(N8839), .A2(N8840), .ZN(n17292));
    NOR2X1 U4421 (.A1(N8841), .A2(N8842), .ZN(n17293));
    NANDX1 U4422 (.A1(N8843), .A2(N8844), .ZN(n17294));
    NANDX1 U4423 (.A1(N8845), .A2(N8846), .ZN(n17295));
    NOR2X1 U4424 (.A1(N8847), .A2(N8848), .ZN(n17296));
    NOR2X1 U4425 (.A1(N8849), .A2(N8850), .ZN(n17297));
    NANDX1 U4426 (.A1(N8851), .A2(N8852), .ZN(n17298));
    NOR2X1 U4427 (.A1(N8853), .A2(N8854), .ZN(n17299));
    NOR2X1 U4428 (.A1(N8855), .A2(N8856), .ZN(n17300));
    NOR2X1 U4429 (.A1(N8857), .A2(N8858), .ZN(N17301));
    NOR2X1 U4430 (.A1(N8859), .A2(N8860), .ZN(n17302));
    NANDX1 U4431 (.A1(N8861), .A2(N8862), .ZN(n17303));
    NANDX1 U4432 (.A1(N8863), .A2(N8864), .ZN(N17304));
    NANDX1 U4433 (.A1(N8865), .A2(N8866), .ZN(n17305));
    NOR2X1 U4434 (.A1(N8867), .A2(N8868), .ZN(n17306));
    NOR2X1 U4435 (.A1(N8869), .A2(N8870), .ZN(n17307));
    NOR2X1 U4436 (.A1(N8871), .A2(N8872), .ZN(n17308));
    NOR2X1 U4437 (.A1(N8873), .A2(N8874), .ZN(n17309));
    NOR2X1 U4438 (.A1(N8875), .A2(N8876), .ZN(N17310));
    NOR2X1 U4439 (.A1(N8877), .A2(N8878), .ZN(n17311));
    NANDX1 U4440 (.A1(N8879), .A2(N8880), .ZN(n17312));
    NANDX1 U4441 (.A1(N8881), .A2(N8882), .ZN(n17313));
    NANDX1 U4442 (.A1(N8883), .A2(N8884), .ZN(n17314));
    NOR2X1 U4443 (.A1(N8885), .A2(N8886), .ZN(n17315));
    NOR2X1 U4444 (.A1(N8887), .A2(N8888), .ZN(n17316));
    NANDX1 U4445 (.A1(N8889), .A2(N8890), .ZN(n17317));
    NANDX1 U4446 (.A1(N8891), .A2(N8892), .ZN(N17318));
    NANDX1 U4447 (.A1(N8893), .A2(N8894), .ZN(n17319));
    NOR2X1 U4448 (.A1(N8895), .A2(N8896), .ZN(n17320));
    NANDX1 U4449 (.A1(N8897), .A2(N8898), .ZN(n17321));
    NANDX1 U4450 (.A1(N8899), .A2(N8900), .ZN(n17322));
    NANDX1 U4451 (.A1(N8901), .A2(N8902), .ZN(N17323));
    NANDX1 U4452 (.A1(N8903), .A2(N8904), .ZN(n17324));
    NOR2X1 U4453 (.A1(N8905), .A2(N8906), .ZN(n17325));
    NOR2X1 U4454 (.A1(N8907), .A2(N8908), .ZN(n17326));
    NANDX1 U4455 (.A1(N8909), .A2(N8910), .ZN(n17327));
    NOR2X1 U4456 (.A1(N8911), .A2(N8912), .ZN(n17328));
    NOR2X1 U4457 (.A1(N8913), .A2(N8914), .ZN(n17329));
    NOR2X1 U4458 (.A1(N8915), .A2(N8916), .ZN(n17330));
    NOR2X1 U4459 (.A1(N8917), .A2(N8918), .ZN(n17331));
    NOR2X1 U4460 (.A1(N8919), .A2(N8920), .ZN(n17332));
    NOR2X1 U4461 (.A1(N8921), .A2(N8922), .ZN(n17333));
    NOR2X1 U4462 (.A1(N8923), .A2(N8924), .ZN(n17334));
    NANDX1 U4463 (.A1(N8925), .A2(N8926), .ZN(N17335));
    NANDX1 U4464 (.A1(N8927), .A2(N8928), .ZN(n17336));
    NOR2X1 U4465 (.A1(N8929), .A2(N8930), .ZN(N17337));
    NANDX1 U4466 (.A1(N8931), .A2(N8932), .ZN(n17338));
    NOR2X1 U4467 (.A1(N8933), .A2(N8934), .ZN(n17339));
    NOR2X1 U4468 (.A1(N8935), .A2(N8936), .ZN(n17340));
    NOR2X1 U4469 (.A1(N8937), .A2(N8938), .ZN(n17341));
    NOR2X1 U4470 (.A1(N8939), .A2(N8940), .ZN(N17342));
    NOR2X1 U4471 (.A1(N8941), .A2(N8942), .ZN(n17343));
    NANDX1 U4472 (.A1(N8943), .A2(N8944), .ZN(n17344));
    NANDX1 U4473 (.A1(N8945), .A2(N8946), .ZN(n17345));
    NOR2X1 U4474 (.A1(N8947), .A2(N8948), .ZN(n17346));
    NANDX1 U4475 (.A1(N8949), .A2(N8950), .ZN(n17347));
    NANDX1 U4476 (.A1(N8951), .A2(N8952), .ZN(n17348));
    NOR2X1 U4477 (.A1(N8953), .A2(N8954), .ZN(n17349));
    NANDX1 U4478 (.A1(N8955), .A2(N8956), .ZN(n17350));
    NANDX1 U4479 (.A1(N8957), .A2(N8958), .ZN(n17351));
    NANDX1 U4480 (.A1(N8959), .A2(N8960), .ZN(n17352));
    NOR2X1 U4481 (.A1(N8961), .A2(N8962), .ZN(n17353));
    NOR2X1 U4482 (.A1(N8963), .A2(N8964), .ZN(n17354));
    NOR2X1 U4483 (.A1(N8965), .A2(N8966), .ZN(n17355));
    NANDX1 U4484 (.A1(N8967), .A2(N8968), .ZN(n17356));
    NANDX1 U4485 (.A1(N8969), .A2(N8970), .ZN(n17357));
    NANDX1 U4486 (.A1(N8971), .A2(N8972), .ZN(n17358));
    NANDX1 U4487 (.A1(N8973), .A2(N8974), .ZN(n17359));
    NANDX1 U4488 (.A1(N8975), .A2(N8976), .ZN(N17360));
    NANDX1 U4489 (.A1(N8977), .A2(N8978), .ZN(n17361));
    NOR2X1 U4490 (.A1(N8979), .A2(N8980), .ZN(N17362));
    NANDX1 U4491 (.A1(N8981), .A2(N8982), .ZN(n17363));
    NANDX1 U4492 (.A1(N8983), .A2(N8984), .ZN(n17364));
    NOR2X1 U4493 (.A1(N8985), .A2(N8986), .ZN(n17365));
    NOR2X1 U4494 (.A1(N8987), .A2(N8988), .ZN(n17366));
    NANDX1 U4495 (.A1(N8989), .A2(N8990), .ZN(N17367));
    NOR2X1 U4496 (.A1(N8991), .A2(N8992), .ZN(n17368));
    NOR2X1 U4497 (.A1(N8993), .A2(N8994), .ZN(N17369));
    NANDX1 U4498 (.A1(N8995), .A2(N8996), .ZN(n17370));
    NANDX1 U4499 (.A1(N8997), .A2(N8998), .ZN(n17371));
    NOR2X1 U4500 (.A1(N8999), .A2(N9000), .ZN(n17372));
    NANDX1 U4501 (.A1(N9001), .A2(N9002), .ZN(n17373));
    NANDX1 U4502 (.A1(N9003), .A2(N9004), .ZN(n17374));
    NANDX1 U4503 (.A1(N9005), .A2(N9006), .ZN(N17375));
    NANDX1 U4504 (.A1(N9007), .A2(N9008), .ZN(n17376));
    NANDX1 U4505 (.A1(N9009), .A2(N9010), .ZN(n17377));
    NANDX1 U4506 (.A1(N9011), .A2(N9012), .ZN(n17378));
    NOR2X1 U4507 (.A1(N9013), .A2(N9014), .ZN(n17379));
    NANDX1 U4508 (.A1(N9015), .A2(N9016), .ZN(n17380));
    NOR2X1 U4509 (.A1(N9017), .A2(N9018), .ZN(n17381));
    NANDX1 U4510 (.A1(N9019), .A2(N9020), .ZN(n17382));
    NOR2X1 U4511 (.A1(N9021), .A2(N9022), .ZN(n17383));
    NOR2X1 U4512 (.A1(N9023), .A2(N9024), .ZN(N17384));
    NOR2X1 U4513 (.A1(N9025), .A2(N9026), .ZN(n17385));
    NOR2X1 U4514 (.A1(N9027), .A2(N9028), .ZN(n17386));
    INVX1 U4515 (.I(N9029), .ZN(n17387));
    INVX1 U4516 (.I(N9030), .ZN(n17388));
    INVX1 U4517 (.I(N9031), .ZN(n17389));
    INVX1 U4518 (.I(N9032), .ZN(n17390));
    INVX1 U4519 (.I(N9033), .ZN(n17391));
    INVX1 U4520 (.I(N9034), .ZN(n17392));
    INVX1 U4521 (.I(N9035), .ZN(N17393));
    INVX1 U4522 (.I(N9036), .ZN(n17394));
    INVX1 U4523 (.I(N9037), .ZN(n17395));
    INVX1 U4524 (.I(N9038), .ZN(n17396));
    INVX1 U4525 (.I(N9039), .ZN(N17397));
    INVX1 U4526 (.I(N9040), .ZN(n17398));
    INVX1 U4527 (.I(N9041), .ZN(N17399));
    INVX1 U4528 (.I(N9042), .ZN(N17400));
    INVX1 U4529 (.I(N9043), .ZN(n17401));
    INVX1 U4530 (.I(N9044), .ZN(n17402));
    INVX1 U4531 (.I(N9045), .ZN(n17403));
    INVX1 U4532 (.I(N9046), .ZN(n17404));
    INVX1 U4533 (.I(N9047), .ZN(n17405));
    INVX1 U4534 (.I(N9048), .ZN(n17406));
    INVX1 U4535 (.I(N9049), .ZN(n17407));
    INVX1 U4536 (.I(N9050), .ZN(n17408));
    INVX1 U4537 (.I(N9051), .ZN(n17409));
    INVX1 U4538 (.I(N9052), .ZN(n17410));
    INVX1 U4539 (.I(N9053), .ZN(n17411));
    INVX1 U4540 (.I(N9054), .ZN(n17412));
    INVX1 U4541 (.I(N9055), .ZN(N17413));
    INVX1 U4542 (.I(N9056), .ZN(n17414));
    INVX1 U4543 (.I(N9057), .ZN(n17415));
    INVX1 U4544 (.I(N9058), .ZN(n17416));
    INVX1 U4545 (.I(N9059), .ZN(n17417));
    INVX1 U4546 (.I(N9060), .ZN(n17418));
    INVX1 U4547 (.I(N9061), .ZN(n17419));
    INVX1 U4548 (.I(N9062), .ZN(n17420));
    INVX1 U4549 (.I(N9063), .ZN(n17421));
    INVX1 U4550 (.I(N9064), .ZN(n17422));
    INVX1 U4551 (.I(N9065), .ZN(n17423));
    INVX1 U4552 (.I(N9066), .ZN(n17424));
    INVX1 U4553 (.I(N9067), .ZN(N17425));
    INVX1 U4554 (.I(N9068), .ZN(n17426));
    INVX1 U4555 (.I(N9069), .ZN(n17427));
    INVX1 U4556 (.I(N9070), .ZN(N17428));
    INVX1 U4557 (.I(N9071), .ZN(n17429));
    INVX1 U4558 (.I(N9072), .ZN(n17430));
    INVX1 U4559 (.I(N9073), .ZN(N17431));
    INVX1 U4560 (.I(N9074), .ZN(n17432));
    INVX1 U4561 (.I(N9075), .ZN(n17433));
    INVX1 U4562 (.I(N9076), .ZN(n17434));
    INVX1 U4563 (.I(N9077), .ZN(n17435));
    INVX1 U4564 (.I(N9078), .ZN(n17436));
    INVX1 U4565 (.I(N9079), .ZN(n17437));
    INVX1 U4566 (.I(N9080), .ZN(n17438));
    INVX1 U4567 (.I(N9081), .ZN(n17439));
    INVX1 U4568 (.I(N9082), .ZN(n17440));
    INVX1 U4569 (.I(N9083), .ZN(n17441));
    INVX1 U4570 (.I(N9084), .ZN(n17442));
    INVX1 U4571 (.I(N9085), .ZN(n17443));
    INVX1 U4572 (.I(N9086), .ZN(N17444));
    INVX1 U4573 (.I(N9087), .ZN(N17445));
    INVX1 U4574 (.I(N9088), .ZN(N17446));
    INVX1 U4575 (.I(N9089), .ZN(n17447));
    INVX1 U4576 (.I(N9090), .ZN(n17448));
    INVX1 U4577 (.I(N9091), .ZN(n17449));
    INVX1 U4578 (.I(N9092), .ZN(n17450));
    INVX1 U4579 (.I(N9093), .ZN(N17451));
    INVX1 U4580 (.I(N9094), .ZN(n17452));
    INVX1 U4581 (.I(N9095), .ZN(n17453));
    INVX1 U4582 (.I(N9096), .ZN(n17454));
    INVX1 U4583 (.I(N9097), .ZN(n17455));
    INVX1 U4584 (.I(N9098), .ZN(n17456));
    INVX1 U4585 (.I(N9099), .ZN(n17457));
    INVX1 U4586 (.I(N9100), .ZN(n17458));
    INVX1 U4587 (.I(N9101), .ZN(N17459));
    INVX1 U4588 (.I(N9102), .ZN(N17460));
    INVX1 U4589 (.I(N9103), .ZN(n17461));
    INVX1 U4590 (.I(N9104), .ZN(n17462));
    INVX1 U4591 (.I(N9105), .ZN(n17463));
    INVX1 U4592 (.I(N9106), .ZN(N17464));
    INVX1 U4593 (.I(N9107), .ZN(n17465));
    INVX1 U4594 (.I(N9108), .ZN(n17466));
    INVX1 U4595 (.I(N9109), .ZN(n17467));
    INVX1 U4596 (.I(N9110), .ZN(n17468));
    INVX1 U4597 (.I(N9111), .ZN(n17469));
    INVX1 U4598 (.I(N9112), .ZN(n17470));
    INVX1 U4599 (.I(N9113), .ZN(n17471));
    INVX1 U4600 (.I(N9114), .ZN(n17472));
    INVX1 U4601 (.I(N9115), .ZN(n17473));
    INVX1 U4602 (.I(N9116), .ZN(n17474));
    INVX1 U4603 (.I(N9117), .ZN(n17475));
    INVX1 U4604 (.I(N9118), .ZN(n17476));
    INVX1 U4605 (.I(N9119), .ZN(n17477));
    INVX1 U4606 (.I(N9120), .ZN(n17478));
    INVX1 U4607 (.I(N9121), .ZN(n17479));
    INVX1 U4608 (.I(N9122), .ZN(N17480));
    INVX1 U4609 (.I(N9123), .ZN(n17481));
    INVX1 U4610 (.I(N9124), .ZN(N17482));
    INVX1 U4611 (.I(N9125), .ZN(n17483));
    INVX1 U4612 (.I(N9126), .ZN(n17484));
    INVX1 U4613 (.I(N9127), .ZN(n17485));
    INVX1 U4614 (.I(N9128), .ZN(n17486));
    INVX1 U4615 (.I(N9129), .ZN(n17487));
    INVX1 U4616 (.I(N9130), .ZN(n17488));
    INVX1 U4617 (.I(N9131), .ZN(n17489));
    INVX1 U4618 (.I(N9132), .ZN(n17490));
    INVX1 U4619 (.I(N9133), .ZN(n17491));
    INVX1 U4620 (.I(N9134), .ZN(n17492));
    INVX1 U4621 (.I(N9135), .ZN(n17493));
    INVX1 U4622 (.I(N9136), .ZN(N17494));
    INVX1 U4623 (.I(N9137), .ZN(N17495));
    INVX1 U4624 (.I(N9138), .ZN(n17496));
    INVX1 U4625 (.I(N9139), .ZN(n17497));
    INVX1 U4626 (.I(N9140), .ZN(n17498));
    INVX1 U4627 (.I(N9141), .ZN(n17499));
    INVX1 U4628 (.I(N9142), .ZN(n17500));
    INVX1 U4629 (.I(N9143), .ZN(n17501));
    INVX1 U4630 (.I(N9144), .ZN(n17502));
    INVX1 U4631 (.I(N9145), .ZN(n17503));
    INVX1 U4632 (.I(N9146), .ZN(n17504));
    INVX1 U4633 (.I(N9147), .ZN(n17505));
    INVX1 U4634 (.I(N9148), .ZN(n17506));
    INVX1 U4635 (.I(N9149), .ZN(n17507));
    INVX1 U4636 (.I(N9150), .ZN(n17508));
    INVX1 U4637 (.I(N9151), .ZN(n17509));
    INVX1 U4638 (.I(N9152), .ZN(n17510));
    INVX1 U4639 (.I(N9153), .ZN(n17511));
    INVX1 U4640 (.I(N9154), .ZN(N17512));
    INVX1 U4641 (.I(N9155), .ZN(n17513));
    INVX1 U4642 (.I(N9156), .ZN(n17514));
    INVX1 U4643 (.I(N9157), .ZN(n17515));
    INVX1 U4644 (.I(N9158), .ZN(n17516));
    INVX1 U4645 (.I(N9159), .ZN(n17517));
    INVX1 U4646 (.I(N9160), .ZN(n17518));
    INVX1 U4647 (.I(N9161), .ZN(n17519));
    INVX1 U4648 (.I(N9162), .ZN(n17520));
    INVX1 U4649 (.I(N9163), .ZN(N17521));
    INVX1 U4650 (.I(N9164), .ZN(n17522));
    INVX1 U4651 (.I(N9165), .ZN(N17523));
    INVX1 U4652 (.I(N9166), .ZN(n17524));
    INVX1 U4653 (.I(N9167), .ZN(n17525));
    INVX1 U4654 (.I(N9168), .ZN(N17526));
    INVX1 U4655 (.I(N9169), .ZN(n17527));
    INVX1 U4656 (.I(N9170), .ZN(n17528));
    INVX1 U4657 (.I(N9171), .ZN(N17529));
    INVX1 U4658 (.I(N9172), .ZN(n17530));
    INVX1 U4659 (.I(N9173), .ZN(n17531));
    INVX1 U4660 (.I(N9174), .ZN(n17532));
    INVX1 U4661 (.I(N9175), .ZN(n17533));
    INVX1 U4662 (.I(N9176), .ZN(n17534));
    INVX1 U4663 (.I(N9177), .ZN(n17535));
    INVX1 U4664 (.I(N9178), .ZN(N17536));
    INVX1 U4665 (.I(N9179), .ZN(N17537));
    INVX1 U4666 (.I(N9180), .ZN(n17538));
    INVX1 U4667 (.I(N9181), .ZN(n17539));
    INVX1 U4668 (.I(N9182), .ZN(n17540));
    INVX1 U4669 (.I(N9183), .ZN(n17541));
    INVX1 U4670 (.I(N9184), .ZN(N17542));
    INVX1 U4671 (.I(N9185), .ZN(n17543));
    INVX1 U4672 (.I(N9186), .ZN(N17544));
    INVX1 U4673 (.I(N9187), .ZN(n17545));
    INVX1 U4674 (.I(N9188), .ZN(n17546));
    INVX1 U4675 (.I(N9189), .ZN(n17547));
    INVX1 U4676 (.I(N9190), .ZN(N17548));
    INVX1 U4677 (.I(N9191), .ZN(n17549));
    INVX1 U4678 (.I(N9192), .ZN(N17550));
    INVX1 U4679 (.I(N9193), .ZN(n17551));
    INVX1 U4680 (.I(N9194), .ZN(n17552));
    INVX1 U4681 (.I(N9195), .ZN(n17553));
    INVX1 U4682 (.I(N9196), .ZN(n17554));
    INVX1 U4683 (.I(N9197), .ZN(N17555));
    INVX1 U4684 (.I(N9198), .ZN(n17556));
    INVX1 U4685 (.I(N9199), .ZN(n17557));
    INVX1 U4686 (.I(N9200), .ZN(n17558));
    INVX1 U4687 (.I(N9201), .ZN(n17559));
    INVX1 U4688 (.I(N9202), .ZN(n17560));
    INVX1 U4689 (.I(N9203), .ZN(n17561));
    INVX1 U4690 (.I(N9204), .ZN(n17562));
    INVX1 U4691 (.I(N9205), .ZN(n17563));
    INVX1 U4692 (.I(N9206), .ZN(n17564));
    INVX1 U4693 (.I(N9207), .ZN(n17565));
    INVX1 U4694 (.I(N9208), .ZN(n17566));
    INVX1 U4695 (.I(N9209), .ZN(n17567));
    INVX1 U4696 (.I(N9210), .ZN(n17568));
    INVX1 U4697 (.I(N9211), .ZN(n17569));
    INVX1 U4698 (.I(N9212), .ZN(n17570));
    INVX1 U4699 (.I(N9213), .ZN(N17571));
    INVX1 U4700 (.I(N9214), .ZN(n17572));
    INVX1 U4701 (.I(N9215), .ZN(n17573));
    INVX1 U4702 (.I(N9216), .ZN(n17574));
    INVX1 U4703 (.I(N9217), .ZN(n17575));
    INVX1 U4704 (.I(N9218), .ZN(n17576));
    INVX1 U4705 (.I(N9219), .ZN(n17577));
    INVX1 U4706 (.I(N9220), .ZN(N17578));
    INVX1 U4707 (.I(N9221), .ZN(N17579));
    INVX1 U4708 (.I(N9222), .ZN(n17580));
    INVX1 U4709 (.I(N9223), .ZN(n17581));
    INVX1 U4710 (.I(N9224), .ZN(N17582));
    INVX1 U4711 (.I(N9225), .ZN(n17583));
    INVX1 U4712 (.I(N9226), .ZN(n17584));
    INVX1 U4713 (.I(N9227), .ZN(n17585));
    INVX1 U4714 (.I(N9228), .ZN(N17586));
    INVX1 U4715 (.I(N9229), .ZN(n17587));
    INVX1 U4716 (.I(N9230), .ZN(n17588));
    INVX1 U4717 (.I(N9231), .ZN(n17589));
    INVX1 U4718 (.I(N9232), .ZN(N17590));
    INVX1 U4719 (.I(N9233), .ZN(N17591));
    INVX1 U4720 (.I(N9234), .ZN(n17592));
    INVX1 U4721 (.I(N9235), .ZN(N17593));
    INVX1 U4722 (.I(N9236), .ZN(n17594));
    INVX1 U4723 (.I(N9237), .ZN(n17595));
    INVX1 U4724 (.I(N9238), .ZN(n17596));
    INVX1 U4725 (.I(N9239), .ZN(n17597));
    INVX1 U4726 (.I(N9240), .ZN(n17598));
    INVX1 U4727 (.I(N9241), .ZN(n17599));
    INVX1 U4728 (.I(N9242), .ZN(n17600));
    INVX1 U4729 (.I(N9243), .ZN(N17601));
    INVX1 U4730 (.I(N9244), .ZN(n17602));
    INVX1 U4731 (.I(N9245), .ZN(n17603));
    INVX1 U4732 (.I(N9246), .ZN(N17604));
    INVX1 U4733 (.I(N9247), .ZN(n17605));
    INVX1 U4734 (.I(N9248), .ZN(n17606));
    INVX1 U4735 (.I(N9249), .ZN(n17607));
    INVX1 U4736 (.I(N9250), .ZN(n17608));
    INVX1 U4737 (.I(N9251), .ZN(N17609));
    INVX1 U4738 (.I(N9252), .ZN(n17610));
    INVX1 U4739 (.I(N9253), .ZN(n17611));
    INVX1 U4740 (.I(N9254), .ZN(N17612));
    INVX1 U4741 (.I(N9255), .ZN(n17613));
    INVX1 U4742 (.I(N9256), .ZN(N17614));
    INVX1 U4743 (.I(N9257), .ZN(n17615));
    INVX1 U4744 (.I(N9258), .ZN(n17616));
    INVX1 U4745 (.I(N9259), .ZN(n17617));
    INVX1 U4746 (.I(N9260), .ZN(n17618));
    INVX1 U4747 (.I(N9261), .ZN(N17619));
    INVX1 U4748 (.I(N9262), .ZN(n17620));
    INVX1 U4749 (.I(N9263), .ZN(n17621));
    INVX1 U4750 (.I(N9264), .ZN(n17622));
    INVX1 U4751 (.I(N9265), .ZN(n17623));
    INVX1 U4752 (.I(N9266), .ZN(n17624));
    INVX1 U4753 (.I(N9267), .ZN(n17625));
    INVX1 U4754 (.I(N9268), .ZN(n17626));
    INVX1 U4755 (.I(N9269), .ZN(n17627));
    INVX1 U4756 (.I(N9270), .ZN(n17628));
    INVX1 U4757 (.I(N9271), .ZN(n17629));
    INVX1 U4758 (.I(N9272), .ZN(n17630));
    INVX1 U4759 (.I(N9273), .ZN(n17631));
    INVX1 U4760 (.I(N9274), .ZN(n17632));
    INVX1 U4761 (.I(N9275), .ZN(N17633));
    INVX1 U4762 (.I(N9276), .ZN(n17634));
    INVX1 U4763 (.I(N9277), .ZN(n17635));
    INVX1 U4764 (.I(N9278), .ZN(n17636));
    INVX1 U4765 (.I(N9279), .ZN(n17637));
    INVX1 U4766 (.I(N9280), .ZN(n17638));
    INVX1 U4767 (.I(N9281), .ZN(n17639));
    INVX1 U4768 (.I(N9282), .ZN(n17640));
    INVX1 U4769 (.I(N9283), .ZN(n17641));
    INVX1 U4770 (.I(N9284), .ZN(N17642));
    INVX1 U4771 (.I(N9285), .ZN(n17643));
    INVX1 U4772 (.I(N9286), .ZN(n17644));
    INVX1 U4773 (.I(N9287), .ZN(n17645));
    INVX1 U4774 (.I(N9288), .ZN(n17646));
    INVX1 U4775 (.I(N9289), .ZN(n17647));
    INVX1 U4776 (.I(N9290), .ZN(n17648));
    INVX1 U4777 (.I(N9291), .ZN(N17649));
    INVX1 U4778 (.I(N9292), .ZN(N17650));
    INVX1 U4779 (.I(N9293), .ZN(n17651));
    INVX1 U4780 (.I(N9294), .ZN(n17652));
    INVX1 U4781 (.I(N9295), .ZN(n17653));
    INVX1 U4782 (.I(N9296), .ZN(n17654));
    INVX1 U4783 (.I(N9297), .ZN(n17655));
    INVX1 U4784 (.I(N9298), .ZN(n17656));
    INVX1 U4785 (.I(N9299), .ZN(n17657));
    INVX1 U4786 (.I(N9300), .ZN(n17658));
    INVX1 U4787 (.I(N9301), .ZN(n17659));
    INVX1 U4788 (.I(N9302), .ZN(n17660));
    INVX1 U4789 (.I(N9303), .ZN(n17661));
    INVX1 U4790 (.I(N9304), .ZN(N17662));
    INVX1 U4791 (.I(N9305), .ZN(n17663));
    INVX1 U4792 (.I(N9306), .ZN(n17664));
    INVX1 U4793 (.I(N9307), .ZN(N17665));
    INVX1 U4794 (.I(N9308), .ZN(n17666));
    INVX1 U4795 (.I(N9309), .ZN(n17667));
    INVX1 U4796 (.I(N9310), .ZN(n17668));
    INVX1 U4797 (.I(N9311), .ZN(n17669));
    INVX1 U4798 (.I(N9312), .ZN(n17670));
    INVX1 U4799 (.I(N9313), .ZN(n17671));
    INVX1 U4800 (.I(N9314), .ZN(n17672));
    INVX1 U4801 (.I(N9315), .ZN(N17673));
    INVX1 U4802 (.I(N9316), .ZN(N17674));
    INVX1 U4803 (.I(N9317), .ZN(N17675));
    INVX1 U4804 (.I(N9318), .ZN(n17676));
    INVX1 U4805 (.I(N9319), .ZN(n17677));
    INVX1 U4806 (.I(N9320), .ZN(n17678));
    INVX1 U4807 (.I(N9321), .ZN(n17679));
    INVX1 U4808 (.I(N9322), .ZN(n17680));
    INVX1 U4809 (.I(N9323), .ZN(n17681));
    INVX1 U4810 (.I(N9324), .ZN(n17682));
    INVX1 U4811 (.I(N9325), .ZN(n17683));
    INVX1 U4812 (.I(N9326), .ZN(n17684));
    INVX1 U4813 (.I(N9327), .ZN(N17685));
    INVX1 U4814 (.I(N9328), .ZN(N17686));
    INVX1 U4815 (.I(N9329), .ZN(n17687));
    INVX1 U4816 (.I(N9330), .ZN(n17688));
    INVX1 U4817 (.I(N9331), .ZN(n17689));
    INVX1 U4818 (.I(N9332), .ZN(n17690));
    INVX1 U4819 (.I(N9333), .ZN(n17691));
    INVX1 U4820 (.I(N9334), .ZN(n17692));
    INVX1 U4821 (.I(N9335), .ZN(n17693));
    INVX1 U4822 (.I(N9336), .ZN(n17694));
    INVX1 U4823 (.I(N9337), .ZN(n17695));
    INVX1 U4824 (.I(N9338), .ZN(n17696));
    INVX1 U4825 (.I(N9339), .ZN(n17697));
    INVX1 U4826 (.I(N9340), .ZN(n17698));
    INVX1 U4827 (.I(N9341), .ZN(n17699));
    INVX1 U4828 (.I(N9342), .ZN(n17700));
    INVX1 U4829 (.I(N9343), .ZN(N17701));
    INVX1 U4830 (.I(N9344), .ZN(n17702));
    INVX1 U4831 (.I(N9345), .ZN(n17703));
    INVX1 U4832 (.I(N9346), .ZN(n17704));
    INVX1 U4833 (.I(N9347), .ZN(n17705));
    INVX1 U4834 (.I(N9348), .ZN(n17706));
    INVX1 U4835 (.I(N9349), .ZN(N17707));
    INVX1 U4836 (.I(N9350), .ZN(n17708));
    INVX1 U4837 (.I(N9351), .ZN(N17709));
    INVX1 U4838 (.I(N9352), .ZN(n17710));
    INVX1 U4839 (.I(N9353), .ZN(N17711));
    INVX1 U4840 (.I(N9354), .ZN(n17712));
    INVX1 U4841 (.I(N9355), .ZN(n17713));
    INVX1 U4842 (.I(N9356), .ZN(n17714));
    INVX1 U4843 (.I(N9357), .ZN(n17715));
    INVX1 U4844 (.I(N9358), .ZN(n17716));
    INVX1 U4845 (.I(N9359), .ZN(n17717));
    INVX1 U4846 (.I(N9360), .ZN(n17718));
    INVX1 U4847 (.I(N9361), .ZN(N17719));
    INVX1 U4848 (.I(N9362), .ZN(n17720));
    INVX1 U4849 (.I(N9363), .ZN(n17721));
    INVX1 U4850 (.I(N9364), .ZN(n17722));
    INVX1 U4851 (.I(N9365), .ZN(N17723));
    INVX1 U4852 (.I(N9366), .ZN(n17724));
    INVX1 U4853 (.I(N9367), .ZN(n17725));
    INVX1 U4854 (.I(N9368), .ZN(n17726));
    INVX1 U4855 (.I(N9369), .ZN(N17727));
    INVX1 U4856 (.I(N9370), .ZN(N17728));
    INVX1 U4857 (.I(N9371), .ZN(n17729));
    INVX1 U4858 (.I(N9372), .ZN(n17730));
    INVX1 U4859 (.I(N9373), .ZN(n17731));
    INVX1 U4860 (.I(N9374), .ZN(n17732));
    INVX1 U4861 (.I(N9375), .ZN(n17733));
    INVX1 U4862 (.I(N9376), .ZN(n17734));
    INVX1 U4863 (.I(N9377), .ZN(N17735));
    INVX1 U4864 (.I(N9378), .ZN(n17736));
    INVX1 U4865 (.I(N9379), .ZN(n17737));
    INVX1 U4866 (.I(N9380), .ZN(n17738));
    INVX1 U4867 (.I(N9381), .ZN(n17739));
    INVX1 U4868 (.I(N9382), .ZN(n17740));
    INVX1 U4869 (.I(N9383), .ZN(n17741));
    INVX1 U4870 (.I(N9384), .ZN(n17742));
    INVX1 U4871 (.I(N9385), .ZN(n17743));
    INVX1 U4872 (.I(N9386), .ZN(n17744));
    INVX1 U4873 (.I(N9387), .ZN(N17745));
    INVX1 U4874 (.I(N9388), .ZN(n17746));
    INVX1 U4875 (.I(N9389), .ZN(n17747));
    INVX1 U4876 (.I(N9390), .ZN(n17748));
    INVX1 U4877 (.I(N9391), .ZN(N17749));
    INVX1 U4878 (.I(N9392), .ZN(n17750));
    INVX1 U4879 (.I(N9393), .ZN(n17751));
    INVX1 U4880 (.I(N9394), .ZN(n17752));
    INVX1 U4881 (.I(N9395), .ZN(N17753));
    INVX1 U4882 (.I(N9396), .ZN(n17754));
    INVX1 U4883 (.I(N9397), .ZN(n17755));
    INVX1 U4884 (.I(N9398), .ZN(n17756));
    INVX1 U4885 (.I(N9399), .ZN(n17757));
    INVX1 U4886 (.I(N9400), .ZN(n17758));
    INVX1 U4887 (.I(N9401), .ZN(n17759));
    INVX1 U4888 (.I(N9402), .ZN(n17760));
    INVX1 U4889 (.I(N9403), .ZN(n17761));
    INVX1 U4890 (.I(N9404), .ZN(n17762));
    INVX1 U4891 (.I(N9405), .ZN(n17763));
    INVX1 U4892 (.I(N9406), .ZN(n17764));
    INVX1 U4893 (.I(N9407), .ZN(n17765));
    INVX1 U4894 (.I(N9408), .ZN(N17766));
    INVX1 U4895 (.I(N9409), .ZN(n17767));
    INVX1 U4896 (.I(N9410), .ZN(n17768));
    INVX1 U4897 (.I(N9411), .ZN(n17769));
    INVX1 U4898 (.I(N9412), .ZN(N17770));
    INVX1 U4899 (.I(N9413), .ZN(n17771));
    INVX1 U4900 (.I(N9414), .ZN(n17772));
    INVX1 U4901 (.I(N9415), .ZN(n17773));
    INVX1 U4902 (.I(N9416), .ZN(n17774));
    INVX1 U4903 (.I(N9417), .ZN(n17775));
    INVX1 U4904 (.I(N9418), .ZN(n17776));
    INVX1 U4905 (.I(N9419), .ZN(n17777));
    INVX1 U4906 (.I(N9420), .ZN(n17778));
    INVX1 U4907 (.I(N9421), .ZN(n17779));
    INVX1 U4908 (.I(N9422), .ZN(n17780));
    INVX1 U4909 (.I(N9423), .ZN(n17781));
    INVX1 U4910 (.I(N9424), .ZN(n17782));
    INVX1 U4911 (.I(N9425), .ZN(n17783));
    INVX1 U4912 (.I(N9426), .ZN(n17784));
    INVX1 U4913 (.I(N9427), .ZN(n17785));
    INVX1 U4914 (.I(N9428), .ZN(n17786));
    INVX1 U4915 (.I(N9429), .ZN(n17787));
    INVX1 U4916 (.I(N9430), .ZN(n17788));
    INVX1 U4917 (.I(N9431), .ZN(n17789));
    INVX1 U4918 (.I(N9432), .ZN(n17790));
    INVX1 U4919 (.I(N9433), .ZN(n17791));
    INVX1 U4920 (.I(N9434), .ZN(n17792));
    INVX1 U4921 (.I(N9435), .ZN(n17793));
    INVX1 U4922 (.I(N9436), .ZN(N17794));
    INVX1 U4923 (.I(N9437), .ZN(n17795));
    INVX1 U4924 (.I(N9438), .ZN(n17796));
    INVX1 U4925 (.I(N9439), .ZN(n17797));
    INVX1 U4926 (.I(N9440), .ZN(n17798));
    INVX1 U4927 (.I(N9441), .ZN(n17799));
    INVX1 U4928 (.I(N9442), .ZN(N17800));
    INVX1 U4929 (.I(N9443), .ZN(n17801));
    INVX1 U4930 (.I(N9444), .ZN(n17802));
    INVX1 U4931 (.I(N9445), .ZN(n17803));
    INVX1 U4932 (.I(N9446), .ZN(N17804));
    INVX1 U4933 (.I(N9447), .ZN(n17805));
    INVX1 U4934 (.I(N9448), .ZN(N17806));
    INVX1 U4935 (.I(N9449), .ZN(n17807));
    INVX1 U4936 (.I(N9450), .ZN(n17808));
    INVX1 U4937 (.I(N9451), .ZN(n17809));
    INVX1 U4938 (.I(N9452), .ZN(n17810));
    INVX1 U4939 (.I(N9453), .ZN(n17811));
    INVX1 U4940 (.I(N9454), .ZN(n17812));
    INVX1 U4941 (.I(N9455), .ZN(n17813));
    INVX1 U4942 (.I(N9456), .ZN(n17814));
    INVX1 U4943 (.I(N9457), .ZN(n17815));
    INVX1 U4944 (.I(N9458), .ZN(n17816));
    INVX1 U4945 (.I(N9459), .ZN(n17817));
    INVX1 U4946 (.I(N9460), .ZN(n17818));
    INVX1 U4947 (.I(N9461), .ZN(n17819));
    INVX1 U4948 (.I(N9462), .ZN(n17820));
    INVX1 U4949 (.I(N9463), .ZN(n17821));
    INVX1 U4950 (.I(N9464), .ZN(n17822));
    INVX1 U4951 (.I(N9465), .ZN(n17823));
    INVX1 U4952 (.I(N9466), .ZN(n17824));
    INVX1 U4953 (.I(N9467), .ZN(n17825));
    INVX1 U4954 (.I(N9468), .ZN(n17826));
    INVX1 U4955 (.I(N9469), .ZN(n17827));
    INVX1 U4956 (.I(N9470), .ZN(n17828));
    INVX1 U4957 (.I(N9471), .ZN(n17829));
    INVX1 U4958 (.I(N9472), .ZN(n17830));
    INVX1 U4959 (.I(N9473), .ZN(n17831));
    INVX1 U4960 (.I(N9474), .ZN(N17832));
    INVX1 U4961 (.I(N9475), .ZN(n17833));
    INVX1 U4962 (.I(N9476), .ZN(n17834));
    INVX1 U4963 (.I(N9477), .ZN(n17835));
    INVX1 U4964 (.I(N9478), .ZN(n17836));
    INVX1 U4965 (.I(N9479), .ZN(n17837));
    INVX1 U4966 (.I(N9480), .ZN(N17838));
    INVX1 U4967 (.I(N9481), .ZN(n17839));
    INVX1 U4968 (.I(N9482), .ZN(n17840));
    INVX1 U4969 (.I(N9483), .ZN(n17841));
    INVX1 U4970 (.I(N9484), .ZN(n17842));
    INVX1 U4971 (.I(N9485), .ZN(N17843));
    INVX1 U4972 (.I(N9486), .ZN(n17844));
    INVX1 U4973 (.I(N9487), .ZN(n17845));
    INVX1 U4974 (.I(N9488), .ZN(n17846));
    INVX1 U4975 (.I(N9489), .ZN(N17847));
    INVX1 U4976 (.I(N9490), .ZN(n17848));
    INVX1 U4977 (.I(N9491), .ZN(n17849));
    INVX1 U4978 (.I(N9492), .ZN(n17850));
    INVX1 U4979 (.I(N9493), .ZN(n17851));
    INVX1 U4980 (.I(N9494), .ZN(N17852));
    INVX1 U4981 (.I(N9495), .ZN(n17853));
    INVX1 U4982 (.I(N9496), .ZN(n17854));
    INVX1 U4983 (.I(N9497), .ZN(n17855));
    INVX1 U4984 (.I(N9498), .ZN(n17856));
    INVX1 U4985 (.I(N9499), .ZN(n17857));
    INVX1 U4986 (.I(N9500), .ZN(N17858));
    INVX1 U4987 (.I(N9501), .ZN(n17859));
    INVX1 U4988 (.I(N9502), .ZN(n17860));
    INVX1 U4989 (.I(N9503), .ZN(n17861));
    INVX1 U4990 (.I(N9504), .ZN(n17862));
    INVX1 U4991 (.I(N9505), .ZN(n17863));
    INVX1 U4992 (.I(N9506), .ZN(n17864));
    INVX1 U4993 (.I(N9507), .ZN(n17865));
    INVX1 U4994 (.I(N9508), .ZN(n17866));
    INVX1 U4995 (.I(N9509), .ZN(n17867));
    INVX1 U4996 (.I(N9510), .ZN(n17868));
    INVX1 U4997 (.I(N9511), .ZN(n17869));
    INVX1 U4998 (.I(N9512), .ZN(n17870));
    INVX1 U4999 (.I(N9513), .ZN(n17871));
    INVX1 U5000 (.I(N9514), .ZN(n17872));
    INVX1 U5001 (.I(N9515), .ZN(n17873));
    INVX1 U5002 (.I(N9516), .ZN(n17874));
    INVX1 U5003 (.I(N9517), .ZN(n17875));
    INVX1 U5004 (.I(N9518), .ZN(n17876));
    INVX1 U5005 (.I(N9519), .ZN(n17877));
    INVX1 U5006 (.I(N9520), .ZN(n17878));
    INVX1 U5007 (.I(N9521), .ZN(n17879));
    INVX1 U5008 (.I(N9522), .ZN(n17880));
    INVX1 U5009 (.I(N9523), .ZN(n17881));
    INVX1 U5010 (.I(N9524), .ZN(n17882));
    INVX1 U5011 (.I(N9525), .ZN(n17883));
    INVX1 U5012 (.I(N9526), .ZN(n17884));
    INVX1 U5013 (.I(N9527), .ZN(N17885));
    INVX1 U5014 (.I(N9528), .ZN(n17886));
    INVX1 U5015 (.I(N9529), .ZN(n17887));
    INVX1 U5016 (.I(N9530), .ZN(N17888));
    INVX1 U5017 (.I(N9531), .ZN(n17889));
    INVX1 U5018 (.I(N9532), .ZN(n17890));
    INVX1 U5019 (.I(N9533), .ZN(n17891));
    INVX1 U5020 (.I(N9534), .ZN(n17892));
    INVX1 U5021 (.I(N9535), .ZN(n17893));
    INVX1 U5022 (.I(N9536), .ZN(N17894));
    INVX1 U5023 (.I(N9537), .ZN(N17895));
    INVX1 U5024 (.I(N9538), .ZN(n17896));
    INVX1 U5025 (.I(N9539), .ZN(N17897));
    INVX1 U5026 (.I(N9540), .ZN(n17898));
    INVX1 U5027 (.I(N9541), .ZN(n17899));
    INVX1 U5028 (.I(N9542), .ZN(n17900));
    INVX1 U5029 (.I(N9543), .ZN(n17901));
    INVX1 U5030 (.I(N9544), .ZN(n17902));
    INVX1 U5031 (.I(N9545), .ZN(N17903));
    INVX1 U5032 (.I(N9546), .ZN(n17904));
    INVX1 U5033 (.I(N9547), .ZN(N17905));
    INVX1 U5034 (.I(N9548), .ZN(n17906));
    INVX1 U5035 (.I(N9549), .ZN(n17907));
    INVX1 U5036 (.I(N9550), .ZN(N17908));
    INVX1 U5037 (.I(N9551), .ZN(n17909));
    INVX1 U5038 (.I(N9552), .ZN(n17910));
    INVX1 U5039 (.I(N9553), .ZN(N17911));
    INVX1 U5040 (.I(N9554), .ZN(N17912));
    INVX1 U5041 (.I(N9555), .ZN(n17913));
    INVX1 U5042 (.I(N9556), .ZN(n17914));
    INVX1 U5043 (.I(N9557), .ZN(n17915));
    INVX1 U5044 (.I(N9558), .ZN(n17916));
    INVX1 U5045 (.I(N9559), .ZN(N17917));
    INVX1 U5046 (.I(N9560), .ZN(N17918));
    INVX1 U5047 (.I(N9561), .ZN(n17919));
    INVX1 U5048 (.I(N9562), .ZN(n17920));
    INVX1 U5049 (.I(N9563), .ZN(n17921));
    INVX1 U5050 (.I(N9564), .ZN(N17922));
    INVX1 U5051 (.I(N9565), .ZN(n17923));
    INVX1 U5052 (.I(N9566), .ZN(n17924));
    INVX1 U5053 (.I(N9567), .ZN(N17925));
    INVX1 U5054 (.I(N9568), .ZN(n17926));
    INVX1 U5055 (.I(N9569), .ZN(N17927));
    INVX1 U5056 (.I(N9570), .ZN(n17928));
    INVX1 U5057 (.I(N9571), .ZN(n17929));
    INVX1 U5058 (.I(N9572), .ZN(n17930));
    INVX1 U5059 (.I(N9573), .ZN(N17931));
    INVX1 U5060 (.I(N9574), .ZN(n17932));
    INVX1 U5061 (.I(N9575), .ZN(n17933));
    INVX1 U5062 (.I(N9576), .ZN(N17934));
    INVX1 U5063 (.I(N9577), .ZN(N17935));
    INVX1 U5064 (.I(N9578), .ZN(n17936));
    INVX1 U5065 (.I(N9579), .ZN(n17937));
    INVX1 U5066 (.I(N9580), .ZN(n17938));
    INVX1 U5067 (.I(N9581), .ZN(n17939));
    INVX1 U5068 (.I(N9582), .ZN(n17940));
    INVX1 U5069 (.I(N9583), .ZN(n17941));
    INVX1 U5070 (.I(N9584), .ZN(n17942));
    INVX1 U5071 (.I(N9585), .ZN(N17943));
    INVX1 U5072 (.I(N9586), .ZN(N17944));
    INVX1 U5073 (.I(N9587), .ZN(N17945));
    INVX1 U5074 (.I(N9588), .ZN(n17946));
    INVX1 U5075 (.I(N9589), .ZN(n17947));
    INVX1 U5076 (.I(N9590), .ZN(N17948));
    INVX1 U5077 (.I(N9591), .ZN(n17949));
    INVX1 U5078 (.I(N9592), .ZN(n17950));
    INVX1 U5079 (.I(N9593), .ZN(n17951));
    INVX1 U5080 (.I(N9594), .ZN(n17952));
    INVX1 U5081 (.I(N9595), .ZN(n17953));
    INVX1 U5082 (.I(N9596), .ZN(n17954));
    INVX1 U5083 (.I(N9597), .ZN(n17955));
    INVX1 U5084 (.I(N9598), .ZN(n17956));
    INVX1 U5085 (.I(N9599), .ZN(n17957));
    INVX1 U5086 (.I(N9600), .ZN(n17958));
    INVX1 U5087 (.I(N9601), .ZN(n17959));
    INVX1 U5088 (.I(N9602), .ZN(n17960));
    INVX1 U5089 (.I(N9603), .ZN(n17961));
    INVX1 U5090 (.I(N9604), .ZN(n17962));
    INVX1 U5091 (.I(N9605), .ZN(n17963));
    INVX1 U5092 (.I(N9606), .ZN(n17964));
    INVX1 U5093 (.I(N9607), .ZN(n17965));
    INVX1 U5094 (.I(N9608), .ZN(N17966));
    INVX1 U5095 (.I(N9609), .ZN(n17967));
    INVX1 U5096 (.I(N9610), .ZN(n17968));
    INVX1 U5097 (.I(N9611), .ZN(n17969));
    INVX1 U5098 (.I(N9612), .ZN(n17970));
    INVX1 U5099 (.I(N9613), .ZN(N17971));
    INVX1 U5100 (.I(N9614), .ZN(N17972));
    INVX1 U5101 (.I(N9615), .ZN(n17973));
    INVX1 U5102 (.I(N9616), .ZN(n17974));
    INVX1 U5103 (.I(N9617), .ZN(n17975));
    INVX1 U5104 (.I(N9618), .ZN(n17976));
    INVX1 U5105 (.I(N9619), .ZN(n17977));
    INVX1 U5106 (.I(N9620), .ZN(n17978));
    INVX1 U5107 (.I(N9621), .ZN(n17979));
    INVX1 U5108 (.I(N9622), .ZN(n17980));
    INVX1 U5109 (.I(N9623), .ZN(n17981));
    INVX1 U5110 (.I(N9624), .ZN(n17982));
    INVX1 U5111 (.I(N9625), .ZN(N17983));
    INVX1 U5112 (.I(N9626), .ZN(n17984));
    INVX1 U5113 (.I(N9627), .ZN(n17985));
    INVX1 U5114 (.I(N9628), .ZN(n17986));
    INVX1 U5115 (.I(N9629), .ZN(n17987));
    INVX1 U5116 (.I(N9630), .ZN(n17988));
    INVX1 U5117 (.I(N9631), .ZN(n17989));
    INVX1 U5118 (.I(N9632), .ZN(n17990));
    INVX1 U5119 (.I(N9633), .ZN(n17991));
    INVX1 U5120 (.I(N9634), .ZN(n17992));
    INVX1 U5121 (.I(N9635), .ZN(N17993));
    INVX1 U5122 (.I(N9636), .ZN(n17994));
    INVX1 U5123 (.I(N9637), .ZN(n17995));
    INVX1 U5124 (.I(N9638), .ZN(n17996));
    INVX1 U5125 (.I(N9639), .ZN(N17997));
    INVX1 U5126 (.I(N9640), .ZN(n17998));
    INVX1 U5127 (.I(N9641), .ZN(N17999));
    INVX1 U5128 (.I(N9642), .ZN(n18000));
    INVX1 U5129 (.I(N9643), .ZN(n18001));
    INVX1 U5130 (.I(N9644), .ZN(n18002));
    INVX1 U5131 (.I(N9645), .ZN(n18003));
    INVX1 U5132 (.I(N9646), .ZN(n18004));
    INVX1 U5133 (.I(N9647), .ZN(N18005));
    INVX1 U5134 (.I(N9648), .ZN(n18006));
    INVX1 U5135 (.I(N9649), .ZN(N18007));
    INVX1 U5136 (.I(N9650), .ZN(n18008));
    INVX1 U5137 (.I(N9651), .ZN(n18009));
    INVX1 U5138 (.I(N9652), .ZN(N18010));
    INVX1 U5139 (.I(N9653), .ZN(n18011));
    INVX1 U5140 (.I(N9654), .ZN(n18012));
    INVX1 U5141 (.I(N9655), .ZN(n18013));
    INVX1 U5142 (.I(N9656), .ZN(n18014));
    INVX1 U5143 (.I(N9657), .ZN(n18015));
    INVX1 U5144 (.I(N9658), .ZN(N18016));
    INVX1 U5145 (.I(N9659), .ZN(n18017));
    INVX1 U5146 (.I(N9660), .ZN(n18018));
    INVX1 U5147 (.I(N9661), .ZN(n18019));
    INVX1 U5148 (.I(N9662), .ZN(n18020));
    INVX1 U5149 (.I(N9663), .ZN(n18021));
    INVX1 U5150 (.I(N9664), .ZN(N18022));
    INVX1 U5151 (.I(N9665), .ZN(n18023));
    INVX1 U5152 (.I(N9666), .ZN(n18024));
    INVX1 U5153 (.I(N9667), .ZN(n18025));
    INVX1 U5154 (.I(N9668), .ZN(n18026));
    INVX1 U5155 (.I(N9669), .ZN(N18027));
    INVX1 U5156 (.I(N9670), .ZN(n18028));
    INVX1 U5157 (.I(N9671), .ZN(N18029));
    INVX1 U5158 (.I(N9672), .ZN(n18030));
    INVX1 U5159 (.I(N9673), .ZN(n18031));
    INVX1 U5160 (.I(N9674), .ZN(n18032));
    INVX1 U5161 (.I(N9675), .ZN(n18033));
    INVX1 U5162 (.I(N9676), .ZN(n18034));
    INVX1 U5163 (.I(N9677), .ZN(n18035));
    INVX1 U5164 (.I(N9678), .ZN(n18036));
    INVX1 U5165 (.I(N9679), .ZN(n18037));
    INVX1 U5166 (.I(N9680), .ZN(n18038));
    INVX1 U5167 (.I(N9681), .ZN(n18039));
    INVX1 U5168 (.I(N9682), .ZN(n18040));
    INVX1 U5169 (.I(N9683), .ZN(n18041));
    INVX1 U5170 (.I(N9684), .ZN(N18042));
    INVX1 U5171 (.I(N9685), .ZN(n18043));
    INVX1 U5172 (.I(N9686), .ZN(n18044));
    INVX1 U5173 (.I(N9687), .ZN(n18045));
    INVX1 U5174 (.I(N9688), .ZN(n18046));
    INVX1 U5175 (.I(N9689), .ZN(n18047));
    INVX1 U5176 (.I(N9690), .ZN(n18048));
    INVX1 U5177 (.I(N9691), .ZN(n18049));
    INVX1 U5178 (.I(N9692), .ZN(n18050));
    INVX1 U5179 (.I(N9693), .ZN(n18051));
    INVX1 U5180 (.I(N9694), .ZN(n18052));
    INVX1 U5181 (.I(N9695), .ZN(n18053));
    INVX1 U5182 (.I(N9696), .ZN(N18054));
    INVX1 U5183 (.I(N9697), .ZN(n18055));
    INVX1 U5184 (.I(N9698), .ZN(n18056));
    INVX1 U5185 (.I(N9699), .ZN(n18057));
    INVX1 U5186 (.I(N9700), .ZN(N18058));
    INVX1 U5187 (.I(N9701), .ZN(n18059));
    INVX1 U5188 (.I(N9702), .ZN(N18060));
    INVX1 U5189 (.I(N9703), .ZN(n18061));
    INVX1 U5190 (.I(N9704), .ZN(n18062));
    INVX1 U5191 (.I(N9705), .ZN(n18063));
    INVX1 U5192 (.I(N9706), .ZN(n18064));
    INVX1 U5193 (.I(N9707), .ZN(n18065));
    INVX1 U5194 (.I(N9708), .ZN(n18066));
    INVX1 U5195 (.I(N9709), .ZN(n18067));
    INVX1 U5196 (.I(N9710), .ZN(n18068));
    INVX1 U5197 (.I(N9711), .ZN(n18069));
    INVX1 U5198 (.I(N9712), .ZN(n18070));
    INVX1 U5199 (.I(N9713), .ZN(n18071));
    INVX1 U5200 (.I(N9714), .ZN(n18072));
    INVX1 U5201 (.I(N9715), .ZN(n18073));
    INVX1 U5202 (.I(N9716), .ZN(n18074));
    INVX1 U5203 (.I(N9717), .ZN(n18075));
    INVX1 U5204 (.I(N9718), .ZN(n18076));
    INVX1 U5205 (.I(N9719), .ZN(n18077));
    INVX1 U5206 (.I(N9720), .ZN(n18078));
    INVX1 U5207 (.I(N9721), .ZN(n18079));
    INVX1 U5208 (.I(N9722), .ZN(n18080));
    INVX1 U5209 (.I(N9723), .ZN(N18081));
    INVX1 U5210 (.I(N9724), .ZN(n18082));
    INVX1 U5211 (.I(N9725), .ZN(n18083));
    INVX1 U5212 (.I(N9726), .ZN(n18084));
    INVX1 U5213 (.I(N9727), .ZN(n18085));
    INVX1 U5214 (.I(N9728), .ZN(n18086));
    INVX1 U5215 (.I(N9729), .ZN(n18087));
    INVX1 U5216 (.I(N9730), .ZN(n18088));
    INVX1 U5217 (.I(N9731), .ZN(n18089));
    INVX1 U5218 (.I(N9732), .ZN(n18090));
    INVX1 U5219 (.I(N9733), .ZN(n18091));
    INVX1 U5220 (.I(N9734), .ZN(n18092));
    INVX1 U5221 (.I(N9735), .ZN(n18093));
    INVX1 U5222 (.I(N9736), .ZN(n18094));
    INVX1 U5223 (.I(N9737), .ZN(n18095));
    INVX1 U5224 (.I(N9738), .ZN(n18096));
    INVX1 U5225 (.I(N9739), .ZN(N18097));
    INVX1 U5226 (.I(N9740), .ZN(n18098));
    INVX1 U5227 (.I(N9741), .ZN(n18099));
    INVX1 U5228 (.I(N9742), .ZN(n18100));
    INVX1 U5229 (.I(N9743), .ZN(N18101));
    INVX1 U5230 (.I(N9744), .ZN(n18102));
    INVX1 U5231 (.I(N9745), .ZN(n18103));
    INVX1 U5232 (.I(N9746), .ZN(n18104));
    INVX1 U5233 (.I(N9747), .ZN(n18105));
    INVX1 U5234 (.I(N9748), .ZN(n18106));
    INVX1 U5235 (.I(N9749), .ZN(n18107));
    INVX1 U5236 (.I(N9750), .ZN(n18108));
    INVX1 U5237 (.I(N9751), .ZN(N18109));
    INVX1 U5238 (.I(N9752), .ZN(N18110));
    INVX1 U5239 (.I(N9753), .ZN(n18111));
    INVX1 U5240 (.I(N9754), .ZN(N18112));
    INVX1 U5241 (.I(N9755), .ZN(n18113));
    INVX1 U5242 (.I(N9756), .ZN(n18114));
    INVX1 U5243 (.I(N9757), .ZN(n18115));
    INVX1 U5244 (.I(N9758), .ZN(n18116));
    INVX1 U5245 (.I(N9759), .ZN(n18117));
    INVX1 U5246 (.I(N9760), .ZN(n18118));
    INVX1 U5247 (.I(N9761), .ZN(n18119));
    INVX1 U5248 (.I(N9762), .ZN(N18120));
    INVX1 U5249 (.I(N9763), .ZN(n18121));
    INVX1 U5250 (.I(N9764), .ZN(n18122));
    INVX1 U5251 (.I(N9765), .ZN(n18123));
    INVX1 U5252 (.I(N9766), .ZN(n18124));
    INVX1 U5253 (.I(N9767), .ZN(n18125));
    INVX1 U5254 (.I(N9768), .ZN(N18126));
    INVX1 U5255 (.I(N9769), .ZN(n18127));
    INVX1 U5256 (.I(N9770), .ZN(n18128));
    INVX1 U5257 (.I(N9771), .ZN(n18129));
    INVX1 U5258 (.I(N9772), .ZN(n18130));
    INVX1 U5259 (.I(N9773), .ZN(n18131));
    INVX1 U5260 (.I(N9774), .ZN(n18132));
    INVX1 U5261 (.I(N9775), .ZN(n18133));
    INVX1 U5262 (.I(N9776), .ZN(n18134));
    INVX1 U5263 (.I(N9777), .ZN(n18135));
    INVX1 U5264 (.I(N9778), .ZN(n18136));
    INVX1 U5265 (.I(N9779), .ZN(n18137));
    INVX1 U5266 (.I(N9780), .ZN(N18138));
    INVX1 U5267 (.I(N9781), .ZN(n18139));
    INVX1 U5268 (.I(N9782), .ZN(n18140));
    INVX1 U5269 (.I(N9783), .ZN(n18141));
    INVX1 U5270 (.I(N9784), .ZN(n18142));
    INVX1 U5271 (.I(N9785), .ZN(n18143));
    INVX1 U5272 (.I(N9786), .ZN(N18144));
    INVX1 U5273 (.I(N9787), .ZN(n18145));
    INVX1 U5274 (.I(N9788), .ZN(n18146));
    INVX1 U5275 (.I(N9789), .ZN(n18147));
    INVX1 U5276 (.I(N9790), .ZN(n18148));
    INVX1 U5277 (.I(N9791), .ZN(N18149));
    INVX1 U5278 (.I(N9792), .ZN(n18150));
    INVX1 U5279 (.I(N9793), .ZN(n18151));
    INVX1 U5280 (.I(N9794), .ZN(n18152));
    INVX1 U5281 (.I(N9795), .ZN(N18153));
    INVX1 U5282 (.I(N9796), .ZN(n18154));
    INVX1 U5283 (.I(N9797), .ZN(n18155));
    INVX1 U5284 (.I(N9798), .ZN(n18156));
    INVX1 U5285 (.I(N9799), .ZN(N18157));
    INVX1 U5286 (.I(N9800), .ZN(n18158));
    INVX1 U5287 (.I(N9801), .ZN(N18159));
    INVX1 U5288 (.I(N9802), .ZN(n18160));
    INVX1 U5289 (.I(N9803), .ZN(n18161));
    INVX1 U5290 (.I(N9804), .ZN(n18162));
    INVX1 U5291 (.I(N9805), .ZN(n18163));
    INVX1 U5292 (.I(N9806), .ZN(n18164));
    INVX1 U5293 (.I(N9807), .ZN(n18165));
    INVX1 U5294 (.I(N9808), .ZN(N18166));
    INVX1 U5295 (.I(N9809), .ZN(n18167));
    INVX1 U5296 (.I(N9810), .ZN(n18168));
    INVX1 U5297 (.I(N9811), .ZN(n18169));
    INVX1 U5298 (.I(N9812), .ZN(n18170));
    INVX1 U5299 (.I(N9813), .ZN(n18171));
    INVX1 U5300 (.I(N9814), .ZN(N18172));
    INVX1 U5301 (.I(N9815), .ZN(N18173));
    INVX1 U5302 (.I(N9816), .ZN(N18174));
    INVX1 U5303 (.I(N9817), .ZN(n18175));
    INVX1 U5304 (.I(N9818), .ZN(n18176));
    INVX1 U5305 (.I(N9819), .ZN(n18177));
    INVX1 U5306 (.I(N9820), .ZN(n18178));
    INVX1 U5307 (.I(N9821), .ZN(n18179));
    INVX1 U5308 (.I(N9822), .ZN(n18180));
    INVX1 U5309 (.I(N9823), .ZN(n18181));
    INVX1 U5310 (.I(N9824), .ZN(n18182));
    INVX1 U5311 (.I(N9825), .ZN(n18183));
    INVX1 U5312 (.I(N9826), .ZN(n18184));
    INVX1 U5313 (.I(N9827), .ZN(n18185));
    INVX1 U5314 (.I(N9828), .ZN(n18186));
    INVX1 U5315 (.I(N9829), .ZN(n18187));
    INVX1 U5316 (.I(N9830), .ZN(n18188));
    INVX1 U5317 (.I(N9831), .ZN(N18189));
    INVX1 U5318 (.I(N9832), .ZN(n18190));
    INVX1 U5319 (.I(N9833), .ZN(n18191));
    INVX1 U5320 (.I(N9834), .ZN(n18192));
    INVX1 U5321 (.I(N9835), .ZN(n18193));
    INVX1 U5322 (.I(N9836), .ZN(n18194));
    INVX1 U5323 (.I(N9837), .ZN(n18195));
    INVX1 U5324 (.I(N9838), .ZN(n18196));
    INVX1 U5325 (.I(N9839), .ZN(n18197));
    INVX1 U5326 (.I(N9840), .ZN(n18198));
    INVX1 U5327 (.I(N9841), .ZN(n18199));
    INVX1 U5328 (.I(N9842), .ZN(n18200));
    INVX1 U5329 (.I(N9843), .ZN(N18201));
    INVX1 U5330 (.I(N9844), .ZN(n18202));
    INVX1 U5331 (.I(N9845), .ZN(N18203));
    INVX1 U5332 (.I(N9846), .ZN(n18204));
    INVX1 U5333 (.I(N9847), .ZN(n18205));
    INVX1 U5334 (.I(N9848), .ZN(n18206));
    INVX1 U5335 (.I(N9849), .ZN(n18207));
    INVX1 U5336 (.I(N9850), .ZN(n18208));
    INVX1 U5337 (.I(N9851), .ZN(n18209));
    INVX1 U5338 (.I(N9852), .ZN(n18210));
    INVX1 U5339 (.I(N9853), .ZN(n18211));
    INVX1 U5340 (.I(N9854), .ZN(n18212));
    INVX1 U5341 (.I(N9855), .ZN(n18213));
    INVX1 U5342 (.I(N9856), .ZN(n18214));
    INVX1 U5343 (.I(N9857), .ZN(n18215));
    INVX1 U5344 (.I(N9858), .ZN(n18216));
    INVX1 U5345 (.I(N9859), .ZN(n18217));
    INVX1 U5346 (.I(N9860), .ZN(n18218));
    INVX1 U5347 (.I(N9861), .ZN(N18219));
    INVX1 U5348 (.I(N9862), .ZN(n18220));
    INVX1 U5349 (.I(N9863), .ZN(n18221));
    INVX1 U5350 (.I(N9864), .ZN(n18222));
    INVX1 U5351 (.I(N9865), .ZN(n18223));
    INVX1 U5352 (.I(N9866), .ZN(n18224));
    INVX1 U5353 (.I(N9867), .ZN(n18225));
    INVX1 U5354 (.I(N9868), .ZN(n18226));
    INVX1 U5355 (.I(N9869), .ZN(n18227));
    INVX1 U5356 (.I(N9870), .ZN(n18228));
    INVX1 U5357 (.I(N9871), .ZN(n18229));
    INVX1 U5358 (.I(N9872), .ZN(n18230));
    INVX1 U5359 (.I(N9873), .ZN(n18231));
    INVX1 U5360 (.I(N9874), .ZN(n18232));
    INVX1 U5361 (.I(N9875), .ZN(n18233));
    INVX1 U5362 (.I(N9876), .ZN(N18234));
    INVX1 U5363 (.I(N9877), .ZN(n18235));
    INVX1 U5364 (.I(N9878), .ZN(n18236));
    INVX1 U5365 (.I(N9879), .ZN(n18237));
    INVX1 U5366 (.I(N9880), .ZN(n18238));
    INVX1 U5367 (.I(N9881), .ZN(n18239));
    INVX1 U5368 (.I(N9882), .ZN(N18240));
    INVX1 U5369 (.I(N9883), .ZN(n18241));
    INVX1 U5370 (.I(N9884), .ZN(n18242));
    INVX1 U5371 (.I(N9885), .ZN(n18243));
    INVX1 U5372 (.I(N9886), .ZN(n18244));
    INVX1 U5373 (.I(N9887), .ZN(N18245));
    INVX1 U5374 (.I(N9888), .ZN(n18246));
    INVX1 U5375 (.I(N9889), .ZN(n18247));
    INVX1 U5376 (.I(N9890), .ZN(n18248));
    INVX1 U5377 (.I(N9891), .ZN(N18249));
    INVX1 U5378 (.I(N9892), .ZN(n18250));
    INVX1 U5379 (.I(N9893), .ZN(n18251));
    INVX1 U5380 (.I(N9894), .ZN(n18252));
    INVX1 U5381 (.I(N9895), .ZN(n18253));
    INVX1 U5382 (.I(N9896), .ZN(n18254));
    INVX1 U5383 (.I(N9897), .ZN(n18255));
    INVX1 U5384 (.I(N9898), .ZN(n18256));
    INVX1 U5385 (.I(N9899), .ZN(n18257));
    INVX1 U5386 (.I(N9900), .ZN(n18258));
    INVX1 U5387 (.I(N9901), .ZN(n18259));
    INVX1 U5388 (.I(N9902), .ZN(n18260));
    INVX1 U5389 (.I(N9903), .ZN(N18261));
    INVX1 U5390 (.I(N9904), .ZN(n18262));
    INVX1 U5391 (.I(N9905), .ZN(n18263));
    INVX1 U5392 (.I(N9906), .ZN(N18264));
    INVX1 U5393 (.I(N9907), .ZN(n18265));
    INVX1 U5394 (.I(N9908), .ZN(n18266));
    INVX1 U5395 (.I(N9909), .ZN(N18267));
    INVX1 U5396 (.I(N9910), .ZN(n18268));
    INVX1 U5397 (.I(N9911), .ZN(n18269));
    INVX1 U5398 (.I(N9912), .ZN(n18270));
    INVX1 U5399 (.I(N9913), .ZN(N18271));
    INVX1 U5400 (.I(N9914), .ZN(n18272));
    INVX1 U5401 (.I(N9915), .ZN(n18273));
    INVX1 U5402 (.I(N9916), .ZN(n18274));
    INVX1 U5403 (.I(N9917), .ZN(n18275));
    INVX1 U5404 (.I(N9918), .ZN(n18276));
    INVX1 U5405 (.I(N9919), .ZN(n18277));
    INVX1 U5406 (.I(N9920), .ZN(n18278));
    INVX1 U5407 (.I(N9921), .ZN(N18279));
    INVX1 U5408 (.I(N9922), .ZN(n18280));
    INVX1 U5409 (.I(N9923), .ZN(N18281));
    INVX1 U5410 (.I(N9924), .ZN(n18282));
    INVX1 U5411 (.I(N9925), .ZN(n18283));
    INVX1 U5412 (.I(N9926), .ZN(n18284));
    INVX1 U5413 (.I(N9927), .ZN(N18285));
    INVX1 U5414 (.I(N9928), .ZN(n18286));
    INVX1 U5415 (.I(N9929), .ZN(n18287));
    INVX1 U5416 (.I(N9930), .ZN(n18288));
    INVX1 U5417 (.I(N9931), .ZN(n18289));
    INVX1 U5418 (.I(N9932), .ZN(n18290));
    INVX1 U5419 (.I(N9933), .ZN(n18291));
    INVX1 U5420 (.I(N9934), .ZN(n18292));
    INVX1 U5421 (.I(N9935), .ZN(n18293));
    INVX1 U5422 (.I(N9936), .ZN(n18294));
    INVX1 U5423 (.I(N9937), .ZN(n18295));
    INVX1 U5424 (.I(N9938), .ZN(n18296));
    INVX1 U5425 (.I(N9939), .ZN(n18297));
    INVX1 U5426 (.I(N9940), .ZN(n18298));
    INVX1 U5427 (.I(N9941), .ZN(n18299));
    INVX1 U5428 (.I(N9942), .ZN(n18300));
    INVX1 U5429 (.I(N9943), .ZN(n18301));
    INVX1 U5430 (.I(N9944), .ZN(n18302));
    INVX1 U5431 (.I(N9945), .ZN(N18303));
    INVX1 U5432 (.I(N9946), .ZN(n18304));
    INVX1 U5433 (.I(N9947), .ZN(n18305));
    INVX1 U5434 (.I(N9948), .ZN(n18306));
    INVX1 U5435 (.I(N9949), .ZN(n18307));
    INVX1 U5436 (.I(N9950), .ZN(n18308));
    INVX1 U5437 (.I(N9951), .ZN(n18309));
    INVX1 U5438 (.I(N9952), .ZN(N18310));
    INVX1 U5439 (.I(N9953), .ZN(n18311));
    INVX1 U5440 (.I(N9954), .ZN(n18312));
    INVX1 U5441 (.I(N9955), .ZN(n18313));
    INVX1 U5442 (.I(N9956), .ZN(n18314));
    INVX1 U5443 (.I(N9957), .ZN(n18315));
    INVX1 U5444 (.I(N9958), .ZN(n18316));
    INVX1 U5445 (.I(N9959), .ZN(n18317));
    INVX1 U5446 (.I(N9960), .ZN(n18318));
    INVX1 U5447 (.I(N9961), .ZN(n18319));
    INVX1 U5448 (.I(N9962), .ZN(n18320));
    INVX1 U5449 (.I(N9963), .ZN(n18321));
    INVX1 U5450 (.I(N9964), .ZN(N18322));
    INVX1 U5451 (.I(N9965), .ZN(n18323));
    INVX1 U5452 (.I(N9966), .ZN(n18324));
    INVX1 U5453 (.I(N9967), .ZN(n18325));
    INVX1 U5454 (.I(N9968), .ZN(n18326));
    INVX1 U5455 (.I(N9969), .ZN(n18327));
    INVX1 U5456 (.I(N9970), .ZN(n18328));
    INVX1 U5457 (.I(N9971), .ZN(n18329));
    INVX1 U5458 (.I(N9972), .ZN(n18330));
    INVX1 U5459 (.I(N9973), .ZN(n18331));
    INVX1 U5460 (.I(N9974), .ZN(n18332));
    INVX1 U5461 (.I(N9975), .ZN(n18333));
    INVX1 U5462 (.I(N9976), .ZN(n18334));
    INVX1 U5463 (.I(N9977), .ZN(n18335));
    INVX1 U5464 (.I(N9978), .ZN(n18336));
    INVX1 U5465 (.I(N9979), .ZN(n18337));
    INVX1 U5466 (.I(N9980), .ZN(N18338));
    INVX1 U5467 (.I(N9981), .ZN(N18339));
    INVX1 U5468 (.I(N9982), .ZN(n18340));
    INVX1 U5469 (.I(N9983), .ZN(n18341));
    INVX1 U5470 (.I(N9984), .ZN(n18342));
    INVX1 U5471 (.I(N9985), .ZN(n18343));
    INVX1 U5472 (.I(N9986), .ZN(n18344));
    INVX1 U5473 (.I(N9987), .ZN(n18345));
    INVX1 U5474 (.I(N9988), .ZN(n18346));
    INVX1 U5475 (.I(N9989), .ZN(n18347));
    INVX1 U5476 (.I(N9990), .ZN(n18348));
    INVX1 U5477 (.I(N9991), .ZN(n18349));
    INVX1 U5478 (.I(N9992), .ZN(N18350));
    INVX1 U5479 (.I(N9993), .ZN(N18351));
    INVX1 U5480 (.I(N9994), .ZN(n18352));
    INVX1 U5481 (.I(N9995), .ZN(n18353));
    INVX1 U5482 (.I(N9996), .ZN(N18354));
    INVX1 U5483 (.I(N9997), .ZN(n18355));
    INVX1 U5484 (.I(N9998), .ZN(n18356));
    INVX1 U5485 (.I(N9999), .ZN(n18357));
    INVX1 U5486 (.I(N10000), .ZN(n18358));
    INVX1 U5487 (.I(N10001), .ZN(n18359));
    INVX1 U5488 (.I(N10002), .ZN(n18360));
    INVX1 U5489 (.I(N10003), .ZN(n18361));
    INVX1 U5490 (.I(N10004), .ZN(N18362));
    INVX1 U5491 (.I(N10005), .ZN(n18363));
    INVX1 U5492 (.I(N10006), .ZN(N18364));
    INVX1 U5493 (.I(N10007), .ZN(n18365));
    INVX1 U5494 (.I(N10008), .ZN(n18366));
    INVX1 U5495 (.I(N10009), .ZN(n18367));
    INVX1 U5496 (.I(N10010), .ZN(n18368));
    INVX1 U5497 (.I(N10011), .ZN(n18369));
    INVX1 U5498 (.I(N10012), .ZN(n18370));
    INVX1 U5499 (.I(N10013), .ZN(n18371));
    INVX1 U5500 (.I(N10014), .ZN(N18372));
    INVX1 U5501 (.I(N10015), .ZN(n18373));
    INVX1 U5502 (.I(N10016), .ZN(n18374));
    INVX1 U5503 (.I(N10017), .ZN(N18375));
    INVX1 U5504 (.I(N10018), .ZN(n18376));
    INVX1 U5505 (.I(N10019), .ZN(n18377));
    INVX1 U5506 (.I(N10020), .ZN(n18378));
    INVX1 U5507 (.I(N10021), .ZN(N18379));
    INVX1 U5508 (.I(N10022), .ZN(n18380));
    INVX1 U5509 (.I(N10023), .ZN(n18381));
    INVX1 U5510 (.I(N10024), .ZN(n18382));
    INVX1 U5511 (.I(N10025), .ZN(n18383));
    INVX1 U5512 (.I(N10026), .ZN(n18384));
    INVX1 U5513 (.I(N10027), .ZN(n18385));
    INVX1 U5514 (.I(N10028), .ZN(n18386));
    INVX1 U5515 (.I(N10029), .ZN(n18387));
    INVX1 U5516 (.I(N10030), .ZN(n18388));
    INVX1 U5517 (.I(N10031), .ZN(n18389));
    INVX1 U5518 (.I(N10032), .ZN(n18390));
    INVX1 U5519 (.I(N10033), .ZN(n18391));
    INVX1 U5520 (.I(N10034), .ZN(n18392));
    INVX1 U5521 (.I(N10035), .ZN(n18393));
    INVX1 U5522 (.I(N10036), .ZN(n18394));
    INVX1 U5523 (.I(N10037), .ZN(n18395));
    INVX1 U5524 (.I(N10038), .ZN(n18396));
    INVX1 U5525 (.I(N10039), .ZN(n18397));
    INVX1 U5526 (.I(N10040), .ZN(n18398));
    INVX1 U5527 (.I(N10041), .ZN(n18399));
    INVX1 U5528 (.I(N10042), .ZN(N18400));
    INVX1 U5529 (.I(N10043), .ZN(n18401));
    INVX1 U5530 (.I(N10044), .ZN(n18402));
    INVX1 U5531 (.I(N10045), .ZN(n18403));
    INVX1 U5532 (.I(N10046), .ZN(n18404));
    INVX1 U5533 (.I(N10047), .ZN(n18405));
    INVX1 U5534 (.I(N10048), .ZN(n18406));
    INVX1 U5535 (.I(N10049), .ZN(n18407));
    INVX1 U5536 (.I(N10050), .ZN(n18408));
    INVX1 U5537 (.I(N10051), .ZN(n18409));
    INVX1 U5538 (.I(N10052), .ZN(n18410));
    INVX1 U5539 (.I(N10053), .ZN(n18411));
    INVX1 U5540 (.I(N10054), .ZN(n18412));
    INVX1 U5541 (.I(N10055), .ZN(n18413));
    INVX1 U5542 (.I(N10056), .ZN(n18414));
    INVX1 U5543 (.I(N10057), .ZN(n18415));
    INVX1 U5544 (.I(N10058), .ZN(N18416));
    INVX1 U5545 (.I(N10059), .ZN(n18417));
    INVX1 U5546 (.I(N10060), .ZN(n18418));
    INVX1 U5547 (.I(N10061), .ZN(n18419));
    INVX1 U5548 (.I(N10062), .ZN(N18420));
    INVX1 U5549 (.I(N10063), .ZN(n18421));
    INVX1 U5550 (.I(N10064), .ZN(n18422));
    INVX1 U5551 (.I(N10065), .ZN(n18423));
    INVX1 U5552 (.I(N10066), .ZN(n18424));
    INVX1 U5553 (.I(N10067), .ZN(n18425));
    INVX1 U5554 (.I(N10068), .ZN(n18426));
    INVX1 U5555 (.I(N10069), .ZN(n18427));
    INVX1 U5556 (.I(N10070), .ZN(n18428));
    INVX1 U5557 (.I(N10071), .ZN(n18429));
    INVX1 U5558 (.I(N10072), .ZN(N18430));
    INVX1 U5559 (.I(N10073), .ZN(n18431));
    INVX1 U5560 (.I(N10074), .ZN(n18432));
    INVX1 U5561 (.I(N10075), .ZN(n18433));
    INVX1 U5562 (.I(N10076), .ZN(n18434));
    INVX1 U5563 (.I(N10077), .ZN(n18435));
    INVX1 U5564 (.I(N10078), .ZN(N18436));
    INVX1 U5565 (.I(N10079), .ZN(n18437));
    INVX1 U5566 (.I(N10080), .ZN(n18438));
    INVX1 U5567 (.I(N10081), .ZN(n18439));
    INVX1 U5568 (.I(N10082), .ZN(n18440));
    INVX1 U5569 (.I(N10083), .ZN(n18441));
    INVX1 U5570 (.I(N10084), .ZN(n18442));
    INVX1 U5571 (.I(N10085), .ZN(n18443));
    INVX1 U5572 (.I(N10086), .ZN(n18444));
    INVX1 U5573 (.I(N10087), .ZN(N18445));
    INVX1 U5574 (.I(N10088), .ZN(n18446));
    INVX1 U5575 (.I(N10089), .ZN(n18447));
    INVX1 U5576 (.I(N10090), .ZN(n18448));
    INVX1 U5577 (.I(N10091), .ZN(n18449));
    INVX1 U5578 (.I(N10092), .ZN(n18450));
    INVX1 U5579 (.I(N10093), .ZN(n18451));
    INVX1 U5580 (.I(N10094), .ZN(n18452));
    INVX1 U5581 (.I(N10095), .ZN(n18453));
    INVX1 U5582 (.I(N10096), .ZN(n18454));
    INVX1 U5583 (.I(N10097), .ZN(n18455));
    INVX1 U5584 (.I(N10098), .ZN(n18456));
    INVX1 U5585 (.I(N10099), .ZN(n18457));
    INVX1 U5586 (.I(N10100), .ZN(n18458));
    INVX1 U5587 (.I(N10101), .ZN(n18459));
    INVX1 U5588 (.I(N10102), .ZN(n18460));
    INVX1 U5589 (.I(N10103), .ZN(N18461));
    INVX1 U5590 (.I(N10104), .ZN(n18462));
    INVX1 U5591 (.I(N10105), .ZN(n18463));
    INVX1 U5592 (.I(N10106), .ZN(N18464));
    INVX1 U5593 (.I(N10107), .ZN(n18465));
    INVX1 U5594 (.I(N10108), .ZN(n18466));
    INVX1 U5595 (.I(N10109), .ZN(N18467));
    INVX1 U5596 (.I(N10110), .ZN(n18468));
    INVX1 U5597 (.I(N10111), .ZN(n18469));
    INVX1 U5598 (.I(N10112), .ZN(n18470));
    INVX1 U5599 (.I(N10113), .ZN(n18471));
    INVX1 U5600 (.I(N10114), .ZN(n18472));
    INVX1 U5601 (.I(N10115), .ZN(n18473));
    INVX1 U5602 (.I(N10116), .ZN(n18474));
    INVX1 U5603 (.I(N10117), .ZN(n18475));
    INVX1 U5604 (.I(N10118), .ZN(n18476));
    INVX1 U5605 (.I(N10119), .ZN(n18477));
    INVX1 U5606 (.I(N10120), .ZN(n18478));
    INVX1 U5607 (.I(N10121), .ZN(n18479));
    INVX1 U5608 (.I(N10122), .ZN(n18480));
    INVX1 U5609 (.I(N10123), .ZN(n18481));
    INVX1 U5610 (.I(N10124), .ZN(n18482));
    INVX1 U5611 (.I(N10125), .ZN(n18483));
    INVX1 U5612 (.I(N10126), .ZN(N18484));
    INVX1 U5613 (.I(N10127), .ZN(n18485));
    INVX1 U5614 (.I(N10128), .ZN(n18486));
    INVX1 U5615 (.I(N10129), .ZN(n18487));
    INVX1 U5616 (.I(N10130), .ZN(N18488));
    INVX1 U5617 (.I(N10131), .ZN(n18489));
    INVX1 U5618 (.I(N10132), .ZN(n18490));
    INVX1 U5619 (.I(N10133), .ZN(n18491));
    INVX1 U5620 (.I(N10134), .ZN(n18492));
    INVX1 U5621 (.I(N10135), .ZN(N18493));
    INVX1 U5622 (.I(N10136), .ZN(n18494));
    INVX1 U5623 (.I(N10137), .ZN(N18495));
    INVX1 U5624 (.I(N10138), .ZN(n18496));
    INVX1 U5625 (.I(N10139), .ZN(n18497));
    INVX1 U5626 (.I(N10140), .ZN(n18498));
    INVX1 U5627 (.I(N10141), .ZN(n18499));
    INVX1 U5628 (.I(N10142), .ZN(n18500));
    INVX1 U5629 (.I(N10143), .ZN(n18501));
    INVX1 U5630 (.I(N10144), .ZN(N18502));
    INVX1 U5631 (.I(N10145), .ZN(n18503));
    INVX1 U5632 (.I(N10146), .ZN(n18504));
    INVX1 U5633 (.I(N10147), .ZN(n18505));
    INVX1 U5634 (.I(N10148), .ZN(N18506));
    INVX1 U5635 (.I(N10149), .ZN(n18507));
    INVX1 U5636 (.I(N10150), .ZN(n18508));
    INVX1 U5637 (.I(N10151), .ZN(n18509));
    INVX1 U5638 (.I(N10152), .ZN(N18510));
    INVX1 U5639 (.I(N10153), .ZN(n18511));
    INVX1 U5640 (.I(N10154), .ZN(n18512));
    INVX1 U5641 (.I(N10155), .ZN(n18513));
    INVX1 U5642 (.I(N10156), .ZN(n18514));
    INVX1 U5643 (.I(N10157), .ZN(n18515));
    INVX1 U5644 (.I(N10158), .ZN(n18516));
    INVX1 U5645 (.I(N10159), .ZN(n18517));
    INVX1 U5646 (.I(N10160), .ZN(n18518));
    INVX1 U5647 (.I(N10161), .ZN(N18519));
    INVX1 U5648 (.I(N10162), .ZN(n18520));
    INVX1 U5649 (.I(N10163), .ZN(n18521));
    INVX1 U5650 (.I(N10164), .ZN(n18522));
    INVX1 U5651 (.I(N10165), .ZN(n18523));
    INVX1 U5652 (.I(N10166), .ZN(N18524));
    INVX1 U5653 (.I(N10167), .ZN(n18525));
    INVX1 U5654 (.I(N10168), .ZN(N18526));
    INVX1 U5655 (.I(N10169), .ZN(n18527));
    INVX1 U5656 (.I(N10170), .ZN(N18528));
    INVX1 U5657 (.I(N10171), .ZN(n18529));
    INVX1 U5658 (.I(N10172), .ZN(n18530));
    INVX1 U5659 (.I(N10173), .ZN(n18531));
    INVX1 U5660 (.I(N10174), .ZN(n18532));
    INVX1 U5661 (.I(N10175), .ZN(n18533));
    INVX1 U5662 (.I(N10176), .ZN(n18534));
    INVX1 U5663 (.I(N10177), .ZN(n18535));
    INVX1 U5664 (.I(N10178), .ZN(n18536));
    INVX1 U5665 (.I(N10179), .ZN(n18537));
    INVX1 U5666 (.I(N10180), .ZN(n18538));
    INVX1 U5667 (.I(N10181), .ZN(n18539));
    INVX1 U5668 (.I(N10182), .ZN(n18540));
    INVX1 U5669 (.I(N10183), .ZN(n18541));
    INVX1 U5670 (.I(N10184), .ZN(n18542));
    INVX1 U5671 (.I(N10185), .ZN(n18543));
    INVX1 U5672 (.I(N10186), .ZN(N18544));
    INVX1 U5673 (.I(N10187), .ZN(n18545));
    INVX1 U5674 (.I(N10188), .ZN(n18546));
    INVX1 U5675 (.I(N10189), .ZN(n18547));
    INVX1 U5676 (.I(N10190), .ZN(n18548));
    INVX1 U5677 (.I(N10191), .ZN(N18549));
    INVX1 U5678 (.I(N10192), .ZN(n18550));
    INVX1 U5679 (.I(N10193), .ZN(n18551));
    INVX1 U5680 (.I(N10194), .ZN(n18552));
    INVX1 U5681 (.I(N10195), .ZN(n18553));
    INVX1 U5682 (.I(N10196), .ZN(n18554));
    INVX1 U5683 (.I(N10197), .ZN(n18555));
    INVX1 U5684 (.I(N10198), .ZN(n18556));
    INVX1 U5685 (.I(N10199), .ZN(n18557));
    INVX1 U5686 (.I(N10200), .ZN(n18558));
    INVX1 U5687 (.I(N10201), .ZN(n18559));
    INVX1 U5688 (.I(N10202), .ZN(n18560));
    INVX1 U5689 (.I(N10203), .ZN(N18561));
    INVX1 U5690 (.I(N10204), .ZN(n18562));
    INVX1 U5691 (.I(N10205), .ZN(N18563));
    INVX1 U5692 (.I(N10206), .ZN(n18564));
    INVX1 U5693 (.I(N10207), .ZN(n18565));
    INVX1 U5694 (.I(N10208), .ZN(N18566));
    INVX1 U5695 (.I(N10209), .ZN(n18567));
    INVX1 U5696 (.I(N10210), .ZN(n18568));
    INVX1 U5697 (.I(N10211), .ZN(n18569));
    INVX1 U5698 (.I(N10212), .ZN(n18570));
    INVX1 U5699 (.I(N10213), .ZN(n18571));
    INVX1 U5700 (.I(N10214), .ZN(n18572));
    INVX1 U5701 (.I(N10215), .ZN(n18573));
    INVX1 U5702 (.I(N10216), .ZN(n18574));
    INVX1 U5703 (.I(N10217), .ZN(n18575));
    INVX1 U5704 (.I(N10218), .ZN(N18576));
    INVX1 U5705 (.I(N10219), .ZN(n18577));
    INVX1 U5706 (.I(N10220), .ZN(N18578));
    INVX1 U5707 (.I(N10221), .ZN(n18579));
    INVX1 U5708 (.I(N10222), .ZN(n18580));
    INVX1 U5709 (.I(N10223), .ZN(n18581));
    INVX1 U5710 (.I(N10224), .ZN(n18582));
    INVX1 U5711 (.I(N10225), .ZN(N18583));
    INVX1 U5712 (.I(N10226), .ZN(n18584));
    INVX1 U5713 (.I(N10227), .ZN(n18585));
    INVX1 U5714 (.I(N10228), .ZN(n18586));
    INVX1 U5715 (.I(N10229), .ZN(N18587));
    INVX1 U5716 (.I(N10230), .ZN(n18588));
    INVX1 U5717 (.I(N10231), .ZN(n18589));
    INVX1 U5718 (.I(N10232), .ZN(n18590));
    INVX1 U5719 (.I(N10233), .ZN(n18591));
    INVX1 U5720 (.I(N10234), .ZN(n18592));
    INVX1 U5721 (.I(N10235), .ZN(n18593));
    INVX1 U5722 (.I(N10236), .ZN(n18594));
    INVX1 U5723 (.I(N10237), .ZN(n18595));
    INVX1 U5724 (.I(N10238), .ZN(n18596));
    INVX1 U5725 (.I(N10239), .ZN(n18597));
    INVX1 U5726 (.I(N10240), .ZN(n18598));
    INVX1 U5727 (.I(N10241), .ZN(n18599));
    INVX1 U5728 (.I(N10242), .ZN(n18600));
    INVX1 U5729 (.I(N10243), .ZN(n18601));
    INVX1 U5730 (.I(N10244), .ZN(n18602));
    INVX1 U5731 (.I(N10245), .ZN(n18603));
    INVX1 U5732 (.I(N10246), .ZN(n18604));
    INVX1 U5733 (.I(N10247), .ZN(n18605));
    INVX1 U5734 (.I(N10248), .ZN(n18606));
    INVX1 U5735 (.I(N10249), .ZN(n18607));
    INVX1 U5736 (.I(N10250), .ZN(n18608));
    INVX1 U5737 (.I(N10251), .ZN(n18609));
    INVX1 U5738 (.I(N10252), .ZN(n18610));
    INVX1 U5739 (.I(N10253), .ZN(n18611));
    INVX1 U5740 (.I(N10254), .ZN(n18612));
    INVX1 U5741 (.I(N10255), .ZN(n18613));
    INVX1 U5742 (.I(N10256), .ZN(n18614));
    INVX1 U5743 (.I(N10257), .ZN(n18615));
    INVX1 U5744 (.I(N10258), .ZN(n18616));
    INVX1 U5745 (.I(N10259), .ZN(n18617));
    INVX1 U5746 (.I(N10260), .ZN(n18618));
    INVX1 U5747 (.I(N10261), .ZN(N18619));
    INVX1 U5748 (.I(N10262), .ZN(n18620));
    INVX1 U5749 (.I(N10263), .ZN(n18621));
    INVX1 U5750 (.I(N10264), .ZN(N18622));
    INVX1 U5751 (.I(N10265), .ZN(n18623));
    INVX1 U5752 (.I(N10266), .ZN(n18624));
    INVX1 U5753 (.I(N10267), .ZN(n18625));
    INVX1 U5754 (.I(N10268), .ZN(n18626));
    INVX1 U5755 (.I(N10269), .ZN(N18627));
    INVX1 U5756 (.I(N10270), .ZN(n18628));
    INVX1 U5757 (.I(N10271), .ZN(n18629));
    INVX1 U5758 (.I(N10272), .ZN(n18630));
    INVX1 U5759 (.I(N10273), .ZN(n18631));
    INVX1 U5760 (.I(N10274), .ZN(n18632));
    INVX1 U5761 (.I(N10275), .ZN(n18633));
    INVX1 U5762 (.I(N10276), .ZN(n18634));
    INVX1 U5763 (.I(N10277), .ZN(n18635));
    INVX1 U5764 (.I(N10278), .ZN(n18636));
    INVX1 U5765 (.I(N10279), .ZN(n18637));
    INVX1 U5766 (.I(N10280), .ZN(n18638));
    INVX1 U5767 (.I(N10281), .ZN(n18639));
    INVX1 U5768 (.I(N10282), .ZN(n18640));
    INVX1 U5769 (.I(N10283), .ZN(N18641));
    INVX1 U5770 (.I(N10284), .ZN(n18642));
    INVX1 U5771 (.I(N10285), .ZN(n18643));
    INVX1 U5772 (.I(N10286), .ZN(n18644));
    INVX1 U5773 (.I(N10287), .ZN(n18645));
    INVX1 U5774 (.I(N10288), .ZN(n18646));
    INVX1 U5775 (.I(N10289), .ZN(n18647));
    INVX1 U5776 (.I(N10290), .ZN(n18648));
    INVX1 U5777 (.I(N10291), .ZN(N18649));
    INVX1 U5778 (.I(N10292), .ZN(n18650));
    INVX1 U5779 (.I(N10293), .ZN(n18651));
    INVX1 U5780 (.I(N10294), .ZN(n18652));
    INVX1 U5781 (.I(N10295), .ZN(n18653));
    INVX1 U5782 (.I(N10296), .ZN(n18654));
    INVX1 U5783 (.I(N10297), .ZN(n18655));
    INVX1 U5784 (.I(N10298), .ZN(n18656));
    INVX1 U5785 (.I(N10299), .ZN(n18657));
    INVX1 U5786 (.I(N10300), .ZN(n18658));
    INVX1 U5787 (.I(N10301), .ZN(n18659));
    INVX1 U5788 (.I(N10302), .ZN(n18660));
    INVX1 U5789 (.I(N10303), .ZN(n18661));
    INVX1 U5790 (.I(N10304), .ZN(n18662));
    INVX1 U5791 (.I(N10305), .ZN(n18663));
    INVX1 U5792 (.I(N10306), .ZN(n18664));
    INVX1 U5793 (.I(N10307), .ZN(N18665));
    INVX1 U5794 (.I(N10308), .ZN(n18666));
    INVX1 U5795 (.I(N10309), .ZN(n18667));
    INVX1 U5796 (.I(N10310), .ZN(N18668));
    INVX1 U5797 (.I(N10311), .ZN(n18669));
    INVX1 U5798 (.I(N10312), .ZN(n18670));
    INVX1 U5799 (.I(N10313), .ZN(N18671));
    INVX1 U5800 (.I(N10314), .ZN(n18672));
    INVX1 U5801 (.I(N10315), .ZN(n18673));
    INVX1 U5802 (.I(N10316), .ZN(n18674));
    INVX1 U5803 (.I(N10317), .ZN(n18675));
    INVX1 U5804 (.I(N10318), .ZN(n18676));
    INVX1 U5805 (.I(N10319), .ZN(n18677));
    INVX1 U5806 (.I(N10320), .ZN(n18678));
    INVX1 U5807 (.I(N10321), .ZN(n18679));
    INVX1 U5808 (.I(N10322), .ZN(n18680));
    INVX1 U5809 (.I(N10323), .ZN(n18681));
    INVX1 U5810 (.I(N10324), .ZN(n18682));
    INVX1 U5811 (.I(N10325), .ZN(n18683));
    INVX1 U5812 (.I(N10326), .ZN(n18684));
    INVX1 U5813 (.I(N10327), .ZN(N18685));
    INVX1 U5814 (.I(N10328), .ZN(n18686));
    INVX1 U5815 (.I(N10329), .ZN(n18687));
    INVX1 U5816 (.I(N10330), .ZN(N18688));
    INVX1 U5817 (.I(N10331), .ZN(n18689));
    INVX1 U5818 (.I(N10332), .ZN(n18690));
    INVX1 U5819 (.I(N10333), .ZN(n18691));
    INVX1 U5820 (.I(N10334), .ZN(n18692));
    INVX1 U5821 (.I(N10335), .ZN(N18693));
    INVX1 U5822 (.I(N10336), .ZN(n18694));
    INVX1 U5823 (.I(N10337), .ZN(n18695));
    INVX1 U5824 (.I(N10338), .ZN(n18696));
    INVX1 U5825 (.I(N10339), .ZN(n18697));
    INVX1 U5826 (.I(N10340), .ZN(n18698));
    INVX1 U5827 (.I(N10341), .ZN(n18699));
    INVX1 U5828 (.I(N10342), .ZN(n18700));
    INVX1 U5829 (.I(N10343), .ZN(n18701));
    INVX1 U5830 (.I(N10344), .ZN(n18702));
    INVX1 U5831 (.I(N10345), .ZN(n18703));
    INVX1 U5832 (.I(N10346), .ZN(n18704));
    INVX1 U5833 (.I(N10347), .ZN(n18705));
    INVX1 U5834 (.I(N10348), .ZN(n18706));
    INVX1 U5835 (.I(N10349), .ZN(n18707));
    INVX1 U5836 (.I(N10350), .ZN(n18708));
    INVX1 U5837 (.I(N10351), .ZN(n18709));
    INVX1 U5838 (.I(N10352), .ZN(n18710));
    INVX1 U5839 (.I(N10353), .ZN(n18711));
    INVX1 U5840 (.I(N10354), .ZN(n18712));
    INVX1 U5841 (.I(N10355), .ZN(n18713));
    INVX1 U5842 (.I(N10356), .ZN(n18714));
    INVX1 U5843 (.I(N10357), .ZN(n18715));
    INVX1 U5844 (.I(N10358), .ZN(n18716));
    INVX1 U5845 (.I(N10359), .ZN(n18717));
    INVX1 U5846 (.I(N10360), .ZN(n18718));
    INVX1 U5847 (.I(N10361), .ZN(n18719));
    INVX1 U5848 (.I(N10362), .ZN(n18720));
    INVX1 U5849 (.I(N10363), .ZN(n18721));
    INVX1 U5850 (.I(N10364), .ZN(n18722));
    INVX1 U5851 (.I(N10365), .ZN(N18723));
    INVX1 U5852 (.I(N10366), .ZN(N18724));
    INVX1 U5853 (.I(N10367), .ZN(n18725));
    INVX1 U5854 (.I(N10368), .ZN(n18726));
    INVX1 U5855 (.I(N10369), .ZN(n18727));
    INVX1 U5856 (.I(N10370), .ZN(n18728));
    INVX1 U5857 (.I(N10371), .ZN(n18729));
    INVX1 U5858 (.I(N10372), .ZN(N18730));
    INVX1 U5859 (.I(N10373), .ZN(n18731));
    INVX1 U5860 (.I(N10374), .ZN(n18732));
    INVX1 U5861 (.I(N10375), .ZN(n18733));
    INVX1 U5862 (.I(N10376), .ZN(n18734));
    INVX1 U5863 (.I(N10377), .ZN(n18735));
    INVX1 U5864 (.I(N10378), .ZN(n18736));
    INVX1 U5865 (.I(N10379), .ZN(N18737));
    INVX1 U5866 (.I(N10380), .ZN(n18738));
    INVX1 U5867 (.I(N10381), .ZN(N18739));
    INVX1 U5868 (.I(N10382), .ZN(n18740));
    INVX1 U5869 (.I(N10383), .ZN(N18741));
    INVX1 U5870 (.I(N10384), .ZN(n18742));
    INVX1 U5871 (.I(N10385), .ZN(N18743));
    INVX1 U5872 (.I(N10386), .ZN(n18744));
    INVX1 U5873 (.I(N10387), .ZN(n18745));
    INVX1 U5874 (.I(N10388), .ZN(n18746));
    INVX1 U5875 (.I(N10389), .ZN(n18747));
    INVX1 U5876 (.I(N10390), .ZN(n18748));
    INVX1 U5877 (.I(N10391), .ZN(n18749));
    INVX1 U5878 (.I(N10392), .ZN(n18750));
    INVX1 U5879 (.I(N10393), .ZN(N18751));
    INVX1 U5880 (.I(N10394), .ZN(n18752));
    INVX1 U5881 (.I(N10395), .ZN(n18753));
    INVX1 U5882 (.I(N10396), .ZN(N18754));
    INVX1 U5883 (.I(N10397), .ZN(n18755));
    INVX1 U5884 (.I(N10398), .ZN(n18756));
    INVX1 U5885 (.I(N10399), .ZN(n18757));
    INVX1 U5886 (.I(N10400), .ZN(n18758));
    INVX1 U5887 (.I(N10401), .ZN(n18759));
    INVX1 U5888 (.I(N10402), .ZN(n18760));
    INVX1 U5889 (.I(N10403), .ZN(n18761));
    INVX1 U5890 (.I(N10404), .ZN(n18762));
    INVX1 U5891 (.I(N10405), .ZN(n18763));
    INVX1 U5892 (.I(N10406), .ZN(n18764));
    INVX1 U5893 (.I(N10407), .ZN(n18765));
    INVX1 U5894 (.I(N10408), .ZN(n18766));
    INVX1 U5895 (.I(N10409), .ZN(n18767));
    INVX1 U5896 (.I(N10410), .ZN(n18768));
    INVX1 U5897 (.I(N10411), .ZN(n18769));
    INVX1 U5898 (.I(N10412), .ZN(n18770));
    INVX1 U5899 (.I(N10413), .ZN(n18771));
    INVX1 U5900 (.I(N10414), .ZN(n18772));
    INVX1 U5901 (.I(N10415), .ZN(n18773));
    INVX1 U5902 (.I(N10416), .ZN(n18774));
    INVX1 U5903 (.I(N10417), .ZN(n18775));
    INVX1 U5904 (.I(N10418), .ZN(N18776));
    INVX1 U5905 (.I(N10419), .ZN(n18777));
    INVX1 U5906 (.I(N10420), .ZN(n18778));
    INVX1 U5907 (.I(N10421), .ZN(n18779));
    INVX1 U5908 (.I(N10422), .ZN(n18780));
    INVX1 U5909 (.I(N10423), .ZN(N18781));
    INVX1 U5910 (.I(N10424), .ZN(n18782));
    INVX1 U5911 (.I(N10425), .ZN(N18783));
    INVX1 U5912 (.I(N10426), .ZN(n18784));
    INVX1 U5913 (.I(N10427), .ZN(n18785));
    INVX1 U5914 (.I(N10428), .ZN(n18786));
    INVX1 U5915 (.I(N10429), .ZN(n18787));
    INVX1 U5916 (.I(N10430), .ZN(n18788));
    INVX1 U5917 (.I(N10431), .ZN(n18789));
    INVX1 U5918 (.I(N10432), .ZN(n18790));
    INVX1 U5919 (.I(N10433), .ZN(n18791));
    INVX1 U5920 (.I(N10434), .ZN(n18792));
    INVX1 U5921 (.I(N10435), .ZN(n18793));
    INVX1 U5922 (.I(N10436), .ZN(n18794));
    INVX1 U5923 (.I(N10437), .ZN(n18795));
    INVX1 U5924 (.I(N10438), .ZN(n18796));
    INVX1 U5925 (.I(N10439), .ZN(n18797));
    INVX1 U5926 (.I(N10440), .ZN(n18798));
    INVX1 U5927 (.I(N10441), .ZN(N18799));
    INVX1 U5928 (.I(N10442), .ZN(n18800));
    INVX1 U5929 (.I(N10443), .ZN(n18801));
    INVX1 U5930 (.I(N10444), .ZN(n18802));
    INVX1 U5931 (.I(N10445), .ZN(n18803));
    INVX1 U5932 (.I(N10446), .ZN(n18804));
    INVX1 U5933 (.I(N10447), .ZN(N18805));
    INVX1 U5934 (.I(N10448), .ZN(n18806));
    INVX1 U5935 (.I(N10449), .ZN(n18807));
    INVX1 U5936 (.I(N10450), .ZN(n18808));
    INVX1 U5937 (.I(N10451), .ZN(n18809));
    INVX1 U5938 (.I(N10452), .ZN(n18810));
    INVX1 U5939 (.I(N10453), .ZN(n18811));
    INVX1 U5940 (.I(N10454), .ZN(n18812));
    INVX1 U5941 (.I(N10455), .ZN(n18813));
    INVX1 U5942 (.I(N10456), .ZN(n18814));
    INVX1 U5943 (.I(N10457), .ZN(n18815));
    INVX1 U5944 (.I(N10458), .ZN(n18816));
    INVX1 U5945 (.I(N10459), .ZN(n18817));
    INVX1 U5946 (.I(N10460), .ZN(n18818));
    INVX1 U5947 (.I(N10461), .ZN(n18819));
    INVX1 U5948 (.I(N10462), .ZN(N18820));
    INVX1 U5949 (.I(N10463), .ZN(n18821));
    INVX1 U5950 (.I(N10464), .ZN(N18822));
    INVX1 U5951 (.I(N10465), .ZN(n18823));
    INVX1 U5952 (.I(N10466), .ZN(n18824));
    INVX1 U5953 (.I(N10467), .ZN(N18825));
    INVX1 U5954 (.I(N10468), .ZN(n18826));
    INVX1 U5955 (.I(N10469), .ZN(n18827));
    INVX1 U5956 (.I(N10470), .ZN(n18828));
    INVX1 U5957 (.I(N10471), .ZN(n18829));
    INVX1 U5958 (.I(N10472), .ZN(n18830));
    INVX1 U5959 (.I(N10473), .ZN(n18831));
    INVX1 U5960 (.I(N10474), .ZN(n18832));
    INVX1 U5961 (.I(N10475), .ZN(n18833));
    INVX1 U5962 (.I(N10476), .ZN(N18834));
    INVX1 U5963 (.I(N10477), .ZN(n18835));
    INVX1 U5964 (.I(N10478), .ZN(n18836));
    INVX1 U5965 (.I(N10479), .ZN(n18837));
    INVX1 U5966 (.I(N10480), .ZN(N18838));
    INVX1 U5967 (.I(N10481), .ZN(n18839));
    INVX1 U5968 (.I(N10482), .ZN(n18840));
    INVX1 U5969 (.I(N10483), .ZN(n18841));
    INVX1 U5970 (.I(N10484), .ZN(n18842));
    INVX1 U5971 (.I(N10485), .ZN(n18843));
    INVX1 U5972 (.I(N10486), .ZN(n18844));
    INVX1 U5973 (.I(N10487), .ZN(n18845));
    INVX1 U5974 (.I(N10488), .ZN(n18846));
    INVX1 U5975 (.I(N10489), .ZN(n18847));
    INVX1 U5976 (.I(N10490), .ZN(N18848));
    INVX1 U5977 (.I(N10491), .ZN(n18849));
    INVX1 U5978 (.I(N10492), .ZN(N18850));
    INVX1 U5979 (.I(N10493), .ZN(n18851));
    INVX1 U5980 (.I(N10494), .ZN(n18852));
    INVX1 U5981 (.I(N10495), .ZN(n18853));
    INVX1 U5982 (.I(N10496), .ZN(n18854));
    INVX1 U5983 (.I(N10497), .ZN(N18855));
    INVX1 U5984 (.I(N10498), .ZN(n18856));
    INVX1 U5985 (.I(N10499), .ZN(n18857));
    INVX1 U5986 (.I(N10500), .ZN(n18858));
    INVX1 U5987 (.I(N10501), .ZN(n18859));
    INVX1 U5988 (.I(N10502), .ZN(n18860));
    INVX1 U5989 (.I(N10503), .ZN(n18861));
    INVX1 U5990 (.I(N10504), .ZN(n18862));
    INVX1 U5991 (.I(N10505), .ZN(n18863));
    INVX1 U5992 (.I(N10506), .ZN(n18864));
    INVX1 U5993 (.I(N10507), .ZN(n18865));
    INVX1 U5994 (.I(N10508), .ZN(N18866));
    INVX1 U5995 (.I(N10509), .ZN(N18867));
    INVX1 U5996 (.I(N10510), .ZN(n18868));
    INVX1 U5997 (.I(N10511), .ZN(n18869));
    INVX1 U5998 (.I(N10512), .ZN(n18870));
    INVX1 U5999 (.I(N10513), .ZN(n18871));
    INVX1 U6000 (.I(N10514), .ZN(n18872));
    INVX1 U6001 (.I(N10515), .ZN(n18873));
    INVX1 U6002 (.I(N10516), .ZN(n18874));
    INVX1 U6003 (.I(N10517), .ZN(n18875));
    INVX1 U6004 (.I(N10518), .ZN(n18876));
    INVX1 U6005 (.I(N10519), .ZN(n18877));
    INVX1 U6006 (.I(N10520), .ZN(n18878));
    INVX1 U6007 (.I(N10521), .ZN(n18879));
    INVX1 U6008 (.I(N10522), .ZN(n18880));
    INVX1 U6009 (.I(N10523), .ZN(N18881));
    INVX1 U6010 (.I(N10524), .ZN(n18882));
    INVX1 U6011 (.I(N10525), .ZN(N18883));
    INVX1 U6012 (.I(N10526), .ZN(N18884));
    INVX1 U6013 (.I(N10527), .ZN(n18885));
    INVX1 U6014 (.I(N10528), .ZN(n18886));
    INVX1 U6015 (.I(N10529), .ZN(N18887));
    INVX1 U6016 (.I(N10530), .ZN(n18888));
    INVX1 U6017 (.I(N10531), .ZN(n18889));
    INVX1 U6018 (.I(N10532), .ZN(n18890));
    INVX1 U6019 (.I(N10533), .ZN(n18891));
    INVX1 U6020 (.I(N10534), .ZN(n18892));
    INVX1 U6021 (.I(N10535), .ZN(n18893));
    INVX1 U6022 (.I(N10536), .ZN(n18894));
    INVX1 U6023 (.I(N10537), .ZN(n18895));
    INVX1 U6024 (.I(N10538), .ZN(n18896));
    INVX1 U6025 (.I(N10539), .ZN(n18897));
    INVX1 U6026 (.I(N10540), .ZN(n18898));
    INVX1 U6027 (.I(N10541), .ZN(N18899));
    INVX1 U6028 (.I(N10542), .ZN(n18900));
    INVX1 U6029 (.I(N10543), .ZN(n18901));
    INVX1 U6030 (.I(N10544), .ZN(n18902));
    INVX1 U6031 (.I(N10545), .ZN(n18903));
    INVX1 U6032 (.I(N10546), .ZN(n18904));
    INVX1 U6033 (.I(N10547), .ZN(n18905));
    INVX1 U6034 (.I(N10548), .ZN(n18906));
    INVX1 U6035 (.I(N10549), .ZN(N18907));
    INVX1 U6036 (.I(N10550), .ZN(n18908));
    INVX1 U6037 (.I(N10551), .ZN(n18909));
    INVX1 U6038 (.I(N10552), .ZN(n18910));
    INVX1 U6039 (.I(N10553), .ZN(n18911));
    INVX1 U6040 (.I(N10554), .ZN(N18912));
    INVX1 U6041 (.I(N10555), .ZN(n18913));
    INVX1 U6042 (.I(N10556), .ZN(n18914));
    INVX1 U6043 (.I(N10557), .ZN(n18915));
    INVX1 U6044 (.I(N10558), .ZN(n18916));
    INVX1 U6045 (.I(N10559), .ZN(n18917));
    INVX1 U6046 (.I(N10560), .ZN(n18918));
    INVX1 U6047 (.I(N10561), .ZN(N18919));
    INVX1 U6048 (.I(N10562), .ZN(n18920));
    INVX1 U6049 (.I(N10563), .ZN(N18921));
    INVX1 U6050 (.I(N10564), .ZN(n18922));
    INVX1 U6051 (.I(N10565), .ZN(n18923));
    INVX1 U6052 (.I(N10566), .ZN(N18924));
    INVX1 U6053 (.I(N10567), .ZN(n18925));
    INVX1 U6054 (.I(N10568), .ZN(n18926));
    INVX1 U6055 (.I(N10569), .ZN(n18927));
    INVX1 U6056 (.I(N10570), .ZN(n18928));
    INVX1 U6057 (.I(N10571), .ZN(N18929));
    INVX1 U6058 (.I(N10572), .ZN(n18930));
    INVX1 U6059 (.I(N10573), .ZN(n18931));
    INVX1 U6060 (.I(N10574), .ZN(n18932));
    INVX1 U6061 (.I(N10575), .ZN(n18933));
    INVX1 U6062 (.I(N10576), .ZN(n18934));
    INVX1 U6063 (.I(N10577), .ZN(n18935));
    INVX1 U6064 (.I(N10578), .ZN(n18936));
    INVX1 U6065 (.I(N10579), .ZN(N18937));
    INVX1 U6066 (.I(N10580), .ZN(n18938));
    INVX1 U6067 (.I(N10581), .ZN(N18939));
    INVX1 U6068 (.I(N10582), .ZN(n18940));
    INVX1 U6069 (.I(N10583), .ZN(n18941));
    INVX1 U6070 (.I(N10584), .ZN(n18942));
    INVX1 U6071 (.I(N10585), .ZN(n18943));
    INVX1 U6072 (.I(N10586), .ZN(N18944));
    INVX1 U6073 (.I(N10587), .ZN(n18945));
    INVX1 U6074 (.I(N10588), .ZN(n18946));
    INVX1 U6075 (.I(N10589), .ZN(n18947));
    INVX1 U6076 (.I(N10590), .ZN(n18948));
    INVX1 U6077 (.I(N10591), .ZN(N18949));
    INVX1 U6078 (.I(N10592), .ZN(n18950));
    INVX1 U6079 (.I(N10593), .ZN(n18951));
    INVX1 U6080 (.I(N10594), .ZN(n18952));
    INVX1 U6081 (.I(N10595), .ZN(n18953));
    INVX1 U6082 (.I(N10596), .ZN(n18954));
    INVX1 U6083 (.I(N10597), .ZN(N18955));
    INVX1 U6084 (.I(N10598), .ZN(n18956));
    INVX1 U6085 (.I(N10599), .ZN(n18957));
    INVX1 U6086 (.I(N10600), .ZN(n18958));
    INVX1 U6087 (.I(N10601), .ZN(n18959));
    INVX1 U6088 (.I(N10602), .ZN(n18960));
    INVX1 U6089 (.I(N10603), .ZN(n18961));
    INVX1 U6090 (.I(N10604), .ZN(n18962));
    INVX1 U6091 (.I(N10605), .ZN(n18963));
    INVX1 U6092 (.I(N10606), .ZN(n18964));
    INVX1 U6093 (.I(N10607), .ZN(n18965));
    INVX1 U6094 (.I(N10608), .ZN(n18966));
    INVX1 U6095 (.I(N10609), .ZN(n18967));
    INVX1 U6096 (.I(N10610), .ZN(n18968));
    INVX1 U6097 (.I(N10611), .ZN(n18969));
    INVX1 U6098 (.I(N10612), .ZN(n18970));
    INVX1 U6099 (.I(N10613), .ZN(N18971));
    INVX1 U6100 (.I(N10614), .ZN(n18972));
    INVX1 U6101 (.I(N10615), .ZN(n18973));
    INVX1 U6102 (.I(N10616), .ZN(n18974));
    INVX1 U6103 (.I(N10617), .ZN(n18975));
    INVX1 U6104 (.I(N10618), .ZN(n18976));
    INVX1 U6105 (.I(N10619), .ZN(n18977));
    INVX1 U6106 (.I(N10620), .ZN(n18978));
    INVX1 U6107 (.I(N10621), .ZN(n18979));
    INVX1 U6108 (.I(N10622), .ZN(N18980));
    INVX1 U6109 (.I(N10623), .ZN(N18981));
    INVX1 U6110 (.I(N10624), .ZN(n18982));
    INVX1 U6111 (.I(N10625), .ZN(N18983));
    INVX1 U6112 (.I(N10626), .ZN(N18984));
    INVX1 U6113 (.I(N10627), .ZN(n18985));
    INVX1 U6114 (.I(N10628), .ZN(n18986));
    INVX1 U6115 (.I(N10629), .ZN(n18987));
    INVX1 U6116 (.I(N10630), .ZN(N18988));
    INVX1 U6117 (.I(N10631), .ZN(n18989));
    INVX1 U6118 (.I(N10632), .ZN(n18990));
    INVX1 U6119 (.I(N10633), .ZN(N18991));
    INVX1 U6120 (.I(N10634), .ZN(n18992));
    INVX1 U6121 (.I(N10635), .ZN(n18993));
    INVX1 U6122 (.I(N10636), .ZN(n18994));
    INVX1 U6123 (.I(N10637), .ZN(n18995));
    INVX1 U6124 (.I(N10638), .ZN(n18996));
    INVX1 U6125 (.I(N10639), .ZN(n18997));
    INVX1 U6126 (.I(N10640), .ZN(n18998));
    INVX1 U6127 (.I(N10641), .ZN(N18999));
    INVX1 U6128 (.I(N10642), .ZN(n19000));
    INVX1 U6129 (.I(N10643), .ZN(n19001));
    INVX1 U6130 (.I(N10644), .ZN(n19002));
    INVX1 U6131 (.I(N10645), .ZN(n19003));
    INVX1 U6132 (.I(N10646), .ZN(n19004));
    INVX1 U6133 (.I(N10647), .ZN(n19005));
    INVX1 U6134 (.I(N10648), .ZN(n19006));
    INVX1 U6135 (.I(N10649), .ZN(N19007));
    INVX1 U6136 (.I(N10650), .ZN(N19008));
    INVX1 U6137 (.I(N10651), .ZN(n19009));
    INVX1 U6138 (.I(N10652), .ZN(n19010));
    INVX1 U6139 (.I(N10653), .ZN(N19011));
    INVX1 U6140 (.I(N10654), .ZN(n19012));
    INVX1 U6141 (.I(N10655), .ZN(n19013));
    INVX1 U6142 (.I(N10656), .ZN(n19014));
    INVX1 U6143 (.I(N10657), .ZN(n19015));
    INVX1 U6144 (.I(N10658), .ZN(n19016));
    INVX1 U6145 (.I(N10659), .ZN(N19017));
    INVX1 U6146 (.I(N10660), .ZN(n19018));
    INVX1 U6147 (.I(N10661), .ZN(n19019));
    INVX1 U6148 (.I(N10662), .ZN(n19020));
    INVX1 U6149 (.I(N10663), .ZN(n19021));
    INVX1 U6150 (.I(N10664), .ZN(n19022));
    INVX1 U6151 (.I(N10665), .ZN(n19023));
    INVX1 U6152 (.I(N10666), .ZN(n19024));
    INVX1 U6153 (.I(N10667), .ZN(n19025));
    INVX1 U6154 (.I(N10668), .ZN(n19026));
    INVX1 U6155 (.I(N10669), .ZN(n19027));
    INVX1 U6156 (.I(N10670), .ZN(n19028));
    INVX1 U6157 (.I(N10671), .ZN(n19029));
    INVX1 U6158 (.I(N10672), .ZN(n19030));
    INVX1 U6159 (.I(N10673), .ZN(n19031));
    INVX1 U6160 (.I(N10674), .ZN(n19032));
    INVX1 U6161 (.I(N10675), .ZN(N19033));
    INVX1 U6162 (.I(N10676), .ZN(n19034));
    INVX1 U6163 (.I(N10677), .ZN(n19035));
    INVX1 U6164 (.I(N10678), .ZN(n19036));
    INVX1 U6165 (.I(N10679), .ZN(n19037));
    INVX1 U6166 (.I(N10680), .ZN(N19038));
    INVX1 U6167 (.I(N10681), .ZN(n19039));
    INVX1 U6168 (.I(N10682), .ZN(n19040));
    INVX1 U6169 (.I(N10683), .ZN(n19041));
    INVX1 U6170 (.I(N10684), .ZN(n19042));
    INVX1 U6171 (.I(N10685), .ZN(n19043));
    INVX1 U6172 (.I(N10686), .ZN(n19044));
    INVX1 U6173 (.I(N10687), .ZN(n19045));
    INVX1 U6174 (.I(N10688), .ZN(n19046));
    INVX1 U6175 (.I(N10689), .ZN(n19047));
    INVX1 U6176 (.I(N10690), .ZN(N19048));
    INVX1 U6177 (.I(N10691), .ZN(n19049));
    INVX1 U6178 (.I(N10692), .ZN(n19050));
    INVX1 U6179 (.I(N10693), .ZN(N19051));
    INVX1 U6180 (.I(N10694), .ZN(n19052));
    INVX1 U6181 (.I(N10695), .ZN(n19053));
    INVX1 U6182 (.I(N10696), .ZN(n19054));
    INVX1 U6183 (.I(N10697), .ZN(n19055));
    INVX1 U6184 (.I(N10698), .ZN(N19056));
    INVX1 U6185 (.I(N10699), .ZN(N19057));
    INVX1 U6186 (.I(N10700), .ZN(N19058));
    INVX1 U6187 (.I(N10701), .ZN(n19059));
    INVX1 U6188 (.I(N10702), .ZN(n19060));
    INVX1 U6189 (.I(N10703), .ZN(n19061));
    INVX1 U6190 (.I(N10704), .ZN(n19062));
    INVX1 U6191 (.I(N10705), .ZN(N19063));
    INVX1 U6192 (.I(N10706), .ZN(n19064));
    INVX1 U6193 (.I(N10707), .ZN(n19065));
    INVX1 U6194 (.I(N10708), .ZN(N19066));
    INVX1 U6195 (.I(N10709), .ZN(n19067));
    INVX1 U6196 (.I(N10710), .ZN(N19068));
    INVX1 U6197 (.I(N10711), .ZN(n19069));
    INVX1 U6198 (.I(N10712), .ZN(N19070));
    INVX1 U6199 (.I(N10713), .ZN(n19071));
    INVX1 U6200 (.I(N10714), .ZN(n19072));
    INVX1 U6201 (.I(N10715), .ZN(n19073));
    INVX1 U6202 (.I(N10716), .ZN(n19074));
    INVX1 U6203 (.I(N10717), .ZN(n19075));
    INVX1 U6204 (.I(N10718), .ZN(N19076));
    INVX1 U6205 (.I(N10719), .ZN(n19077));
    INVX1 U6206 (.I(N10720), .ZN(n19078));
    INVX1 U6207 (.I(N10721), .ZN(n19079));
    INVX1 U6208 (.I(N10722), .ZN(n19080));
    INVX1 U6209 (.I(N10723), .ZN(n19081));
    INVX1 U6210 (.I(N10724), .ZN(n19082));
    INVX1 U6211 (.I(N10725), .ZN(n19083));
    INVX1 U6212 (.I(N10726), .ZN(n19084));
    INVX1 U6213 (.I(N10727), .ZN(n19085));
    INVX1 U6214 (.I(N10728), .ZN(n19086));
    INVX1 U6215 (.I(N10729), .ZN(N19087));
    INVX1 U6216 (.I(N10730), .ZN(N19088));
    INVX1 U6217 (.I(N10731), .ZN(n19089));
    INVX1 U6218 (.I(N10732), .ZN(n19090));
    INVX1 U6219 (.I(N10733), .ZN(n19091));
    INVX1 U6220 (.I(N10734), .ZN(n19092));
    INVX1 U6221 (.I(N10735), .ZN(n19093));
    INVX1 U6222 (.I(N10736), .ZN(n19094));
    INVX1 U6223 (.I(N10737), .ZN(N19095));
    INVX1 U6224 (.I(N10738), .ZN(n19096));
    INVX1 U6225 (.I(N10739), .ZN(N19097));
    INVX1 U6226 (.I(N10740), .ZN(n19098));
    INVX1 U6227 (.I(N10741), .ZN(n19099));
    INVX1 U6228 (.I(N10742), .ZN(N19100));
    INVX1 U6229 (.I(N10743), .ZN(n19101));
    INVX1 U6230 (.I(N10744), .ZN(n19102));
    INVX1 U6231 (.I(N10745), .ZN(n19103));
    INVX1 U6232 (.I(N10746), .ZN(N19104));
    INVX1 U6233 (.I(N10747), .ZN(N19105));
    INVX1 U6234 (.I(N10748), .ZN(n19106));
    INVX1 U6235 (.I(N10749), .ZN(n19107));
    INVX1 U6236 (.I(N10750), .ZN(N19108));
    INVX1 U6237 (.I(N10751), .ZN(N19109));
    INVX1 U6238 (.I(N10752), .ZN(n19110));
    INVX1 U6239 (.I(N10753), .ZN(n19111));
    INVX1 U6240 (.I(N10754), .ZN(N19112));
    INVX1 U6241 (.I(N10755), .ZN(N19113));
    INVX1 U6242 (.I(N10756), .ZN(n19114));
    INVX1 U6243 (.I(N10757), .ZN(n19115));
    INVX1 U6244 (.I(N10758), .ZN(N19116));
    INVX1 U6245 (.I(N10759), .ZN(n19117));
    INVX1 U6246 (.I(N10760), .ZN(n19118));
    INVX1 U6247 (.I(N10761), .ZN(n19119));
    INVX1 U6248 (.I(N10762), .ZN(n19120));
    INVX1 U6249 (.I(N10763), .ZN(n19121));
    INVX1 U6250 (.I(N10764), .ZN(n19122));
    INVX1 U6251 (.I(N10765), .ZN(n19123));
    INVX1 U6252 (.I(N10766), .ZN(n19124));
    INVX1 U6253 (.I(N10767), .ZN(n19125));
    INVX1 U6254 (.I(N10768), .ZN(n19126));
    INVX1 U6255 (.I(N10769), .ZN(n19127));
    INVX1 U6256 (.I(N10770), .ZN(n19128));
    INVX1 U6257 (.I(N10771), .ZN(N19129));
    INVX1 U6258 (.I(N10772), .ZN(N19130));
    INVX1 U6259 (.I(N10773), .ZN(n19131));
    INVX1 U6260 (.I(N10774), .ZN(n19132));
    INVX1 U6261 (.I(N10775), .ZN(n19133));
    INVX1 U6262 (.I(N10776), .ZN(n19134));
    INVX1 U6263 (.I(N10777), .ZN(n19135));
    INVX1 U6264 (.I(N10778), .ZN(n19136));
    INVX1 U6265 (.I(N10779), .ZN(n19137));
    INVX1 U6266 (.I(N10780), .ZN(n19138));
    INVX1 U6267 (.I(N10781), .ZN(N19139));
    INVX1 U6268 (.I(N10782), .ZN(n19140));
    INVX1 U6269 (.I(N10783), .ZN(n19141));
    INVX1 U6270 (.I(N10784), .ZN(n19142));
    INVX1 U6271 (.I(N10785), .ZN(n19143));
    INVX1 U6272 (.I(N10786), .ZN(n19144));
    INVX1 U6273 (.I(N10787), .ZN(n19145));
    INVX1 U6274 (.I(N10788), .ZN(n19146));
    INVX1 U6275 (.I(N10789), .ZN(n19147));
    INVX1 U6276 (.I(N10790), .ZN(n19148));
    INVX1 U6277 (.I(N10791), .ZN(n19149));
    INVX1 U6278 (.I(N10792), .ZN(n19150));
    INVX1 U6279 (.I(N10793), .ZN(n19151));
    INVX1 U6280 (.I(N10794), .ZN(n19152));
    INVX1 U6281 (.I(N10795), .ZN(n19153));
    INVX1 U6282 (.I(N10796), .ZN(n19154));
    INVX1 U6283 (.I(N10797), .ZN(n19155));
    INVX1 U6284 (.I(N10798), .ZN(n19156));
    INVX1 U6285 (.I(N10799), .ZN(n19157));
    INVX1 U6286 (.I(N10800), .ZN(n19158));
    INVX1 U6287 (.I(N10801), .ZN(n19159));
    INVX1 U6288 (.I(N10802), .ZN(N19160));
    INVX1 U6289 (.I(N10803), .ZN(n19161));
    INVX1 U6290 (.I(N10804), .ZN(n19162));
    INVX1 U6291 (.I(N10805), .ZN(n19163));
    INVX1 U6292 (.I(N10806), .ZN(n19164));
    INVX1 U6293 (.I(N10807), .ZN(n19165));
    INVX1 U6294 (.I(N10808), .ZN(n19166));
    INVX1 U6295 (.I(N10809), .ZN(n19167));
    INVX1 U6296 (.I(N10810), .ZN(n19168));
    INVX1 U6297 (.I(N10811), .ZN(n19169));
    INVX1 U6298 (.I(N10812), .ZN(n19170));
    INVX1 U6299 (.I(N10813), .ZN(n19171));
    INVX1 U6300 (.I(N10814), .ZN(n19172));
    INVX1 U6301 (.I(N10815), .ZN(n19173));
    INVX1 U6302 (.I(N10816), .ZN(N19174));
    INVX1 U6303 (.I(N10817), .ZN(N19175));
    INVX1 U6304 (.I(N10818), .ZN(n19176));
    INVX1 U6305 (.I(N10819), .ZN(n19177));
    INVX1 U6306 (.I(N10820), .ZN(N19178));
    INVX1 U6307 (.I(N10821), .ZN(n19179));
    INVX1 U6308 (.I(N10822), .ZN(n19180));
    INVX1 U6309 (.I(N10823), .ZN(n19181));
    INVX1 U6310 (.I(N10824), .ZN(N19182));
    INVX1 U6311 (.I(N10825), .ZN(n19183));
    INVX1 U6312 (.I(N10826), .ZN(n19184));
    INVX1 U6313 (.I(N10827), .ZN(n19185));
    INVX1 U6314 (.I(N10828), .ZN(n19186));
    INVX1 U6315 (.I(N10829), .ZN(N19187));
    INVX1 U6316 (.I(N10830), .ZN(n19188));
    INVX1 U6317 (.I(N10831), .ZN(n19189));
    INVX1 U6318 (.I(N10832), .ZN(N19190));
    INVX1 U6319 (.I(N10833), .ZN(n19191));
    INVX1 U6320 (.I(N10834), .ZN(n19192));
    INVX1 U6321 (.I(N10835), .ZN(n19193));
    INVX1 U6322 (.I(N10836), .ZN(N19194));
    INVX1 U6323 (.I(N10837), .ZN(n19195));
    INVX1 U6324 (.I(N10838), .ZN(n19196));
    INVX1 U6325 (.I(N10839), .ZN(n19197));
    INVX1 U6326 (.I(N10840), .ZN(n19198));
    INVX1 U6327 (.I(N10841), .ZN(n19199));
    INVX1 U6328 (.I(N10842), .ZN(n19200));
    INVX1 U6329 (.I(N10843), .ZN(n19201));
    INVX1 U6330 (.I(N10844), .ZN(n19202));
    INVX1 U6331 (.I(N10845), .ZN(n19203));
    INVX1 U6332 (.I(N10846), .ZN(n19204));
    INVX1 U6333 (.I(N10847), .ZN(n19205));
    INVX1 U6334 (.I(N10848), .ZN(n19206));
    INVX1 U6335 (.I(N10849), .ZN(N19207));
    INVX1 U6336 (.I(N10850), .ZN(n19208));
    INVX1 U6337 (.I(N10851), .ZN(N19209));
    INVX1 U6338 (.I(N10852), .ZN(n19210));
    INVX1 U6339 (.I(N10853), .ZN(n19211));
    INVX1 U6340 (.I(N10854), .ZN(N19212));
    INVX1 U6341 (.I(N10855), .ZN(N19213));
    INVX1 U6342 (.I(N10856), .ZN(n19214));
    INVX1 U6343 (.I(N10857), .ZN(N19215));
    INVX1 U6344 (.I(N10858), .ZN(n19216));
    INVX1 U6345 (.I(N10859), .ZN(n19217));
    INVX1 U6346 (.I(N10860), .ZN(n19218));
    INVX1 U6347 (.I(N10861), .ZN(n19219));
    INVX1 U6348 (.I(N10862), .ZN(N19220));
    INVX1 U6349 (.I(N10863), .ZN(n19221));
    INVX1 U6350 (.I(N10864), .ZN(n19222));
    INVX1 U6351 (.I(N10865), .ZN(n19223));
    INVX1 U6352 (.I(N10866), .ZN(N19224));
    INVX1 U6353 (.I(N10867), .ZN(n19225));
    INVX1 U6354 (.I(N10868), .ZN(n19226));
    INVX1 U6355 (.I(N10869), .ZN(n19227));
    INVX1 U6356 (.I(N10870), .ZN(n19228));
    INVX1 U6357 (.I(N10871), .ZN(n19229));
    INVX1 U6358 (.I(N10872), .ZN(n19230));
    INVX1 U6359 (.I(N10873), .ZN(n19231));
    INVX1 U6360 (.I(N10874), .ZN(n19232));
    INVX1 U6361 (.I(N10875), .ZN(n19233));
    INVX1 U6362 (.I(N10876), .ZN(n19234));
    INVX1 U6363 (.I(N10877), .ZN(n19235));
    INVX1 U6364 (.I(N10878), .ZN(n19236));
    INVX1 U6365 (.I(N10879), .ZN(n19237));
    INVX1 U6366 (.I(N10880), .ZN(n19238));
    INVX1 U6367 (.I(N10881), .ZN(n19239));
    INVX1 U6368 (.I(N10882), .ZN(n19240));
    INVX1 U6369 (.I(N10883), .ZN(N19241));
    INVX1 U6370 (.I(N10884), .ZN(N19242));
    INVX1 U6371 (.I(N10885), .ZN(n19243));
    INVX1 U6372 (.I(N10886), .ZN(n19244));
    INVX1 U6373 (.I(N10887), .ZN(n19245));
    INVX1 U6374 (.I(N10888), .ZN(N19246));
    INVX1 U6375 (.I(N10889), .ZN(N19247));
    INVX1 U6376 (.I(N10890), .ZN(N19248));
    INVX1 U6377 (.I(N10891), .ZN(n19249));
    INVX1 U6378 (.I(N10892), .ZN(n19250));
    INVX1 U6379 (.I(N10893), .ZN(N19251));
    INVX1 U6380 (.I(N10894), .ZN(n19252));
    INVX1 U6381 (.I(N10895), .ZN(n19253));
    INVX1 U6382 (.I(N10896), .ZN(n19254));
    INVX1 U6383 (.I(N10897), .ZN(n19255));
    INVX1 U6384 (.I(N10898), .ZN(n19256));
    INVX1 U6385 (.I(N10899), .ZN(n19257));
    INVX1 U6386 (.I(N10900), .ZN(n19258));
    INVX1 U6387 (.I(N10901), .ZN(n19259));
    INVX1 U6388 (.I(N10902), .ZN(n19260));
    INVX1 U6389 (.I(N10903), .ZN(n19261));
    INVX1 U6390 (.I(N10904), .ZN(n19262));
    INVX1 U6391 (.I(N10905), .ZN(n19263));
    INVX1 U6392 (.I(N10906), .ZN(n19264));
    INVX1 U6393 (.I(N10907), .ZN(N19265));
    INVX1 U6394 (.I(N10908), .ZN(n19266));
    INVX1 U6395 (.I(N10909), .ZN(n19267));
    INVX1 U6396 (.I(N10910), .ZN(n19268));
    INVX1 U6397 (.I(N10911), .ZN(n19269));
    INVX1 U6398 (.I(N10912), .ZN(n19270));
    INVX1 U6399 (.I(N10913), .ZN(n19271));
    INVX1 U6400 (.I(N10914), .ZN(n19272));
    INVX1 U6401 (.I(N10915), .ZN(n19273));
    INVX1 U6402 (.I(N10916), .ZN(N19274));
    INVX1 U6403 (.I(N10917), .ZN(n19275));
    INVX1 U6404 (.I(N10918), .ZN(n19276));
    INVX1 U6405 (.I(N10919), .ZN(N19277));
    INVX1 U6406 (.I(N10920), .ZN(n19278));
    INVX1 U6407 (.I(N10921), .ZN(N19279));
    INVX1 U6408 (.I(N10922), .ZN(n19280));
    INVX1 U6409 (.I(N10923), .ZN(n19281));
    INVX1 U6410 (.I(N10924), .ZN(n19282));
    INVX1 U6411 (.I(N10925), .ZN(n19283));
    INVX1 U6412 (.I(N10926), .ZN(n19284));
    INVX1 U6413 (.I(N10927), .ZN(n19285));
    INVX1 U6414 (.I(N10928), .ZN(n19286));
    INVX1 U6415 (.I(N10929), .ZN(n19287));
    INVX1 U6416 (.I(N10930), .ZN(n19288));
    INVX1 U6417 (.I(N10931), .ZN(n19289));
    INVX1 U6418 (.I(N10932), .ZN(n19290));
    INVX1 U6419 (.I(N10933), .ZN(n19291));
    INVX1 U6420 (.I(N10934), .ZN(n19292));
    INVX1 U6421 (.I(N10935), .ZN(n19293));
    INVX1 U6422 (.I(N10936), .ZN(n19294));
    INVX1 U6423 (.I(N10937), .ZN(n19295));
    INVX1 U6424 (.I(N10938), .ZN(N19296));
    INVX1 U6425 (.I(N10939), .ZN(n19297));
    INVX1 U6426 (.I(N10940), .ZN(n19298));
    INVX1 U6427 (.I(N10941), .ZN(n19299));
    INVX1 U6428 (.I(N10942), .ZN(n19300));
    INVX1 U6429 (.I(N10943), .ZN(n19301));
    INVX1 U6430 (.I(N10944), .ZN(n19302));
    INVX1 U6431 (.I(N10945), .ZN(N19303));
    INVX1 U6432 (.I(N10946), .ZN(n19304));
    INVX1 U6433 (.I(N10947), .ZN(n19305));
    INVX1 U6434 (.I(N10948), .ZN(N19306));
    INVX1 U6435 (.I(N10949), .ZN(n19307));
    INVX1 U6436 (.I(N10950), .ZN(n19308));
    INVX1 U6437 (.I(N10951), .ZN(n19309));
    INVX1 U6438 (.I(N10952), .ZN(n19310));
    INVX1 U6439 (.I(N10953), .ZN(n19311));
    INVX1 U6440 (.I(N10954), .ZN(n19312));
    INVX1 U6441 (.I(N10955), .ZN(n19313));
    INVX1 U6442 (.I(N10956), .ZN(N19314));
    INVX1 U6443 (.I(N10957), .ZN(n19315));
    INVX1 U6444 (.I(N10958), .ZN(n19316));
    INVX1 U6445 (.I(N10959), .ZN(n19317));
    INVX1 U6446 (.I(N10960), .ZN(n19318));
    INVX1 U6447 (.I(N10961), .ZN(n19319));
    INVX1 U6448 (.I(N10962), .ZN(n19320));
    INVX1 U6449 (.I(N10963), .ZN(n19321));
    INVX1 U6450 (.I(N10964), .ZN(n19322));
    INVX1 U6451 (.I(N10965), .ZN(n19323));
    INVX1 U6452 (.I(N10966), .ZN(N19324));
    INVX1 U6453 (.I(N10967), .ZN(n19325));
    INVX1 U6454 (.I(N10968), .ZN(N19326));
    INVX1 U6455 (.I(N10969), .ZN(n19327));
    INVX1 U6456 (.I(N10970), .ZN(n19328));
    INVX1 U6457 (.I(N10971), .ZN(N19329));
    INVX1 U6458 (.I(N10972), .ZN(n19330));
    INVX1 U6459 (.I(N10973), .ZN(n19331));
    INVX1 U6460 (.I(N10974), .ZN(n19332));
    INVX1 U6461 (.I(N10975), .ZN(n19333));
    INVX1 U6462 (.I(N10976), .ZN(N19334));
    INVX1 U6463 (.I(N10977), .ZN(n19335));
    INVX1 U6464 (.I(N10978), .ZN(n19336));
    INVX1 U6465 (.I(N10979), .ZN(n19337));
    INVX1 U6466 (.I(N10980), .ZN(n19338));
    INVX1 U6467 (.I(N10981), .ZN(n19339));
    INVX1 U6468 (.I(N10982), .ZN(N19340));
    INVX1 U6469 (.I(N10983), .ZN(N19341));
    INVX1 U6470 (.I(N10984), .ZN(n19342));
    INVX1 U6471 (.I(N10985), .ZN(n19343));
    INVX1 U6472 (.I(N10986), .ZN(n19344));
    INVX1 U6473 (.I(N10987), .ZN(n19345));
    INVX1 U6474 (.I(N10988), .ZN(N19346));
    INVX1 U6475 (.I(N10989), .ZN(N19347));
    INVX1 U6476 (.I(N10990), .ZN(n19348));
    INVX1 U6477 (.I(N10991), .ZN(n19349));
    INVX1 U6478 (.I(N10992), .ZN(N19350));
    INVX1 U6479 (.I(N10993), .ZN(n19351));
    INVX1 U6480 (.I(N10994), .ZN(n19352));
    INVX1 U6481 (.I(N10995), .ZN(n19353));
    INVX1 U6482 (.I(N10996), .ZN(n19354));
    INVX1 U6483 (.I(N10997), .ZN(n19355));
    INVX1 U6484 (.I(N10998), .ZN(n19356));
    INVX1 U6485 (.I(N10999), .ZN(n19357));
    INVX1 U6486 (.I(N11000), .ZN(n19358));
    INVX1 U6487 (.I(N11001), .ZN(n19359));
    INVX1 U6488 (.I(N11002), .ZN(n19360));
    INVX1 U6489 (.I(N11003), .ZN(n19361));
    INVX1 U6490 (.I(N11004), .ZN(n19362));
    INVX1 U6491 (.I(N11005), .ZN(n19363));
    INVX1 U6492 (.I(N11006), .ZN(n19364));
    INVX1 U6493 (.I(N11007), .ZN(n19365));
    INVX1 U6494 (.I(N11008), .ZN(n19366));
    INVX1 U6495 (.I(N11009), .ZN(n19367));
    INVX1 U6496 (.I(N11010), .ZN(n19368));
    INVX1 U6497 (.I(N11011), .ZN(n19369));
    INVX1 U6498 (.I(N11012), .ZN(n19370));
    INVX1 U6499 (.I(N11013), .ZN(n19371));
    INVX1 U6500 (.I(N11014), .ZN(n19372));
    INVX1 U6501 (.I(N11015), .ZN(n19373));
    INVX1 U6502 (.I(N11016), .ZN(n19374));
    INVX1 U6503 (.I(N11017), .ZN(N19375));
    INVX1 U6504 (.I(N11018), .ZN(n19376));
    INVX1 U6505 (.I(N11019), .ZN(n19377));
    INVX1 U6506 (.I(N11020), .ZN(n19378));
    INVX1 U6507 (.I(N11021), .ZN(n19379));
    INVX1 U6508 (.I(N11022), .ZN(N19380));
    INVX1 U6509 (.I(N11023), .ZN(n19381));
    INVX1 U6510 (.I(N11024), .ZN(n19382));
    INVX1 U6511 (.I(N11025), .ZN(n19383));
    INVX1 U6512 (.I(N11026), .ZN(n19384));
    INVX1 U6513 (.I(N11027), .ZN(n19385));
    INVX1 U6514 (.I(N11028), .ZN(N19386));
    INVX1 U6515 (.I(N11029), .ZN(n19387));
    INVX1 U6516 (.I(N11030), .ZN(N19388));
    INVX1 U6517 (.I(N11031), .ZN(n19389));
    INVX1 U6518 (.I(N11032), .ZN(n19390));
    INVX1 U6519 (.I(N11033), .ZN(n19391));
    INVX1 U6520 (.I(N11034), .ZN(n19392));
    INVX1 U6521 (.I(N11035), .ZN(n19393));
    INVX1 U6522 (.I(N11036), .ZN(n19394));
    INVX1 U6523 (.I(N11037), .ZN(n19395));
    INVX1 U6524 (.I(N11038), .ZN(n19396));
    INVX1 U6525 (.I(N11039), .ZN(n19397));
    INVX1 U6526 (.I(N11040), .ZN(n19398));
    INVX1 U6527 (.I(N11041), .ZN(N19399));
    INVX1 U6528 (.I(N11042), .ZN(n19400));
    INVX1 U6529 (.I(N11043), .ZN(n19401));
    INVX1 U6530 (.I(N11044), .ZN(N19402));
    INVX1 U6531 (.I(N11045), .ZN(n19403));
    INVX1 U6532 (.I(N11046), .ZN(n19404));
    INVX1 U6533 (.I(N11047), .ZN(n19405));
    INVX1 U6534 (.I(N11048), .ZN(n19406));
    INVX1 U6535 (.I(N11049), .ZN(n19407));
    INVX1 U6536 (.I(N11050), .ZN(n19408));
    INVX1 U6537 (.I(N11051), .ZN(N19409));
    INVX1 U6538 (.I(N11052), .ZN(n19410));
    INVX1 U6539 (.I(N11053), .ZN(n19411));
    INVX1 U6540 (.I(N11054), .ZN(n19412));
    INVX1 U6541 (.I(N11055), .ZN(n19413));
    INVX1 U6542 (.I(N11056), .ZN(n19414));
    INVX1 U6543 (.I(N11057), .ZN(n19415));
    INVX1 U6544 (.I(N11058), .ZN(n19416));
    INVX1 U6545 (.I(N11059), .ZN(n19417));
    INVX1 U6546 (.I(N11060), .ZN(n19418));
    INVX1 U6547 (.I(N11061), .ZN(n19419));
    INVX1 U6548 (.I(N11062), .ZN(n19420));
    INVX1 U6549 (.I(N11063), .ZN(n19421));
    INVX1 U6550 (.I(N11064), .ZN(n19422));
    INVX1 U6551 (.I(N11065), .ZN(n19423));
    INVX1 U6552 (.I(N11066), .ZN(n19424));
    INVX1 U6553 (.I(N11067), .ZN(n19425));
    INVX1 U6554 (.I(N11068), .ZN(n19426));
    INVX1 U6555 (.I(N11069), .ZN(n19427));
    INVX1 U6556 (.I(N11070), .ZN(n19428));
    INVX1 U6557 (.I(N11071), .ZN(n19429));
    INVX1 U6558 (.I(N11072), .ZN(N19430));
    INVX1 U6559 (.I(N11073), .ZN(n19431));
    INVX1 U6560 (.I(N11074), .ZN(n19432));
    INVX1 U6561 (.I(N11075), .ZN(n19433));
    INVX1 U6562 (.I(N11076), .ZN(n19434));
    INVX1 U6563 (.I(N11077), .ZN(n19435));
    INVX1 U6564 (.I(N11078), .ZN(n19436));
    INVX1 U6565 (.I(N11079), .ZN(n19437));
    INVX1 U6566 (.I(N11080), .ZN(n19438));
    INVX1 U6567 (.I(N11081), .ZN(n19439));
    INVX1 U6568 (.I(N11082), .ZN(n19440));
    INVX1 U6569 (.I(N11083), .ZN(n19441));
    INVX1 U6570 (.I(N11084), .ZN(n19442));
    INVX1 U6571 (.I(N11085), .ZN(n19443));
    INVX1 U6572 (.I(N11086), .ZN(n19444));
    INVX1 U6573 (.I(N11087), .ZN(N19445));
    INVX1 U6574 (.I(N11088), .ZN(n19446));
    INVX1 U6575 (.I(N11089), .ZN(N19447));
    INVX1 U6576 (.I(N11090), .ZN(n19448));
    INVX1 U6577 (.I(N11091), .ZN(n19449));
    INVX1 U6578 (.I(N11092), .ZN(n19450));
    INVX1 U6579 (.I(N11093), .ZN(n19451));
    INVX1 U6580 (.I(N11094), .ZN(n19452));
    INVX1 U6581 (.I(N11095), .ZN(n19453));
    INVX1 U6582 (.I(N11096), .ZN(n19454));
    INVX1 U6583 (.I(N11097), .ZN(n19455));
    INVX1 U6584 (.I(N11098), .ZN(n19456));
    INVX1 U6585 (.I(N11099), .ZN(N19457));
    INVX1 U6586 (.I(N11100), .ZN(n19458));
    INVX1 U6587 (.I(N11101), .ZN(N19459));
    INVX1 U6588 (.I(N11102), .ZN(n19460));
    INVX1 U6589 (.I(N11103), .ZN(n19461));
    INVX1 U6590 (.I(N11104), .ZN(n19462));
    INVX1 U6591 (.I(N11105), .ZN(n19463));
    INVX1 U6592 (.I(N11106), .ZN(n19464));
    INVX1 U6593 (.I(N11107), .ZN(n19465));
    INVX1 U6594 (.I(N11108), .ZN(n19466));
    INVX1 U6595 (.I(N11109), .ZN(n19467));
    INVX1 U6596 (.I(N11110), .ZN(n19468));
    INVX1 U6597 (.I(N11111), .ZN(n19469));
    INVX1 U6598 (.I(N11112), .ZN(n19470));
    INVX1 U6599 (.I(N11113), .ZN(n19471));
    INVX1 U6600 (.I(N11114), .ZN(n19472));
    INVX1 U6601 (.I(N11115), .ZN(n19473));
    INVX1 U6602 (.I(N11116), .ZN(N19474));
    INVX1 U6603 (.I(N11117), .ZN(n19475));
    INVX1 U6604 (.I(N11118), .ZN(n19476));
    INVX1 U6605 (.I(N11119), .ZN(n19477));
    INVX1 U6606 (.I(N11120), .ZN(n19478));
    INVX1 U6607 (.I(N11121), .ZN(n19479));
    INVX1 U6608 (.I(N11122), .ZN(n19480));
    INVX1 U6609 (.I(N11123), .ZN(N19481));
    INVX1 U6610 (.I(N11124), .ZN(N19482));
    INVX1 U6611 (.I(N11125), .ZN(n19483));
    INVX1 U6612 (.I(N11126), .ZN(N19484));
    INVX1 U6613 (.I(N11127), .ZN(n19485));
    INVX1 U6614 (.I(N11128), .ZN(n19486));
    INVX1 U6615 (.I(N11129), .ZN(n19487));
    INVX1 U6616 (.I(N11130), .ZN(n19488));
    INVX1 U6617 (.I(N11131), .ZN(n19489));
    INVX1 U6618 (.I(N11132), .ZN(n19490));
    INVX1 U6619 (.I(N11133), .ZN(n19491));
    INVX1 U6620 (.I(N11134), .ZN(n19492));
    INVX1 U6621 (.I(N11135), .ZN(N19493));
    INVX1 U6622 (.I(N11136), .ZN(n19494));
    INVX1 U6623 (.I(N11137), .ZN(n19495));
    INVX1 U6624 (.I(N11138), .ZN(n19496));
    INVX1 U6625 (.I(N11139), .ZN(n19497));
    INVX1 U6626 (.I(N11140), .ZN(n19498));
    INVX1 U6627 (.I(N11141), .ZN(N19499));
    INVX1 U6628 (.I(N11142), .ZN(n19500));
    INVX1 U6629 (.I(N11143), .ZN(n19501));
    INVX1 U6630 (.I(N11144), .ZN(n19502));
    INVX1 U6631 (.I(N11145), .ZN(n19503));
    INVX1 U6632 (.I(N11146), .ZN(n19504));
    INVX1 U6633 (.I(N11147), .ZN(n19505));
    INVX1 U6634 (.I(N11148), .ZN(n19506));
    INVX1 U6635 (.I(N11149), .ZN(n19507));
    INVX1 U6636 (.I(N11150), .ZN(n19508));
    INVX1 U6637 (.I(N11151), .ZN(n19509));
    INVX1 U6638 (.I(N11152), .ZN(n19510));
    INVX1 U6639 (.I(N11153), .ZN(n19511));
    INVX1 U6640 (.I(N11154), .ZN(n19512));
    INVX1 U6641 (.I(N11155), .ZN(n19513));
    INVX1 U6642 (.I(N11156), .ZN(n19514));
    INVX1 U6643 (.I(N11157), .ZN(n19515));
    INVX1 U6644 (.I(N11158), .ZN(n19516));
    INVX1 U6645 (.I(N11159), .ZN(n19517));
    INVX1 U6646 (.I(N11160), .ZN(n19518));
    INVX1 U6647 (.I(N11161), .ZN(n19519));
    INVX1 U6648 (.I(N11162), .ZN(n19520));
    INVX1 U6649 (.I(N11163), .ZN(n19521));
    INVX1 U6650 (.I(N11164), .ZN(n19522));
    INVX1 U6651 (.I(N11165), .ZN(n19523));
    INVX1 U6652 (.I(N11166), .ZN(N19524));
    INVX1 U6653 (.I(N11167), .ZN(n19525));
    INVX1 U6654 (.I(N11168), .ZN(n19526));
    INVX1 U6655 (.I(N11169), .ZN(N19527));
    INVX1 U6656 (.I(N11170), .ZN(n19528));
    INVX1 U6657 (.I(N11171), .ZN(n19529));
    INVX1 U6658 (.I(N11172), .ZN(n19530));
    INVX1 U6659 (.I(N11173), .ZN(N19531));
    INVX1 U6660 (.I(N11174), .ZN(N19532));
    INVX1 U6661 (.I(N11175), .ZN(n19533));
    INVX1 U6662 (.I(N11176), .ZN(N19534));
    INVX1 U6663 (.I(N11177), .ZN(n19535));
    INVX1 U6664 (.I(N11178), .ZN(N19536));
    INVX1 U6665 (.I(N11179), .ZN(N19537));
    INVX1 U6666 (.I(N11180), .ZN(n19538));
    INVX1 U6667 (.I(N11181), .ZN(n19539));
    INVX1 U6668 (.I(N11182), .ZN(n19540));
    INVX1 U6669 (.I(N11183), .ZN(n19541));
    INVX1 U6670 (.I(N11184), .ZN(n19542));
    INVX1 U6671 (.I(N11185), .ZN(N19543));
    INVX1 U6672 (.I(N11186), .ZN(n19544));
    INVX1 U6673 (.I(N11187), .ZN(n19545));
    INVX1 U6674 (.I(N11188), .ZN(n19546));
    INVX1 U6675 (.I(N11189), .ZN(n19547));
    INVX1 U6676 (.I(N11190), .ZN(n19548));
    INVX1 U6677 (.I(N11191), .ZN(N19549));
    INVX1 U6678 (.I(N11192), .ZN(n19550));
    INVX1 U6679 (.I(N11193), .ZN(n19551));
    INVX1 U6680 (.I(N11194), .ZN(n19552));
    INVX1 U6681 (.I(N11195), .ZN(n19553));
    INVX1 U6682 (.I(N11196), .ZN(n19554));
    INVX1 U6683 (.I(N11197), .ZN(n19555));
    INVX1 U6684 (.I(N11198), .ZN(n19556));
    INVX1 U6685 (.I(N11199), .ZN(n19557));
    INVX1 U6686 (.I(N11200), .ZN(n19558));
    INVX1 U6687 (.I(N11201), .ZN(n19559));
    INVX1 U6688 (.I(N11202), .ZN(n19560));
    INVX1 U6689 (.I(N11203), .ZN(N19561));
    INVX1 U6690 (.I(N11204), .ZN(n19562));
    INVX1 U6691 (.I(N11205), .ZN(n19563));
    INVX1 U6692 (.I(N11206), .ZN(N19564));
    INVX1 U6693 (.I(N11207), .ZN(n19565));
    INVX1 U6694 (.I(N11208), .ZN(n19566));
    INVX1 U6695 (.I(N11209), .ZN(N19567));
    INVX1 U6696 (.I(N11210), .ZN(N19568));
    INVX1 U6697 (.I(N11211), .ZN(n19569));
    INVX1 U6698 (.I(N11212), .ZN(N19570));
    INVX1 U6699 (.I(N11213), .ZN(n19571));
    INVX1 U6700 (.I(N11214), .ZN(n19572));
    INVX1 U6701 (.I(N11215), .ZN(n19573));
    INVX1 U6702 (.I(N11216), .ZN(n19574));
    INVX1 U6703 (.I(N11217), .ZN(n19575));
    INVX1 U6704 (.I(N11218), .ZN(n19576));
    INVX1 U6705 (.I(N11219), .ZN(N19577));
    INVX1 U6706 (.I(N11220), .ZN(n19578));
    INVX1 U6707 (.I(N11221), .ZN(n19579));
    INVX1 U6708 (.I(N11222), .ZN(n19580));
    INVX1 U6709 (.I(N11223), .ZN(n19581));
    INVX1 U6710 (.I(N11224), .ZN(n19582));
    INVX1 U6711 (.I(N11225), .ZN(N19583));
    INVX1 U6712 (.I(N11226), .ZN(n19584));
    INVX1 U6713 (.I(N11227), .ZN(N19585));
    INVX1 U6714 (.I(N11228), .ZN(n19586));
    INVX1 U6715 (.I(N11229), .ZN(n19587));
    INVX1 U6716 (.I(N11230), .ZN(n19588));
    INVX1 U6717 (.I(N11231), .ZN(n19589));
    INVX1 U6718 (.I(N11232), .ZN(n19590));
    INVX1 U6719 (.I(N11233), .ZN(n19591));
    INVX1 U6720 (.I(N11234), .ZN(n19592));
    INVX1 U6721 (.I(N11235), .ZN(N19593));
    INVX1 U6722 (.I(N11236), .ZN(n19594));
    INVX1 U6723 (.I(N11237), .ZN(n19595));
    INVX1 U6724 (.I(N11238), .ZN(N19596));
    INVX1 U6725 (.I(N11239), .ZN(n19597));
    INVX1 U6726 (.I(N11240), .ZN(n19598));
    INVX1 U6727 (.I(N11241), .ZN(n19599));
    INVX1 U6728 (.I(N11242), .ZN(n19600));
    INVX1 U6729 (.I(N11243), .ZN(n19601));
    INVX1 U6730 (.I(N11244), .ZN(n19602));
    INVX1 U6731 (.I(N11245), .ZN(n19603));
    INVX1 U6732 (.I(N11246), .ZN(n19604));
    INVX1 U6733 (.I(N11247), .ZN(n19605));
    INVX1 U6734 (.I(N11248), .ZN(n19606));
    INVX1 U6735 (.I(N11249), .ZN(n19607));
    INVX1 U6736 (.I(N11250), .ZN(n19608));
    INVX1 U6737 (.I(N11251), .ZN(n19609));
    INVX1 U6738 (.I(N11252), .ZN(n19610));
    INVX1 U6739 (.I(N11253), .ZN(n19611));
    INVX1 U6740 (.I(N11254), .ZN(n19612));
    INVX1 U6741 (.I(N11255), .ZN(n19613));
    INVX1 U6742 (.I(N11256), .ZN(n19614));
    INVX1 U6743 (.I(N11257), .ZN(n19615));
    INVX1 U6744 (.I(N11258), .ZN(n19616));
    INVX1 U6745 (.I(N11259), .ZN(N19617));
    INVX1 U6746 (.I(N11260), .ZN(n19618));
    INVX1 U6747 (.I(N11261), .ZN(n19619));
    INVX1 U6748 (.I(N11262), .ZN(n19620));
    INVX1 U6749 (.I(N11263), .ZN(n19621));
    INVX1 U6750 (.I(N11264), .ZN(N19622));
    INVX1 U6751 (.I(N11265), .ZN(N19623));
    INVX1 U6752 (.I(N11266), .ZN(n19624));
    INVX1 U6753 (.I(N11267), .ZN(n19625));
    INVX1 U6754 (.I(N11268), .ZN(n19626));
    INVX1 U6755 (.I(N11269), .ZN(n19627));
    INVX1 U6756 (.I(N11270), .ZN(n19628));
    INVX1 U6757 (.I(N11271), .ZN(n19629));
    INVX1 U6758 (.I(N11272), .ZN(N19630));
    INVX1 U6759 (.I(N11273), .ZN(n19631));
    INVX1 U6760 (.I(N11274), .ZN(n19632));
    INVX1 U6761 (.I(N11275), .ZN(N19633));
    INVX1 U6762 (.I(N11276), .ZN(n19634));
    INVX1 U6763 (.I(N11277), .ZN(n19635));
    INVX1 U6764 (.I(N11278), .ZN(n19636));
    INVX1 U6765 (.I(N11279), .ZN(n19637));
    INVX1 U6766 (.I(N11280), .ZN(n19638));
    INVX1 U6767 (.I(N11281), .ZN(n19639));
    INVX1 U6768 (.I(N11282), .ZN(n19640));
    INVX1 U6769 (.I(N11283), .ZN(n19641));
    INVX1 U6770 (.I(N11284), .ZN(n19642));
    INVX1 U6771 (.I(N11285), .ZN(n19643));
    INVX1 U6772 (.I(N11286), .ZN(n19644));
    INVX1 U6773 (.I(N11287), .ZN(n19645));
    INVX1 U6774 (.I(N11288), .ZN(n19646));
    INVX1 U6775 (.I(N11289), .ZN(n19647));
    INVX1 U6776 (.I(N11290), .ZN(n19648));
    INVX1 U6777 (.I(N11291), .ZN(n19649));
    INVX1 U6778 (.I(N11292), .ZN(n19650));
    INVX1 U6779 (.I(N11293), .ZN(n19651));
    INVX1 U6780 (.I(N11294), .ZN(n19652));
    INVX1 U6781 (.I(N11295), .ZN(n19653));
    INVX1 U6782 (.I(N11296), .ZN(n19654));
    INVX1 U6783 (.I(N11297), .ZN(n19655));
    INVX1 U6784 (.I(N11298), .ZN(n19656));
    INVX1 U6785 (.I(N11299), .ZN(N19657));
    INVX1 U6786 (.I(N11300), .ZN(N19658));
    INVX1 U6787 (.I(N11301), .ZN(n19659));
    INVX1 U6788 (.I(N11302), .ZN(n19660));
    INVX1 U6789 (.I(N11303), .ZN(n19661));
    INVX1 U6790 (.I(N11304), .ZN(n19662));
    INVX1 U6791 (.I(N11305), .ZN(n19663));
    INVX1 U6792 (.I(N11306), .ZN(n19664));
    INVX1 U6793 (.I(N11307), .ZN(n19665));
    INVX1 U6794 (.I(N11308), .ZN(n19666));
    INVX1 U6795 (.I(N11309), .ZN(n19667));
    INVX1 U6796 (.I(N11310), .ZN(N19668));
    INVX1 U6797 (.I(N11311), .ZN(n19669));
    INVX1 U6798 (.I(N11312), .ZN(N19670));
    INVX1 U6799 (.I(N11313), .ZN(n19671));
    INVX1 U6800 (.I(N11314), .ZN(n19672));
    INVX1 U6801 (.I(N11315), .ZN(N19673));
    INVX1 U6802 (.I(N11316), .ZN(n19674));
    INVX1 U6803 (.I(N11317), .ZN(n19675));
    INVX1 U6804 (.I(N11318), .ZN(N19676));
    INVX1 U6805 (.I(N11319), .ZN(n19677));
    INVX1 U6806 (.I(N11320), .ZN(N19678));
    INVX1 U6807 (.I(N11321), .ZN(n19679));
    INVX1 U6808 (.I(N11322), .ZN(n19680));
    INVX1 U6809 (.I(N11323), .ZN(n19681));
    INVX1 U6810 (.I(N11324), .ZN(n19682));
    INVX1 U6811 (.I(N11325), .ZN(n19683));
    INVX1 U6812 (.I(N11326), .ZN(n19684));
    INVX1 U6813 (.I(N11327), .ZN(n19685));
    INVX1 U6814 (.I(N11328), .ZN(N19686));
    INVX1 U6815 (.I(N11329), .ZN(n19687));
    INVX1 U6816 (.I(N11330), .ZN(n19688));
    INVX1 U6817 (.I(N11331), .ZN(n19689));
    INVX1 U6818 (.I(N11332), .ZN(n19690));
    INVX1 U6819 (.I(N11333), .ZN(n19691));
    INVX1 U6820 (.I(N11334), .ZN(n19692));
    INVX1 U6821 (.I(N11335), .ZN(N19693));
    INVX1 U6822 (.I(N11336), .ZN(n19694));
    INVX1 U6823 (.I(N11337), .ZN(n19695));
    INVX1 U6824 (.I(N11338), .ZN(N19696));
    INVX1 U6825 (.I(N11339), .ZN(n19697));
    INVX1 U6826 (.I(N11340), .ZN(n19698));
    INVX1 U6827 (.I(N11341), .ZN(n19699));
    INVX1 U6828 (.I(N11342), .ZN(n19700));
    INVX1 U6829 (.I(N11343), .ZN(n19701));
    INVX1 U6830 (.I(N11344), .ZN(n19702));
    INVX1 U6831 (.I(N11345), .ZN(n19703));
    INVX1 U6832 (.I(N11346), .ZN(n19704));
    INVX1 U6833 (.I(N11347), .ZN(n19705));
    INVX1 U6834 (.I(N11348), .ZN(n19706));
    INVX1 U6835 (.I(N11349), .ZN(n19707));
    INVX1 U6836 (.I(N11350), .ZN(n19708));
    INVX1 U6837 (.I(N11351), .ZN(n19709));
    INVX1 U6838 (.I(N11352), .ZN(n19710));
    INVX1 U6839 (.I(N11353), .ZN(n19711));
    INVX1 U6840 (.I(N11354), .ZN(n19712));
    INVX1 U6841 (.I(N11355), .ZN(n19713));
    INVX1 U6842 (.I(N11356), .ZN(N19714));
    INVX1 U6843 (.I(N11357), .ZN(n19715));
    INVX1 U6844 (.I(N11358), .ZN(n19716));
    INVX1 U6845 (.I(N11359), .ZN(n19717));
    INVX1 U6846 (.I(N11360), .ZN(n19718));
    INVX1 U6847 (.I(N11361), .ZN(n19719));
    INVX1 U6848 (.I(N11362), .ZN(n19720));
    INVX1 U6849 (.I(N11363), .ZN(n19721));
    INVX1 U6850 (.I(N11364), .ZN(n19722));
    INVX1 U6851 (.I(N11365), .ZN(n19723));
    INVX1 U6852 (.I(N11366), .ZN(n19724));
    INVX1 U6853 (.I(N11367), .ZN(n19725));
    INVX1 U6854 (.I(N11368), .ZN(n19726));
    INVX1 U6855 (.I(N11369), .ZN(n19727));
    INVX1 U6856 (.I(N11370), .ZN(n19728));
    INVX1 U6857 (.I(N11371), .ZN(N19729));
    INVX1 U6858 (.I(N11372), .ZN(n19730));
    INVX1 U6859 (.I(N11373), .ZN(n19731));
    INVX1 U6860 (.I(N11374), .ZN(n19732));
    INVX1 U6861 (.I(N11375), .ZN(n19733));
    INVX1 U6862 (.I(N11376), .ZN(n19734));
    INVX1 U6863 (.I(N11377), .ZN(n19735));
    INVX1 U6864 (.I(N11378), .ZN(n19736));
    INVX1 U6865 (.I(N11379), .ZN(n19737));
    INVX1 U6866 (.I(N11380), .ZN(n19738));
    INVX1 U6867 (.I(N11381), .ZN(n19739));
    INVX1 U6868 (.I(N11382), .ZN(n19740));
    INVX1 U6869 (.I(N11383), .ZN(n19741));
    INVX1 U6870 (.I(N11384), .ZN(n19742));
    INVX1 U6871 (.I(N11385), .ZN(N19743));
    INVX1 U6872 (.I(N11386), .ZN(N19744));
    INVX1 U6873 (.I(N11387), .ZN(n19745));
    INVX1 U6874 (.I(N11388), .ZN(N19746));
    INVX1 U6875 (.I(N11389), .ZN(N19747));
    INVX1 U6876 (.I(N11390), .ZN(N19748));
    INVX1 U6877 (.I(N11391), .ZN(n19749));
    INVX1 U6878 (.I(N11392), .ZN(n19750));
    INVX1 U6879 (.I(N11393), .ZN(N19751));
    INVX1 U6880 (.I(N11394), .ZN(n19752));
    INVX1 U6881 (.I(N11395), .ZN(n19753));
    INVX1 U6882 (.I(N11396), .ZN(n19754));
    INVX1 U6883 (.I(N11397), .ZN(n19755));
    INVX1 U6884 (.I(N11398), .ZN(n19756));
    INVX1 U6885 (.I(N11399), .ZN(n19757));
    INVX1 U6886 (.I(N11400), .ZN(n19758));
    INVX1 U6887 (.I(N11401), .ZN(n19759));
    INVX1 U6888 (.I(N11402), .ZN(n19760));
    INVX1 U6889 (.I(N11403), .ZN(n19761));
    INVX1 U6890 (.I(N11404), .ZN(n19762));
    INVX1 U6891 (.I(N11405), .ZN(N19763));
    INVX1 U6892 (.I(N11406), .ZN(n19764));
    INVX1 U6893 (.I(N11407), .ZN(n19765));
    INVX1 U6894 (.I(N11408), .ZN(n19766));
    INVX1 U6895 (.I(N11409), .ZN(n19767));
    INVX1 U6896 (.I(N11410), .ZN(n19768));
    INVX1 U6897 (.I(N11411), .ZN(n19769));
    INVX1 U6898 (.I(N11412), .ZN(n19770));
    INVX1 U6899 (.I(N11413), .ZN(n19771));
    INVX1 U6900 (.I(N11414), .ZN(n19772));
    INVX1 U6901 (.I(N11415), .ZN(n19773));
    INVX1 U6902 (.I(N11416), .ZN(n19774));
    INVX1 U6903 (.I(N11417), .ZN(n19775));
    INVX1 U6904 (.I(N11418), .ZN(n19776));
    INVX1 U6905 (.I(N11419), .ZN(n19777));
    INVX1 U6906 (.I(N11420), .ZN(n19778));
    INVX1 U6907 (.I(N11421), .ZN(n19779));
    INVX1 U6908 (.I(N11422), .ZN(N19780));
    INVX1 U6909 (.I(N11423), .ZN(n19781));
    INVX1 U6910 (.I(N11424), .ZN(n19782));
    INVX1 U6911 (.I(N11425), .ZN(n19783));
    INVX1 U6912 (.I(N11426), .ZN(n19784));
    INVX1 U6913 (.I(N11427), .ZN(N19785));
    INVX1 U6914 (.I(N11428), .ZN(n19786));
    INVX1 U6915 (.I(N11429), .ZN(n19787));
    INVX1 U6916 (.I(N11430), .ZN(n19788));
    INVX1 U6917 (.I(N11431), .ZN(n19789));
    INVX1 U6918 (.I(N11432), .ZN(n19790));
    INVX1 U6919 (.I(N11433), .ZN(n19791));
    INVX1 U6920 (.I(N11434), .ZN(n19792));
    INVX1 U6921 (.I(N11435), .ZN(n19793));
    INVX1 U6922 (.I(N11436), .ZN(n19794));
    INVX1 U6923 (.I(N11437), .ZN(n19795));
    INVX1 U6924 (.I(N11438), .ZN(n19796));
    INVX1 U6925 (.I(N11439), .ZN(n19797));
    INVX1 U6926 (.I(N11440), .ZN(n19798));
    INVX1 U6927 (.I(N11441), .ZN(n19799));
    INVX1 U6928 (.I(N11442), .ZN(n19800));
    INVX1 U6929 (.I(N11443), .ZN(n19801));
    INVX1 U6930 (.I(N11444), .ZN(n19802));
    INVX1 U6931 (.I(N11445), .ZN(n19803));
    INVX1 U6932 (.I(N11446), .ZN(n19804));
    INVX1 U6933 (.I(N11447), .ZN(n19805));
    INVX1 U6934 (.I(N11448), .ZN(n19806));
    INVX1 U6935 (.I(N11449), .ZN(n19807));
    INVX1 U6936 (.I(N11450), .ZN(n19808));
    INVX1 U6937 (.I(N11451), .ZN(n19809));
    INVX1 U6938 (.I(N11452), .ZN(n19810));
    INVX1 U6939 (.I(N11453), .ZN(n19811));
    INVX1 U6940 (.I(N11454), .ZN(n19812));
    INVX1 U6941 (.I(N11455), .ZN(n19813));
    INVX1 U6942 (.I(N11456), .ZN(n19814));
    INVX1 U6943 (.I(N11457), .ZN(n19815));
    INVX1 U6944 (.I(N11458), .ZN(N19816));
    INVX1 U6945 (.I(N11459), .ZN(n19817));
    INVX1 U6946 (.I(N11460), .ZN(n19818));
    INVX1 U6947 (.I(N11461), .ZN(N19819));
    INVX1 U6948 (.I(N11462), .ZN(n19820));
    INVX1 U6949 (.I(N11463), .ZN(n19821));
    INVX1 U6950 (.I(N11464), .ZN(N19822));
    INVX1 U6951 (.I(N11465), .ZN(N19823));
    INVX1 U6952 (.I(N11466), .ZN(N19824));
    INVX1 U6953 (.I(N11467), .ZN(n19825));
    INVX1 U6954 (.I(N11468), .ZN(n19826));
    INVX1 U6955 (.I(N11469), .ZN(n19827));
    INVX1 U6956 (.I(N11470), .ZN(n19828));
    INVX1 U6957 (.I(N11471), .ZN(N19829));
    INVX1 U6958 (.I(N11472), .ZN(n19830));
    INVX1 U6959 (.I(N11473), .ZN(n19831));
    INVX1 U6960 (.I(N11474), .ZN(N19832));
    INVX1 U6961 (.I(N11475), .ZN(n19833));
    INVX1 U6962 (.I(N11476), .ZN(n19834));
    INVX1 U6963 (.I(N11477), .ZN(n19835));
    INVX1 U6964 (.I(N11478), .ZN(n19836));
    INVX1 U6965 (.I(N11479), .ZN(n19837));
    INVX1 U6966 (.I(N11480), .ZN(n19838));
    INVX1 U6967 (.I(N11481), .ZN(N19839));
    INVX1 U6968 (.I(N11482), .ZN(n19840));
    INVX1 U6969 (.I(N11483), .ZN(n19841));
    INVX1 U6970 (.I(N11484), .ZN(n19842));
    INVX1 U6971 (.I(N11485), .ZN(n19843));
    INVX1 U6972 (.I(N11486), .ZN(N19844));
    INVX1 U6973 (.I(N11487), .ZN(n19845));
    INVX1 U6974 (.I(N11488), .ZN(n19846));
    INVX1 U6975 (.I(N11489), .ZN(n19847));
    INVX1 U6976 (.I(N11490), .ZN(n19848));
    INVX1 U6977 (.I(N11491), .ZN(n19849));
    INVX1 U6978 (.I(N11492), .ZN(n19850));
    INVX1 U6979 (.I(N11493), .ZN(N19851));
    INVX1 U6980 (.I(N11494), .ZN(N19852));
    INVX1 U6981 (.I(N11495), .ZN(n19853));
    INVX1 U6982 (.I(N11496), .ZN(n19854));
    INVX1 U6983 (.I(N11497), .ZN(n19855));
    INVX1 U6984 (.I(N11498), .ZN(n19856));
    INVX1 U6985 (.I(N11499), .ZN(n19857));
    INVX1 U6986 (.I(N11500), .ZN(n19858));
    INVX1 U6987 (.I(N11501), .ZN(N19859));
    INVX1 U6988 (.I(N11502), .ZN(n19860));
    INVX1 U6989 (.I(N11503), .ZN(n19861));
    INVX1 U6990 (.I(N11504), .ZN(n19862));
    INVX1 U6991 (.I(N11505), .ZN(n19863));
    INVX1 U6992 (.I(N11506), .ZN(N19864));
    INVX1 U6993 (.I(N11507), .ZN(n19865));
    INVX1 U6994 (.I(N11508), .ZN(n19866));
    INVX1 U6995 (.I(N11509), .ZN(n19867));
    INVX1 U6996 (.I(N11510), .ZN(n19868));
    INVX1 U6997 (.I(N11511), .ZN(n19869));
    INVX1 U6998 (.I(N11512), .ZN(N19870));
    INVX1 U6999 (.I(N11513), .ZN(N19871));
    INVX1 U7000 (.I(N11514), .ZN(N19872));
    INVX1 U7001 (.I(N11515), .ZN(n19873));
    INVX1 U7002 (.I(N11516), .ZN(n19874));
    INVX1 U7003 (.I(N11517), .ZN(n19875));
    INVX1 U7004 (.I(N11518), .ZN(n19876));
    INVX1 U7005 (.I(N11519), .ZN(n19877));
    INVX1 U7006 (.I(N11520), .ZN(n19878));
    INVX1 U7007 (.I(N11521), .ZN(n19879));
    INVX1 U7008 (.I(N11522), .ZN(n19880));
    INVX1 U7009 (.I(N11523), .ZN(N19881));
    INVX1 U7010 (.I(N11524), .ZN(n19882));
    INVX1 U7011 (.I(N11525), .ZN(n19883));
    INVX1 U7012 (.I(N11526), .ZN(n19884));
    INVX1 U7013 (.I(N11527), .ZN(n19885));
    INVX1 U7014 (.I(N11528), .ZN(n19886));
    INVX1 U7015 (.I(N11529), .ZN(n19887));
    INVX1 U7016 (.I(N11530), .ZN(n19888));
    INVX1 U7017 (.I(N11531), .ZN(n19889));
    INVX1 U7018 (.I(N11532), .ZN(n19890));
    INVX1 U7019 (.I(N11533), .ZN(n19891));
    INVX1 U7020 (.I(N11534), .ZN(N19892));
    INVX1 U7021 (.I(N11535), .ZN(N19893));
    INVX1 U7022 (.I(N11536), .ZN(n19894));
    INVX1 U7023 (.I(N11537), .ZN(n19895));
    INVX1 U7024 (.I(N11538), .ZN(n19896));
    INVX1 U7025 (.I(N11539), .ZN(N19897));
    INVX1 U7026 (.I(N11540), .ZN(n19898));
    INVX1 U7027 (.I(N11541), .ZN(n19899));
    INVX1 U7028 (.I(N11542), .ZN(n19900));
    INVX1 U7029 (.I(N11543), .ZN(n19901));
    INVX1 U7030 (.I(N11544), .ZN(n19902));
    INVX1 U7031 (.I(N11545), .ZN(n19903));
    INVX1 U7032 (.I(N11546), .ZN(n19904));
    INVX1 U7033 (.I(N11547), .ZN(N19905));
    INVX1 U7034 (.I(N11548), .ZN(n19906));
    INVX1 U7035 (.I(N11549), .ZN(n19907));
    INVX1 U7036 (.I(N11550), .ZN(n19908));
    INVX1 U7037 (.I(N11551), .ZN(N19909));
    INVX1 U7038 (.I(N11552), .ZN(n19910));
    INVX1 U7039 (.I(N11553), .ZN(n19911));
    INVX1 U7040 (.I(N11554), .ZN(n19912));
    INVX1 U7041 (.I(N11555), .ZN(n19913));
    INVX1 U7042 (.I(N11556), .ZN(n19914));
    INVX1 U7043 (.I(N11557), .ZN(n19915));
    INVX1 U7044 (.I(N11558), .ZN(n19916));
    INVX1 U7045 (.I(N11559), .ZN(n19917));
    INVX1 U7046 (.I(N11560), .ZN(N19918));
    INVX1 U7047 (.I(N11561), .ZN(n19919));
    INVX1 U7048 (.I(N11562), .ZN(N19920));
    INVX1 U7049 (.I(N11563), .ZN(N19921));
    INVX1 U7050 (.I(N11564), .ZN(n19922));
    INVX1 U7051 (.I(N11565), .ZN(n19923));
    INVX1 U7052 (.I(N11566), .ZN(n19924));
    INVX1 U7053 (.I(N11567), .ZN(n19925));
    INVX1 U7054 (.I(N11568), .ZN(n19926));
    INVX1 U7055 (.I(N11569), .ZN(N19927));
    INVX1 U7056 (.I(N11570), .ZN(n19928));
    INVX1 U7057 (.I(N11571), .ZN(n19929));
    INVX1 U7058 (.I(N11572), .ZN(n19930));
    INVX1 U7059 (.I(N11573), .ZN(n19931));
    INVX1 U7060 (.I(N11574), .ZN(n19932));
    INVX1 U7061 (.I(N11575), .ZN(n19933));
    INVX1 U7062 (.I(N11576), .ZN(n19934));
    INVX1 U7063 (.I(N11577), .ZN(n19935));
    INVX1 U7064 (.I(N11578), .ZN(n19936));
    INVX1 U7065 (.I(N11579), .ZN(N19937));
    INVX1 U7066 (.I(N11580), .ZN(N19938));
    INVX1 U7067 (.I(N11581), .ZN(N19939));
    INVX1 U7068 (.I(N11582), .ZN(n19940));
    INVX1 U7069 (.I(N11583), .ZN(n19941));
    INVX1 U7070 (.I(N11584), .ZN(N19942));
    INVX1 U7071 (.I(N11585), .ZN(n19943));
    INVX1 U7072 (.I(N11586), .ZN(n19944));
    INVX1 U7073 (.I(N11587), .ZN(n19945));
    INVX1 U7074 (.I(N11588), .ZN(n19946));
    INVX1 U7075 (.I(N11589), .ZN(n19947));
    INVX1 U7076 (.I(N11590), .ZN(N19948));
    INVX1 U7077 (.I(N11591), .ZN(n19949));
    INVX1 U7078 (.I(N11592), .ZN(n19950));
    INVX1 U7079 (.I(N11593), .ZN(N19951));
    INVX1 U7080 (.I(N11594), .ZN(n19952));
    INVX1 U7081 (.I(N11595), .ZN(N19953));
    INVX1 U7082 (.I(N11596), .ZN(n19954));
    INVX1 U7083 (.I(N11597), .ZN(n19955));
    INVX1 U7084 (.I(N11598), .ZN(n19956));
    INVX1 U7085 (.I(N11599), .ZN(n19957));
    INVX1 U7086 (.I(N11600), .ZN(n19958));
    INVX1 U7087 (.I(N11601), .ZN(n19959));
    INVX1 U7088 (.I(N11602), .ZN(N19960));
    INVX1 U7089 (.I(N11603), .ZN(n19961));
    INVX1 U7090 (.I(N11604), .ZN(n19962));
    INVX1 U7091 (.I(N11605), .ZN(n19963));
    INVX1 U7092 (.I(N11606), .ZN(n19964));
    INVX1 U7093 (.I(N11607), .ZN(n19965));
    INVX1 U7094 (.I(N11608), .ZN(n19966));
    INVX1 U7095 (.I(N11609), .ZN(n19967));
    INVX1 U7096 (.I(N11610), .ZN(N19968));
    INVX1 U7097 (.I(N11611), .ZN(N19969));
    INVX1 U7098 (.I(N11612), .ZN(n19970));
    INVX1 U7099 (.I(N11613), .ZN(n19971));
    INVX1 U7100 (.I(N11614), .ZN(n19972));
    INVX1 U7101 (.I(N11615), .ZN(n19973));
    INVX1 U7102 (.I(N11616), .ZN(n19974));
    INVX1 U7103 (.I(N11617), .ZN(n19975));
    INVX1 U7104 (.I(N11618), .ZN(n19976));
    INVX1 U7105 (.I(N11619), .ZN(n19977));
    INVX1 U7106 (.I(N11620), .ZN(N19978));
    INVX1 U7107 (.I(N11621), .ZN(n19979));
    INVX1 U7108 (.I(N11622), .ZN(n19980));
    INVX1 U7109 (.I(N11623), .ZN(n19981));
    INVX1 U7110 (.I(N11624), .ZN(n19982));
    INVX1 U7111 (.I(N11625), .ZN(n19983));
    INVX1 U7112 (.I(N11626), .ZN(n19984));
    INVX1 U7113 (.I(N11627), .ZN(n19985));
    INVX1 U7114 (.I(N11628), .ZN(N19986));
    INVX1 U7115 (.I(N11629), .ZN(n19987));
    INVX1 U7116 (.I(N11630), .ZN(N19988));
    INVX1 U7117 (.I(N11631), .ZN(n19989));
    INVX1 U7118 (.I(N11632), .ZN(n19990));
    INVX1 U7119 (.I(N11633), .ZN(n19991));
    INVX1 U7120 (.I(N11634), .ZN(n19992));
    INVX1 U7121 (.I(N11635), .ZN(n19993));
    INVX1 U7122 (.I(N11636), .ZN(n19994));
    INVX1 U7123 (.I(N11637), .ZN(N19995));
    INVX1 U7124 (.I(N11638), .ZN(n19996));
    INVX1 U7125 (.I(N11639), .ZN(n19997));
    INVX1 U7126 (.I(N11640), .ZN(N19998));
    INVX1 U7127 (.I(N11641), .ZN(n19999));
    INVX1 U7128 (.I(N11642), .ZN(n20000));
    INVX1 U7129 (.I(N11643), .ZN(n20001));
    INVX1 U7130 (.I(N11644), .ZN(N20002));
    INVX1 U7131 (.I(N11645), .ZN(N20003));
    INVX1 U7132 (.I(N11646), .ZN(n20004));
    INVX1 U7133 (.I(N11647), .ZN(n20005));
    INVX1 U7134 (.I(N11648), .ZN(n20006));
    INVX1 U7135 (.I(N11649), .ZN(N20007));
    INVX1 U7136 (.I(N11650), .ZN(n20008));
    INVX1 U7137 (.I(N11651), .ZN(n20009));
    INVX1 U7138 (.I(N11652), .ZN(N20010));
    INVX1 U7139 (.I(N11653), .ZN(n20011));
    INVX1 U7140 (.I(N11654), .ZN(n20012));
    INVX1 U7141 (.I(N11655), .ZN(n20013));
    INVX1 U7142 (.I(N11656), .ZN(n20014));
    INVX1 U7143 (.I(N11657), .ZN(n20015));
    INVX1 U7144 (.I(N11658), .ZN(n20016));
    INVX1 U7145 (.I(N11659), .ZN(n20017));
    INVX1 U7146 (.I(N11660), .ZN(N20018));
    INVX1 U7147 (.I(N11661), .ZN(N20019));
    INVX1 U7148 (.I(N11662), .ZN(n20020));
    INVX1 U7149 (.I(N11663), .ZN(n20021));
    INVX1 U7150 (.I(N11664), .ZN(n20022));
    INVX1 U7151 (.I(N11665), .ZN(n20023));
    INVX1 U7152 (.I(N11666), .ZN(n20024));
    INVX1 U7153 (.I(N11667), .ZN(n20025));
    INVX1 U7154 (.I(N11668), .ZN(n20026));
    INVX1 U7155 (.I(N11669), .ZN(n20027));
    INVX1 U7156 (.I(N11670), .ZN(n20028));
    INVX1 U7157 (.I(N11671), .ZN(n20029));
    INVX1 U7158 (.I(N11672), .ZN(n20030));
    INVX1 U7159 (.I(N11673), .ZN(n20031));
    INVX1 U7160 (.I(N11674), .ZN(n20032));
    INVX1 U7161 (.I(N11675), .ZN(n20033));
    INVX1 U7162 (.I(N11676), .ZN(n20034));
    INVX1 U7163 (.I(N11677), .ZN(n20035));
    INVX1 U7164 (.I(N11678), .ZN(N20036));
    INVX1 U7165 (.I(N11679), .ZN(n20037));
    INVX1 U7166 (.I(N11680), .ZN(n20038));
    INVX1 U7167 (.I(N11681), .ZN(n20039));
    INVX1 U7168 (.I(N11682), .ZN(n20040));
    INVX1 U7169 (.I(N11683), .ZN(n20041));
    INVX1 U7170 (.I(N11684), .ZN(N20042));
    INVX1 U7171 (.I(N11685), .ZN(n20043));
    INVX1 U7172 (.I(N11686), .ZN(n20044));
    INVX1 U7173 (.I(N11687), .ZN(n20045));
    INVX1 U7174 (.I(N11688), .ZN(n20046));
    INVX1 U7175 (.I(N11689), .ZN(N20047));
    INVX1 U7176 (.I(N11690), .ZN(N20048));
    INVX1 U7177 (.I(N11691), .ZN(n20049));
    INVX1 U7178 (.I(N11692), .ZN(n20050));
    INVX1 U7179 (.I(N11693), .ZN(n20051));
    INVX1 U7180 (.I(N11694), .ZN(n20052));
    INVX1 U7181 (.I(N11695), .ZN(n20053));
    INVX1 U7182 (.I(N11696), .ZN(n20054));
    INVX1 U7183 (.I(N11697), .ZN(N20055));
    INVX1 U7184 (.I(N11698), .ZN(n20056));
    INVX1 U7185 (.I(N11699), .ZN(N20057));
    INVX1 U7186 (.I(N11700), .ZN(n20058));
    INVX1 U7187 (.I(N11701), .ZN(N20059));
    INVX1 U7188 (.I(N11702), .ZN(N20060));
    INVX1 U7189 (.I(N11703), .ZN(n20061));
    INVX1 U7190 (.I(N11704), .ZN(n20062));
    INVX1 U7191 (.I(N11705), .ZN(n20063));
    INVX1 U7192 (.I(N11706), .ZN(n20064));
    INVX1 U7193 (.I(N11707), .ZN(n20065));
    INVX1 U7194 (.I(N11708), .ZN(N20066));
    INVX1 U7195 (.I(N11709), .ZN(n20067));
    INVX1 U7196 (.I(N11710), .ZN(N20068));
    INVX1 U7197 (.I(N11711), .ZN(N20069));
    INVX1 U7198 (.I(N11712), .ZN(n20070));
    INVX1 U7199 (.I(N11713), .ZN(n20071));
    INVX1 U7200 (.I(N11714), .ZN(N20072));
    INVX1 U7201 (.I(N11715), .ZN(n20073));
    INVX1 U7202 (.I(N11716), .ZN(N20074));
    INVX1 U7203 (.I(N11717), .ZN(n20075));
    INVX1 U7204 (.I(N11718), .ZN(n20076));
    INVX1 U7205 (.I(N11719), .ZN(N20077));
    INVX1 U7206 (.I(N11720), .ZN(n20078));
    INVX1 U7207 (.I(N11721), .ZN(n20079));
    INVX1 U7208 (.I(N11722), .ZN(n20080));
    INVX1 U7209 (.I(N11723), .ZN(n20081));
    INVX1 U7210 (.I(N11724), .ZN(N20082));
    INVX1 U7211 (.I(N11725), .ZN(n20083));
    INVX1 U7212 (.I(N11726), .ZN(n20084));
    INVX1 U7213 (.I(N11727), .ZN(n20085));
    INVX1 U7214 (.I(N11728), .ZN(n20086));
    INVX1 U7215 (.I(N11729), .ZN(N20087));
    INVX1 U7216 (.I(N11730), .ZN(n20088));
    INVX1 U7217 (.I(N11731), .ZN(N20089));
    INVX1 U7218 (.I(N11732), .ZN(n20090));
    INVX1 U7219 (.I(N11733), .ZN(n20091));
    INVX1 U7220 (.I(N11734), .ZN(n20092));
    INVX1 U7221 (.I(N11735), .ZN(n20093));
    INVX1 U7222 (.I(N11736), .ZN(n20094));
    INVX1 U7223 (.I(N11737), .ZN(n20095));
    INVX1 U7224 (.I(N11738), .ZN(n20096));
    INVX1 U7225 (.I(N11739), .ZN(n20097));
    INVX1 U7226 (.I(N11740), .ZN(n20098));
    INVX1 U7227 (.I(N11741), .ZN(N20099));
    INVX1 U7228 (.I(N11742), .ZN(n20100));
    INVX1 U7229 (.I(N11743), .ZN(n20101));
    INVX1 U7230 (.I(N11744), .ZN(n20102));
    INVX1 U7231 (.I(N11745), .ZN(n20103));
    INVX1 U7232 (.I(N11746), .ZN(n20104));
    INVX1 U7233 (.I(N11747), .ZN(N20105));
    INVX1 U7234 (.I(N11748), .ZN(n20106));
    INVX1 U7235 (.I(N11749), .ZN(n20107));
    INVX1 U7236 (.I(N11750), .ZN(N20108));
    INVX1 U7237 (.I(N11751), .ZN(n20109));
    INVX1 U7238 (.I(N11752), .ZN(n20110));
    INVX1 U7239 (.I(N11753), .ZN(n20111));
    INVX1 U7240 (.I(N11754), .ZN(n20112));
    INVX1 U7241 (.I(N11755), .ZN(n20113));
    INVX1 U7242 (.I(N11756), .ZN(n20114));
    INVX1 U7243 (.I(N11757), .ZN(n20115));
    INVX1 U7244 (.I(N11758), .ZN(n20116));
    INVX1 U7245 (.I(N11759), .ZN(n20117));
    INVX1 U7246 (.I(N11760), .ZN(n20118));
    INVX1 U7247 (.I(N11761), .ZN(N20119));
    INVX1 U7248 (.I(N11762), .ZN(n20120));
    INVX1 U7249 (.I(N11763), .ZN(n20121));
    INVX1 U7250 (.I(N11764), .ZN(n20122));
    INVX1 U7251 (.I(N11765), .ZN(N20123));
    INVX1 U7252 (.I(N11766), .ZN(n20124));
    INVX1 U7253 (.I(N11767), .ZN(N20125));
    INVX1 U7254 (.I(N11768), .ZN(n20126));
    INVX1 U7255 (.I(N11769), .ZN(n20127));
    INVX1 U7256 (.I(N11770), .ZN(n20128));
    INVX1 U7257 (.I(N11771), .ZN(n20129));
    INVX1 U7258 (.I(N11772), .ZN(n20130));
    INVX1 U7259 (.I(N11773), .ZN(n20131));
    INVX1 U7260 (.I(N11774), .ZN(n20132));
    INVX1 U7261 (.I(N11775), .ZN(n20133));
    INVX1 U7262 (.I(N11776), .ZN(n20134));
    INVX1 U7263 (.I(N11777), .ZN(N20135));
    INVX1 U7264 (.I(N11778), .ZN(n20136));
    INVX1 U7265 (.I(N11779), .ZN(n20137));
    INVX1 U7266 (.I(N11780), .ZN(N20138));
    INVX1 U7267 (.I(N11781), .ZN(n20139));
    INVX1 U7268 (.I(N11782), .ZN(n20140));
    INVX1 U7269 (.I(N11783), .ZN(n20141));
    INVX1 U7270 (.I(N11784), .ZN(n20142));
    INVX1 U7271 (.I(N11785), .ZN(n20143));
    INVX1 U7272 (.I(N11786), .ZN(n20144));
    INVX1 U7273 (.I(N11787), .ZN(n20145));
    INVX1 U7274 (.I(N11788), .ZN(N20146));
    INVX1 U7275 (.I(N11789), .ZN(n20147));
    INVX1 U7276 (.I(N11790), .ZN(n20148));
    INVX1 U7277 (.I(N11791), .ZN(n20149));
    INVX1 U7278 (.I(N11792), .ZN(n20150));
    INVX1 U7279 (.I(N11793), .ZN(n20151));
    INVX1 U7280 (.I(N11794), .ZN(n20152));
    INVX1 U7281 (.I(N11795), .ZN(n20153));
    INVX1 U7282 (.I(N11796), .ZN(N20154));
    INVX1 U7283 (.I(N11797), .ZN(n20155));
    INVX1 U7284 (.I(N11798), .ZN(n20156));
    INVX1 U7285 (.I(N11799), .ZN(n20157));
    INVX1 U7286 (.I(N11800), .ZN(N20158));
    INVX1 U7287 (.I(N11801), .ZN(n20159));
    INVX1 U7288 (.I(N11802), .ZN(n20160));
    INVX1 U7289 (.I(N11803), .ZN(n20161));
    INVX1 U7290 (.I(N11804), .ZN(n20162));
    INVX1 U7291 (.I(N11805), .ZN(n20163));
    INVX1 U7292 (.I(N11806), .ZN(N20164));
    INVX1 U7293 (.I(N11807), .ZN(n20165));
    INVX1 U7294 (.I(N11808), .ZN(n20166));
    INVX1 U7295 (.I(N11809), .ZN(n20167));
    INVX1 U7296 (.I(N11810), .ZN(n20168));
    INVX1 U7297 (.I(N11811), .ZN(n20169));
    INVX1 U7298 (.I(N11812), .ZN(n20170));
    INVX1 U7299 (.I(N11813), .ZN(n20171));
    INVX1 U7300 (.I(N11814), .ZN(n20172));
    INVX1 U7301 (.I(N11815), .ZN(n20173));
    INVX1 U7302 (.I(N11816), .ZN(n20174));
    INVX1 U7303 (.I(N11817), .ZN(n20175));
    INVX1 U7304 (.I(N11818), .ZN(n20176));
    INVX1 U7305 (.I(N11819), .ZN(n20177));
    INVX1 U7306 (.I(N11820), .ZN(n20178));
    INVX1 U7307 (.I(N11821), .ZN(n20179));
    INVX1 U7308 (.I(N11822), .ZN(n20180));
    INVX1 U7309 (.I(N11823), .ZN(n20181));
    INVX1 U7310 (.I(N11824), .ZN(n20182));
    INVX1 U7311 (.I(N11825), .ZN(n20183));
    INVX1 U7312 (.I(N11826), .ZN(n20184));
    INVX1 U7313 (.I(N11827), .ZN(n20185));
    INVX1 U7314 (.I(N11828), .ZN(N20186));
    INVX1 U7315 (.I(N11829), .ZN(n20187));
    INVX1 U7316 (.I(N11830), .ZN(n20188));
    INVX1 U7317 (.I(N11831), .ZN(N20189));
    INVX1 U7318 (.I(N11832), .ZN(N20190));
    INVX1 U7319 (.I(N11833), .ZN(N20191));
    INVX1 U7320 (.I(N11834), .ZN(N20192));
    INVX1 U7321 (.I(N11835), .ZN(n20193));
    INVX1 U7322 (.I(N11836), .ZN(n20194));
    INVX1 U7323 (.I(N11837), .ZN(n20195));
    INVX1 U7324 (.I(N11838), .ZN(n20196));
    INVX1 U7325 (.I(N11839), .ZN(N20197));
    INVX1 U7326 (.I(N11840), .ZN(n20198));
    INVX1 U7327 (.I(N11841), .ZN(N20199));
    INVX1 U7328 (.I(N11842), .ZN(n20200));
    INVX1 U7329 (.I(N11843), .ZN(n20201));
    INVX1 U7330 (.I(N11844), .ZN(n20202));
    INVX1 U7331 (.I(N11845), .ZN(N20203));
    INVX1 U7332 (.I(N11846), .ZN(n20204));
    INVX1 U7333 (.I(N11847), .ZN(n20205));
    INVX1 U7334 (.I(N11848), .ZN(n20206));
    INVX1 U7335 (.I(N11849), .ZN(n20207));
    INVX1 U7336 (.I(N11850), .ZN(N20208));
    INVX1 U7337 (.I(N11851), .ZN(n20209));
    INVX1 U7338 (.I(N11852), .ZN(n20210));
    INVX1 U7339 (.I(N11853), .ZN(n20211));
    INVX1 U7340 (.I(N11854), .ZN(n20212));
    INVX1 U7341 (.I(N11855), .ZN(n20213));
    INVX1 U7342 (.I(N11856), .ZN(n20214));
    INVX1 U7343 (.I(N11857), .ZN(n20215));
    INVX1 U7344 (.I(N11858), .ZN(n20216));
    INVX1 U7345 (.I(N11859), .ZN(N20217));
    INVX1 U7346 (.I(N11860), .ZN(N20218));
    INVX1 U7347 (.I(N11861), .ZN(n20219));
    INVX1 U7348 (.I(N11862), .ZN(n20220));
    INVX1 U7349 (.I(N11863), .ZN(n20221));
    INVX1 U7350 (.I(N11864), .ZN(n20222));
    INVX1 U7351 (.I(N11865), .ZN(n20223));
    INVX1 U7352 (.I(N11866), .ZN(n20224));
    INVX1 U7353 (.I(N11867), .ZN(n20225));
    INVX1 U7354 (.I(N11868), .ZN(n20226));
    INVX1 U7355 (.I(N11869), .ZN(N20227));
    INVX1 U7356 (.I(N11870), .ZN(n20228));
    INVX1 U7357 (.I(N11871), .ZN(n20229));
    INVX1 U7358 (.I(N11872), .ZN(n20230));
    INVX1 U7359 (.I(N11873), .ZN(n20231));
    INVX1 U7360 (.I(N11874), .ZN(n20232));
    INVX1 U7361 (.I(N11875), .ZN(n20233));
    INVX1 U7362 (.I(N11876), .ZN(n20234));
    INVX1 U7363 (.I(N11877), .ZN(n20235));
    INVX1 U7364 (.I(N11878), .ZN(n20236));
    INVX1 U7365 (.I(N11879), .ZN(n20237));
    INVX1 U7366 (.I(N11880), .ZN(n20238));
    INVX1 U7367 (.I(N11881), .ZN(n20239));
    INVX1 U7368 (.I(N11882), .ZN(n20240));
    INVX1 U7369 (.I(N11883), .ZN(n20241));
    INVX1 U7370 (.I(N11884), .ZN(n20242));
    INVX1 U7371 (.I(N11885), .ZN(n20243));
    INVX1 U7372 (.I(N11886), .ZN(n20244));
    INVX1 U7373 (.I(N11887), .ZN(n20245));
    INVX1 U7374 (.I(N11888), .ZN(n20246));
    INVX1 U7375 (.I(N11889), .ZN(n20247));
    INVX1 U7376 (.I(N11890), .ZN(n20248));
    INVX1 U7377 (.I(N11891), .ZN(N20249));
    INVX1 U7378 (.I(N11892), .ZN(n20250));
    INVX1 U7379 (.I(N11893), .ZN(n20251));
    INVX1 U7380 (.I(N11894), .ZN(n20252));
    INVX1 U7381 (.I(N11895), .ZN(n20253));
    INVX1 U7382 (.I(N11896), .ZN(n20254));
    INVX1 U7383 (.I(N11897), .ZN(n20255));
    INVX1 U7384 (.I(N11898), .ZN(n20256));
    INVX1 U7385 (.I(N11899), .ZN(n20257));
    INVX1 U7386 (.I(N11900), .ZN(n20258));
    INVX1 U7387 (.I(N11901), .ZN(n20259));
    INVX1 U7388 (.I(N11902), .ZN(n20260));
    INVX1 U7389 (.I(N11903), .ZN(n20261));
    INVX1 U7390 (.I(N11904), .ZN(n20262));
    INVX1 U7391 (.I(N11905), .ZN(n20263));
    INVX1 U7392 (.I(N11906), .ZN(n20264));
    INVX1 U7393 (.I(N11907), .ZN(n20265));
    INVX1 U7394 (.I(N11908), .ZN(n20266));
    INVX1 U7395 (.I(N11909), .ZN(n20267));
    INVX1 U7396 (.I(N11910), .ZN(n20268));
    INVX1 U7397 (.I(N11911), .ZN(n20269));
    INVX1 U7398 (.I(N11912), .ZN(N20270));
    INVX1 U7399 (.I(N11913), .ZN(n20271));
    INVX1 U7400 (.I(N11914), .ZN(n20272));
    INVX1 U7401 (.I(N11915), .ZN(n20273));
    INVX1 U7402 (.I(N11916), .ZN(n20274));
    INVX1 U7403 (.I(N11917), .ZN(n20275));
    INVX1 U7404 (.I(N11918), .ZN(n20276));
    INVX1 U7405 (.I(N11919), .ZN(N20277));
    INVX1 U7406 (.I(N11920), .ZN(N20278));
    INVX1 U7407 (.I(N11921), .ZN(N20279));
    INVX1 U7408 (.I(N11922), .ZN(n20280));
    INVX1 U7409 (.I(N11923), .ZN(N20281));
    INVX1 U7410 (.I(N11924), .ZN(n20282));
    INVX1 U7411 (.I(N11925), .ZN(n20283));
    INVX1 U7412 (.I(N11926), .ZN(N20284));
    INVX1 U7413 (.I(N11927), .ZN(n20285));
    INVX1 U7414 (.I(N11928), .ZN(N20286));
    INVX1 U7415 (.I(N11929), .ZN(N20287));
    INVX1 U7416 (.I(N11930), .ZN(n20288));
    INVX1 U7417 (.I(N11931), .ZN(n20289));
    INVX1 U7418 (.I(N11932), .ZN(n20290));
    INVX1 U7419 (.I(N11933), .ZN(N20291));
    INVX1 U7420 (.I(N11934), .ZN(N20292));
    INVX1 U7421 (.I(N11935), .ZN(n20293));
    INVX1 U7422 (.I(N11936), .ZN(n20294));
    INVX1 U7423 (.I(N11937), .ZN(N20295));
    INVX1 U7424 (.I(N11938), .ZN(n20296));
    INVX1 U7425 (.I(N11939), .ZN(n20297));
    INVX1 U7426 (.I(N11940), .ZN(n20298));
    INVX1 U7427 (.I(N11941), .ZN(N20299));
    INVX1 U7428 (.I(N11942), .ZN(N20300));
    INVX1 U7429 (.I(N11943), .ZN(n20301));
    INVX1 U7430 (.I(N11944), .ZN(n20302));
    INVX1 U7431 (.I(N11945), .ZN(n20303));
    INVX1 U7432 (.I(N11946), .ZN(n20304));
    INVX1 U7433 (.I(N11947), .ZN(n20305));
    INVX1 U7434 (.I(N11948), .ZN(n20306));
    INVX1 U7435 (.I(N11949), .ZN(n20307));
    INVX1 U7436 (.I(N11950), .ZN(n20308));
    INVX1 U7437 (.I(N11951), .ZN(N20309));
    INVX1 U7438 (.I(N11952), .ZN(n20310));
    INVX1 U7439 (.I(N11953), .ZN(n20311));
    INVX1 U7440 (.I(N11954), .ZN(n20312));
    INVX1 U7441 (.I(N11955), .ZN(n20313));
    INVX1 U7442 (.I(N11956), .ZN(N20314));
    INVX1 U7443 (.I(N11957), .ZN(n20315));
    INVX1 U7444 (.I(N11958), .ZN(n20316));
    INVX1 U7445 (.I(N11959), .ZN(n20317));
    INVX1 U7446 (.I(N11960), .ZN(n20318));
    INVX1 U7447 (.I(N11961), .ZN(n20319));
    INVX1 U7448 (.I(N11962), .ZN(n20320));
    INVX1 U7449 (.I(N11963), .ZN(n20321));
    INVX1 U7450 (.I(N11964), .ZN(n20322));
    INVX1 U7451 (.I(N11965), .ZN(n20323));
    INVX1 U7452 (.I(N11966), .ZN(n20324));
    INVX1 U7453 (.I(N11967), .ZN(n20325));
    INVX1 U7454 (.I(N11968), .ZN(n20326));
    INVX1 U7455 (.I(N11969), .ZN(n20327));
    INVX1 U7456 (.I(N11970), .ZN(n20328));
    INVX1 U7457 (.I(N11971), .ZN(n20329));
    INVX1 U7458 (.I(N11972), .ZN(n20330));
    INVX1 U7459 (.I(N11973), .ZN(n20331));
    INVX1 U7460 (.I(N11974), .ZN(n20332));
    INVX1 U7461 (.I(N11975), .ZN(N20333));
    INVX1 U7462 (.I(N11976), .ZN(n20334));
    INVX1 U7463 (.I(N11977), .ZN(n20335));
    INVX1 U7464 (.I(N11978), .ZN(n20336));
    INVX1 U7465 (.I(N11979), .ZN(n20337));
    INVX1 U7466 (.I(N11980), .ZN(n20338));
    INVX1 U7467 (.I(N11981), .ZN(n20339));
    INVX1 U7468 (.I(N11982), .ZN(n20340));
    INVX1 U7469 (.I(N11983), .ZN(n20341));
    INVX1 U7470 (.I(N11984), .ZN(n20342));
    INVX1 U7471 (.I(N11985), .ZN(n20343));
    INVX1 U7472 (.I(N11986), .ZN(n20344));
    INVX1 U7473 (.I(N11987), .ZN(N20345));
    INVX1 U7474 (.I(N11988), .ZN(n20346));
    INVX1 U7475 (.I(N11989), .ZN(n20347));
    INVX1 U7476 (.I(N11990), .ZN(n20348));
    INVX1 U7477 (.I(N11991), .ZN(n20349));
    INVX1 U7478 (.I(N11992), .ZN(n20350));
    INVX1 U7479 (.I(N11993), .ZN(n20351));
    INVX1 U7480 (.I(N11994), .ZN(n20352));
    INVX1 U7481 (.I(N11995), .ZN(n20353));
    INVX1 U7482 (.I(N11996), .ZN(N20354));
    INVX1 U7483 (.I(N11997), .ZN(n20355));
    INVX1 U7484 (.I(N11998), .ZN(n20356));
    INVX1 U7485 (.I(N11999), .ZN(n20357));
    INVX1 U7486 (.I(N12000), .ZN(n20358));
    INVX1 U7487 (.I(N12001), .ZN(N20359));
    INVX1 U7488 (.I(N12002), .ZN(N20360));
    INVX1 U7489 (.I(N12003), .ZN(n20361));
    INVX1 U7490 (.I(N12004), .ZN(n20362));
    INVX1 U7491 (.I(N12005), .ZN(n20363));
    INVX1 U7492 (.I(N12006), .ZN(n20364));
    INVX1 U7493 (.I(N12007), .ZN(n20365));
    INVX1 U7494 (.I(N12008), .ZN(n20366));
    INVX1 U7495 (.I(N12009), .ZN(N20367));
    INVX1 U7496 (.I(N12010), .ZN(n20368));
    INVX1 U7497 (.I(N12011), .ZN(N20369));
    INVX1 U7498 (.I(N12012), .ZN(n20370));
    INVX1 U7499 (.I(N12013), .ZN(n20371));
    INVX1 U7500 (.I(N12014), .ZN(n20372));
    INVX1 U7501 (.I(N12015), .ZN(n20373));
    INVX1 U7502 (.I(N12016), .ZN(n20374));
    INVX1 U7503 (.I(N12017), .ZN(n20375));
    INVX1 U7504 (.I(N12018), .ZN(N20376));
    INVX1 U7505 (.I(N12019), .ZN(n20377));
    INVX1 U7506 (.I(N12020), .ZN(n20378));
    INVX1 U7507 (.I(N12021), .ZN(n20379));
    INVX1 U7508 (.I(N12022), .ZN(n20380));
    INVX1 U7509 (.I(N12023), .ZN(n20381));
    INVX1 U7510 (.I(N12024), .ZN(n20382));
    INVX1 U7511 (.I(N12025), .ZN(n20383));
    INVX1 U7512 (.I(N12026), .ZN(n20384));
    INVX1 U7513 (.I(N12027), .ZN(n20385));
    INVX1 U7514 (.I(N12028), .ZN(n20386));
    INVX1 U7515 (.I(N12029), .ZN(n20387));
    INVX1 U7516 (.I(N12030), .ZN(n20388));
    INVX1 U7517 (.I(N12031), .ZN(n20389));
    INVX1 U7518 (.I(N12032), .ZN(n20390));
    INVX1 U7519 (.I(N12033), .ZN(n20391));
    INVX1 U7520 (.I(N12034), .ZN(n20392));
    INVX1 U7521 (.I(N12035), .ZN(n20393));
    INVX1 U7522 (.I(N12036), .ZN(N20394));
    INVX1 U7523 (.I(N12037), .ZN(n20395));
    INVX1 U7524 (.I(N12038), .ZN(N20396));
    INVX1 U7525 (.I(N12039), .ZN(n20397));
    INVX1 U7526 (.I(N12040), .ZN(n20398));
    INVX1 U7527 (.I(N12041), .ZN(n20399));
    INVX1 U7528 (.I(N12042), .ZN(n20400));
    INVX1 U7529 (.I(N12043), .ZN(n20401));
    INVX1 U7530 (.I(N12044), .ZN(n20402));
    INVX1 U7531 (.I(N12045), .ZN(N20403));
    INVX1 U7532 (.I(N12046), .ZN(N20404));
    INVX1 U7533 (.I(N12047), .ZN(n20405));
    INVX1 U7534 (.I(N12048), .ZN(n20406));
    INVX1 U7535 (.I(N12049), .ZN(N20407));
    INVX1 U7536 (.I(N12050), .ZN(N20408));
    INVX1 U7537 (.I(N12051), .ZN(N20409));
    INVX1 U7538 (.I(N12052), .ZN(n20410));
    INVX1 U7539 (.I(N12053), .ZN(N20411));
    INVX1 U7540 (.I(N12054), .ZN(n20412));
    INVX1 U7541 (.I(N12055), .ZN(N20413));
    INVX1 U7542 (.I(N12056), .ZN(n20414));
    INVX1 U7543 (.I(N12057), .ZN(n20415));
    INVX1 U7544 (.I(N12058), .ZN(n20416));
    INVX1 U7545 (.I(N12059), .ZN(n20417));
    INVX1 U7546 (.I(N12060), .ZN(n20418));
    INVX1 U7547 (.I(N12061), .ZN(n20419));
    INVX1 U7548 (.I(N12062), .ZN(n20420));
    INVX1 U7549 (.I(N12063), .ZN(n20421));
    INVX1 U7550 (.I(N12064), .ZN(N20422));
    INVX1 U7551 (.I(N12065), .ZN(n20423));
    INVX1 U7552 (.I(N12066), .ZN(n20424));
    INVX1 U7553 (.I(N12067), .ZN(N20425));
    INVX1 U7554 (.I(N12068), .ZN(n20426));
    INVX1 U7555 (.I(N12069), .ZN(n20427));
    INVX1 U7556 (.I(N12070), .ZN(n20428));
    INVX1 U7557 (.I(N12071), .ZN(N20429));
    INVX1 U7558 (.I(N12072), .ZN(n20430));
    INVX1 U7559 (.I(N12073), .ZN(n20431));
    INVX1 U7560 (.I(N12074), .ZN(n20432));
    INVX1 U7561 (.I(N12075), .ZN(n20433));
    INVX1 U7562 (.I(N12076), .ZN(n20434));
    INVX1 U7563 (.I(N12077), .ZN(n20435));
    INVX1 U7564 (.I(N12078), .ZN(n20436));
    INVX1 U7565 (.I(N12079), .ZN(n20437));
    INVX1 U7566 (.I(N12080), .ZN(n20438));
    INVX1 U7567 (.I(N12081), .ZN(n20439));
    INVX1 U7568 (.I(N12082), .ZN(n20440));
    INVX1 U7569 (.I(N12083), .ZN(n20441));
    INVX1 U7570 (.I(N12084), .ZN(n20442));
    INVX1 U7571 (.I(N12085), .ZN(n20443));
    INVX1 U7572 (.I(N12086), .ZN(n20444));
    INVX1 U7573 (.I(N12087), .ZN(N20445));
    INVX1 U7574 (.I(N12088), .ZN(n20446));
    INVX1 U7575 (.I(N12089), .ZN(n20447));
    INVX1 U7576 (.I(N12090), .ZN(n20448));
    INVX1 U7577 (.I(N12091), .ZN(n20449));
    INVX1 U7578 (.I(N12092), .ZN(n20450));
    INVX1 U7579 (.I(N12093), .ZN(n20451));
    INVX1 U7580 (.I(N12094), .ZN(n20452));
    INVX1 U7581 (.I(N12095), .ZN(n20453));
    INVX1 U7582 (.I(N12096), .ZN(n20454));
    INVX1 U7583 (.I(N12097), .ZN(N20455));
    INVX1 U7584 (.I(N12098), .ZN(n20456));
    INVX1 U7585 (.I(N12099), .ZN(n20457));
    INVX1 U7586 (.I(N12100), .ZN(N20458));
    INVX1 U7587 (.I(N12101), .ZN(n20459));
    INVX1 U7588 (.I(N12102), .ZN(n20460));
    INVX1 U7589 (.I(N12103), .ZN(n20461));
    INVX1 U7590 (.I(N12104), .ZN(n20462));
    INVX1 U7591 (.I(N12105), .ZN(n20463));
    INVX1 U7592 (.I(N12106), .ZN(n20464));
    INVX1 U7593 (.I(N12107), .ZN(n20465));
    INVX1 U7594 (.I(N12108), .ZN(n20466));
    INVX1 U7595 (.I(N12109), .ZN(n20467));
    INVX1 U7596 (.I(N12110), .ZN(n20468));
    INVX1 U7597 (.I(N12111), .ZN(n20469));
    INVX1 U7598 (.I(N12112), .ZN(n20470));
    INVX1 U7599 (.I(N12113), .ZN(n20471));
    INVX1 U7600 (.I(N12114), .ZN(n20472));
    INVX1 U7601 (.I(N12115), .ZN(n20473));
    INVX1 U7602 (.I(N12116), .ZN(n20474));
    INVX1 U7603 (.I(N12117), .ZN(n20475));
    INVX1 U7604 (.I(N12118), .ZN(n20476));
    INVX1 U7605 (.I(N12119), .ZN(n20477));
    INVX1 U7606 (.I(N12120), .ZN(n20478));
    INVX1 U7607 (.I(N12121), .ZN(N20479));
    INVX1 U7608 (.I(N12122), .ZN(n20480));
    INVX1 U7609 (.I(N12123), .ZN(n20481));
    INVX1 U7610 (.I(N12124), .ZN(n20482));
    INVX1 U7611 (.I(N12125), .ZN(n20483));
    INVX1 U7612 (.I(N12126), .ZN(N20484));
    INVX1 U7613 (.I(N12127), .ZN(n20485));
    INVX1 U7614 (.I(N12128), .ZN(n20486));
    INVX1 U7615 (.I(N12129), .ZN(n20487));
    INVX1 U7616 (.I(N12130), .ZN(n20488));
    INVX1 U7617 (.I(N12131), .ZN(n20489));
    INVX1 U7618 (.I(N12132), .ZN(n20490));
    INVX1 U7619 (.I(N12133), .ZN(n20491));
    INVX1 U7620 (.I(N12134), .ZN(n20492));
    INVX1 U7621 (.I(N12135), .ZN(N20493));
    INVX1 U7622 (.I(N12136), .ZN(n20494));
    INVX1 U7623 (.I(N12137), .ZN(N20495));
    INVX1 U7624 (.I(N12138), .ZN(n20496));
    INVX1 U7625 (.I(N12139), .ZN(n20497));
    INVX1 U7626 (.I(N12140), .ZN(n20498));
    INVX1 U7627 (.I(N12141), .ZN(n20499));
    INVX1 U7628 (.I(N12142), .ZN(n20500));
    INVX1 U7629 (.I(N12143), .ZN(n20501));
    INVX1 U7630 (.I(N12144), .ZN(n20502));
    INVX1 U7631 (.I(N12145), .ZN(n20503));
    INVX1 U7632 (.I(N12146), .ZN(n20504));
    INVX1 U7633 (.I(N12147), .ZN(n20505));
    INVX1 U7634 (.I(N12148), .ZN(n20506));
    INVX1 U7635 (.I(N12149), .ZN(N20507));
    INVX1 U7636 (.I(N12150), .ZN(N20508));
    INVX1 U7637 (.I(N12151), .ZN(n20509));
    INVX1 U7638 (.I(N12152), .ZN(n20510));
    INVX1 U7639 (.I(N12153), .ZN(n20511));
    INVX1 U7640 (.I(N12154), .ZN(n20512));
    INVX1 U7641 (.I(N12155), .ZN(n20513));
    INVX1 U7642 (.I(N12156), .ZN(n20514));
    INVX1 U7643 (.I(N12157), .ZN(N20515));
    INVX1 U7644 (.I(N12158), .ZN(n20516));
    INVX1 U7645 (.I(N12159), .ZN(n20517));
    INVX1 U7646 (.I(N12160), .ZN(n20518));
    INVX1 U7647 (.I(N12161), .ZN(n20519));
    INVX1 U7648 (.I(N12162), .ZN(n20520));
    INVX1 U7649 (.I(N12163), .ZN(n20521));
    INVX1 U7650 (.I(N12164), .ZN(N20522));
    INVX1 U7651 (.I(N12165), .ZN(N20523));
    INVX1 U7652 (.I(N12166), .ZN(n20524));
    INVX1 U7653 (.I(N12167), .ZN(n20525));
    INVX1 U7654 (.I(N12168), .ZN(n20526));
    INVX1 U7655 (.I(N12169), .ZN(n20527));
    INVX1 U7656 (.I(N12170), .ZN(n20528));
    INVX1 U7657 (.I(N12171), .ZN(n20529));
    INVX1 U7658 (.I(N12172), .ZN(n20530));
    INVX1 U7659 (.I(N12173), .ZN(n20531));
    INVX1 U7660 (.I(N12174), .ZN(n20532));
    INVX1 U7661 (.I(N12175), .ZN(N20533));
    INVX1 U7662 (.I(N12176), .ZN(N20534));
    INVX1 U7663 (.I(N12177), .ZN(n20535));
    INVX1 U7664 (.I(N12178), .ZN(N20536));
    INVX1 U7665 (.I(N12179), .ZN(n20537));
    INVX1 U7666 (.I(N12180), .ZN(n20538));
    INVX1 U7667 (.I(N12181), .ZN(n20539));
    INVX1 U7668 (.I(N12182), .ZN(n20540));
    INVX1 U7669 (.I(N12183), .ZN(N20541));
    INVX1 U7670 (.I(N12184), .ZN(n20542));
    INVX1 U7671 (.I(N12185), .ZN(n20543));
    INVX1 U7672 (.I(N12186), .ZN(n20544));
    INVX1 U7673 (.I(N12187), .ZN(N20545));
    INVX1 U7674 (.I(N12188), .ZN(n20546));
    INVX1 U7675 (.I(N12189), .ZN(N20547));
    INVX1 U7676 (.I(N12190), .ZN(n20548));
    INVX1 U7677 (.I(N12191), .ZN(n20549));
    INVX1 U7678 (.I(N12192), .ZN(n20550));
    INVX1 U7679 (.I(N12193), .ZN(n20551));
    INVX1 U7680 (.I(N12194), .ZN(n20552));
    INVX1 U7681 (.I(N12195), .ZN(n20553));
    INVX1 U7682 (.I(N12196), .ZN(n20554));
    INVX1 U7683 (.I(N12197), .ZN(n20555));
    INVX1 U7684 (.I(N12198), .ZN(n20556));
    INVX1 U7685 (.I(N12199), .ZN(n20557));
    INVX1 U7686 (.I(N12200), .ZN(n20558));
    INVX1 U7687 (.I(N12201), .ZN(n20559));
    INVX1 U7688 (.I(N12202), .ZN(n20560));
    INVX1 U7689 (.I(N12203), .ZN(n20561));
    INVX1 U7690 (.I(N12204), .ZN(n20562));
    INVX1 U7691 (.I(N12205), .ZN(n20563));
    INVX1 U7692 (.I(N12206), .ZN(n20564));
    INVX1 U7693 (.I(N12207), .ZN(n20565));
    INVX1 U7694 (.I(N12208), .ZN(n20566));
    INVX1 U7695 (.I(N12209), .ZN(N20567));
    INVX1 U7696 (.I(N12210), .ZN(n20568));
    INVX1 U7697 (.I(N12211), .ZN(n20569));
    INVX1 U7698 (.I(N12212), .ZN(n20570));
    INVX1 U7699 (.I(N12213), .ZN(n20571));
    INVX1 U7700 (.I(N12214), .ZN(n20572));
    INVX1 U7701 (.I(N12215), .ZN(n20573));
    INVX1 U7702 (.I(N12216), .ZN(n20574));
    INVX1 U7703 (.I(N12217), .ZN(n20575));
    INVX1 U7704 (.I(N12218), .ZN(N20576));
    INVX1 U7705 (.I(N12219), .ZN(N20577));
    INVX1 U7706 (.I(N12220), .ZN(n20578));
    INVX1 U7707 (.I(N12221), .ZN(n20579));
    INVX1 U7708 (.I(N12222), .ZN(n20580));
    INVX1 U7709 (.I(N12223), .ZN(n20581));
    INVX1 U7710 (.I(N12224), .ZN(n20582));
    INVX1 U7711 (.I(N12225), .ZN(n20583));
    INVX1 U7712 (.I(N12226), .ZN(n20584));
    INVX1 U7713 (.I(N12227), .ZN(n20585));
    INVX1 U7714 (.I(N12228), .ZN(N20586));
    INVX1 U7715 (.I(N12229), .ZN(n20587));
    INVX1 U7716 (.I(N12230), .ZN(N20588));
    INVX1 U7717 (.I(N12231), .ZN(n20589));
    INVX1 U7718 (.I(N12232), .ZN(n20590));
    INVX1 U7719 (.I(N12233), .ZN(n20591));
    INVX1 U7720 (.I(N12234), .ZN(n20592));
    INVX1 U7721 (.I(N12235), .ZN(n20593));
    INVX1 U7722 (.I(N12236), .ZN(N20594));
    INVX1 U7723 (.I(N12237), .ZN(n20595));
    INVX1 U7724 (.I(N12238), .ZN(n20596));
    INVX1 U7725 (.I(N12239), .ZN(n20597));
    INVX1 U7726 (.I(N12240), .ZN(N20598));
    INVX1 U7727 (.I(N12241), .ZN(n20599));
    INVX1 U7728 (.I(N12242), .ZN(n20600));
    INVX1 U7729 (.I(N12243), .ZN(N20601));
    INVX1 U7730 (.I(N12244), .ZN(N20602));
    INVX1 U7731 (.I(N12245), .ZN(n20603));
    INVX1 U7732 (.I(N12246), .ZN(N20604));
    INVX1 U7733 (.I(N12247), .ZN(n20605));
    INVX1 U7734 (.I(N12248), .ZN(N20606));
    INVX1 U7735 (.I(N12249), .ZN(N20607));
    INVX1 U7736 (.I(N12250), .ZN(n20608));
    INVX1 U7737 (.I(N12251), .ZN(n20609));
    INVX1 U7738 (.I(N12252), .ZN(N20610));
    INVX1 U7739 (.I(N12253), .ZN(n20611));
    INVX1 U7740 (.I(N12254), .ZN(n20612));
    INVX1 U7741 (.I(N12255), .ZN(N20613));
    INVX1 U7742 (.I(N12256), .ZN(n20614));
    INVX1 U7743 (.I(N12257), .ZN(n20615));
    INVX1 U7744 (.I(N12258), .ZN(n20616));
    INVX1 U7745 (.I(N12259), .ZN(n20617));
    INVX1 U7746 (.I(N12260), .ZN(N20618));
    INVX1 U7747 (.I(N12261), .ZN(N20619));
    INVX1 U7748 (.I(N12262), .ZN(n20620));
    INVX1 U7749 (.I(N12263), .ZN(n20621));
    INVX1 U7750 (.I(N12264), .ZN(n20622));
    INVX1 U7751 (.I(N12265), .ZN(n20623));
    INVX1 U7752 (.I(N12266), .ZN(n20624));
    INVX1 U7753 (.I(N12267), .ZN(n20625));
    INVX1 U7754 (.I(N12268), .ZN(n20626));
    INVX1 U7755 (.I(N12269), .ZN(n20627));
    INVX1 U7756 (.I(N12270), .ZN(n20628));
    INVX1 U7757 (.I(N12271), .ZN(N20629));
    INVX1 U7758 (.I(N12272), .ZN(n20630));
    INVX1 U7759 (.I(N12273), .ZN(n20631));
    INVX1 U7760 (.I(N12274), .ZN(n20632));
    INVX1 U7761 (.I(N12275), .ZN(n20633));
    INVX1 U7762 (.I(N12276), .ZN(n20634));
    INVX1 U7763 (.I(N12277), .ZN(n20635));
    INVX1 U7764 (.I(N12278), .ZN(n20636));
    INVX1 U7765 (.I(N12279), .ZN(N20637));
    INVX1 U7766 (.I(N12280), .ZN(N20638));
    INVX1 U7767 (.I(N12281), .ZN(n20639));
    INVX1 U7768 (.I(N12282), .ZN(N20640));
    INVX1 U7769 (.I(N12283), .ZN(n20641));
    INVX1 U7770 (.I(N12284), .ZN(n20642));
    INVX1 U7771 (.I(N12285), .ZN(n20643));
    INVX1 U7772 (.I(N12286), .ZN(n20644));
    INVX1 U7773 (.I(N12287), .ZN(n20645));
    INVX1 U7774 (.I(N12288), .ZN(n20646));
    INVX1 U7775 (.I(N12289), .ZN(n20647));
    INVX1 U7776 (.I(N12290), .ZN(n20648));
    INVX1 U7777 (.I(N12291), .ZN(n20649));
    INVX1 U7778 (.I(N12292), .ZN(N20650));
    INVX1 U7779 (.I(N12293), .ZN(n20651));
    INVX1 U7780 (.I(N12294), .ZN(N20652));
    INVX1 U7781 (.I(N12295), .ZN(N20653));
    INVX1 U7782 (.I(N12296), .ZN(n20654));
    INVX1 U7783 (.I(N12297), .ZN(n20655));
    INVX1 U7784 (.I(N12298), .ZN(n20656));
    INVX1 U7785 (.I(N12299), .ZN(n20657));
    INVX1 U7786 (.I(N12300), .ZN(n20658));
    INVX1 U7787 (.I(N12301), .ZN(n20659));
    INVX1 U7788 (.I(N12302), .ZN(n20660));
    INVX1 U7789 (.I(N12303), .ZN(N20661));
    INVX1 U7790 (.I(N12304), .ZN(n20662));
    INVX1 U7791 (.I(N12305), .ZN(N20663));
    INVX1 U7792 (.I(N12306), .ZN(n20664));
    INVX1 U7793 (.I(N12307), .ZN(n20665));
    INVX1 U7794 (.I(N12308), .ZN(n20666));
    INVX1 U7795 (.I(N12309), .ZN(n20667));
    INVX1 U7796 (.I(N12310), .ZN(N20668));
    INVX1 U7797 (.I(N12311), .ZN(n20669));
    INVX1 U7798 (.I(N12312), .ZN(n20670));
    INVX1 U7799 (.I(N12313), .ZN(n20671));
    INVX1 U7800 (.I(N12314), .ZN(n20672));
    INVX1 U7801 (.I(N12315), .ZN(n20673));
    INVX1 U7802 (.I(N12316), .ZN(n20674));
    INVX1 U7803 (.I(N12317), .ZN(n20675));
    INVX1 U7804 (.I(N12318), .ZN(n20676));
    INVX1 U7805 (.I(N12319), .ZN(n20677));
    INVX1 U7806 (.I(N12320), .ZN(n20678));
    INVX1 U7807 (.I(N12321), .ZN(n20679));
    INVX1 U7808 (.I(N12322), .ZN(N20680));
    INVX1 U7809 (.I(N12323), .ZN(n20681));
    INVX1 U7810 (.I(N12324), .ZN(n20682));
    INVX1 U7811 (.I(N12325), .ZN(n20683));
    INVX1 U7812 (.I(N12326), .ZN(n20684));
    INVX1 U7813 (.I(N12327), .ZN(N20685));
    INVX1 U7814 (.I(N12328), .ZN(n20686));
    INVX1 U7815 (.I(N12329), .ZN(n20687));
    INVX1 U7816 (.I(N12330), .ZN(n20688));
    INVX1 U7817 (.I(N12331), .ZN(n20689));
    INVX1 U7818 (.I(N12332), .ZN(n20690));
    INVX1 U7819 (.I(N12333), .ZN(n20691));
    INVX1 U7820 (.I(N12334), .ZN(N20692));
    INVX1 U7821 (.I(N12335), .ZN(n20693));
    INVX1 U7822 (.I(N12336), .ZN(n20694));
    INVX1 U7823 (.I(N12337), .ZN(n20695));
    INVX1 U7824 (.I(N12338), .ZN(n20696));
    INVX1 U7825 (.I(N12339), .ZN(n20697));
    INVX1 U7826 (.I(N12340), .ZN(n20698));
    INVX1 U7827 (.I(N12341), .ZN(n20699));
    INVX1 U7828 (.I(N12342), .ZN(n20700));
    INVX1 U7829 (.I(N12343), .ZN(n20701));
    INVX1 U7830 (.I(N12344), .ZN(n20702));
    INVX1 U7831 (.I(N12345), .ZN(N20703));
    INVX1 U7832 (.I(N12346), .ZN(n20704));
    INVX1 U7833 (.I(N12347), .ZN(n20705));
    INVX1 U7834 (.I(N12348), .ZN(n20706));
    INVX1 U7835 (.I(N12349), .ZN(n20707));
    INVX1 U7836 (.I(N12350), .ZN(n20708));
    INVX1 U7837 (.I(N12351), .ZN(n20709));
    INVX1 U7838 (.I(N12352), .ZN(N20710));
    INVX1 U7839 (.I(N12353), .ZN(n20711));
    INVX1 U7840 (.I(N12354), .ZN(n20712));
    INVX1 U7841 (.I(N12355), .ZN(n20713));
    INVX1 U7842 (.I(N12356), .ZN(n20714));
    INVX1 U7843 (.I(N12357), .ZN(n20715));
    INVX1 U7844 (.I(N12358), .ZN(n20716));
    INVX1 U7845 (.I(N12359), .ZN(n20717));
    INVX1 U7846 (.I(N12360), .ZN(n20718));
    INVX1 U7847 (.I(N12361), .ZN(n20719));
    INVX1 U7848 (.I(N12362), .ZN(n20720));
    INVX1 U7849 (.I(N12363), .ZN(n20721));
    INVX1 U7850 (.I(N12364), .ZN(n20722));
    INVX1 U7851 (.I(N12365), .ZN(n20723));
    INVX1 U7852 (.I(N12366), .ZN(n20724));
    INVX1 U7853 (.I(N12367), .ZN(n20725));
    INVX1 U7854 (.I(N12368), .ZN(n20726));
    INVX1 U7855 (.I(N12369), .ZN(N20727));
    INVX1 U7856 (.I(N12370), .ZN(n20728));
    INVX1 U7857 (.I(N12371), .ZN(n20729));
    INVX1 U7858 (.I(N12372), .ZN(n20730));
    INVX1 U7859 (.I(N12373), .ZN(n20731));
    INVX1 U7860 (.I(N12374), .ZN(n20732));
    INVX1 U7861 (.I(N12375), .ZN(n20733));
    INVX1 U7862 (.I(N12376), .ZN(n20734));
    INVX1 U7863 (.I(N12377), .ZN(n20735));
    INVX1 U7864 (.I(N12378), .ZN(n20736));
    INVX1 U7865 (.I(N12379), .ZN(n20737));
    INVX1 U7866 (.I(N12380), .ZN(n20738));
    INVX1 U7867 (.I(N12381), .ZN(n20739));
    INVX1 U7868 (.I(N12382), .ZN(n20740));
    INVX1 U7869 (.I(N12383), .ZN(n20741));
    INVX1 U7870 (.I(N12384), .ZN(n20742));
    INVX1 U7871 (.I(N12385), .ZN(n20743));
    INVX1 U7872 (.I(N12386), .ZN(N20744));
    INVX1 U7873 (.I(N12387), .ZN(n20745));
    INVX1 U7874 (.I(N12388), .ZN(n20746));
    INVX1 U7875 (.I(N12389), .ZN(N20747));
    INVX1 U7876 (.I(N12390), .ZN(N20748));
    INVX1 U7877 (.I(N12391), .ZN(n20749));
    INVX1 U7878 (.I(N12392), .ZN(n20750));
    INVX1 U7879 (.I(N12393), .ZN(n20751));
    INVX1 U7880 (.I(N12394), .ZN(n20752));
    INVX1 U7881 (.I(N12395), .ZN(n20753));
    INVX1 U7882 (.I(N12396), .ZN(n20754));
    INVX1 U7883 (.I(N12397), .ZN(n20755));
    INVX1 U7884 (.I(N12398), .ZN(n20756));
    INVX1 U7885 (.I(N12399), .ZN(n20757));
    INVX1 U7886 (.I(N12400), .ZN(n20758));
    INVX1 U7887 (.I(N12401), .ZN(n20759));
    INVX1 U7888 (.I(N12402), .ZN(n20760));
    INVX1 U7889 (.I(N12403), .ZN(n20761));
    INVX1 U7890 (.I(N12404), .ZN(n20762));
    INVX1 U7891 (.I(N12405), .ZN(n20763));
    INVX1 U7892 (.I(N12406), .ZN(n20764));
    INVX1 U7893 (.I(N12407), .ZN(n20765));
    INVX1 U7894 (.I(N12408), .ZN(n20766));
    INVX1 U7895 (.I(N12409), .ZN(n20767));
    INVX1 U7896 (.I(N12410), .ZN(n20768));
    INVX1 U7897 (.I(N12411), .ZN(n20769));
    INVX1 U7898 (.I(N12412), .ZN(n20770));
    INVX1 U7899 (.I(N12413), .ZN(N20771));
    INVX1 U7900 (.I(N12414), .ZN(n20772));
    INVX1 U7901 (.I(N12415), .ZN(N20773));
    INVX1 U7902 (.I(N12416), .ZN(n20774));
    INVX1 U7903 (.I(N12417), .ZN(n20775));
    INVX1 U7904 (.I(N12418), .ZN(N20776));
    INVX1 U7905 (.I(N12419), .ZN(n20777));
    INVX1 U7906 (.I(N12420), .ZN(n20778));
    INVX1 U7907 (.I(N12421), .ZN(n20779));
    INVX1 U7908 (.I(N12422), .ZN(n20780));
    INVX1 U7909 (.I(N12423), .ZN(n20781));
    INVX1 U7910 (.I(N12424), .ZN(n20782));
    INVX1 U7911 (.I(N12425), .ZN(N20783));
    INVX1 U7912 (.I(N12426), .ZN(n20784));
    INVX1 U7913 (.I(N12427), .ZN(n20785));
    INVX1 U7914 (.I(N12428), .ZN(n20786));
    INVX1 U7915 (.I(N12429), .ZN(N20787));
    INVX1 U7916 (.I(N12430), .ZN(n20788));
    INVX1 U7917 (.I(N12431), .ZN(n20789));
    INVX1 U7918 (.I(N12432), .ZN(n20790));
    INVX1 U7919 (.I(N12433), .ZN(N20791));
    INVX1 U7920 (.I(N12434), .ZN(n20792));
    INVX1 U7921 (.I(N12435), .ZN(n20793));
    INVX1 U7922 (.I(N12436), .ZN(n20794));
    INVX1 U7923 (.I(N12437), .ZN(n20795));
    INVX1 U7924 (.I(N12438), .ZN(n20796));
    INVX1 U7925 (.I(N12439), .ZN(n20797));
    INVX1 U7926 (.I(N12440), .ZN(n20798));
    INVX1 U7927 (.I(N12441), .ZN(N20799));
    INVX1 U7928 (.I(N12442), .ZN(n20800));
    INVX1 U7929 (.I(N12443), .ZN(n20801));
    INVX1 U7930 (.I(N12444), .ZN(n20802));
    INVX1 U7931 (.I(N12445), .ZN(N20803));
    INVX1 U7932 (.I(N12446), .ZN(n20804));
    INVX1 U7933 (.I(N12447), .ZN(n20805));
    INVX1 U7934 (.I(N12448), .ZN(N20806));
    INVX1 U7935 (.I(N12449), .ZN(N20807));
    INVX1 U7936 (.I(N12450), .ZN(N20808));
    INVX1 U7937 (.I(N12451), .ZN(n20809));
    INVX1 U7938 (.I(N12452), .ZN(n20810));
    INVX1 U7939 (.I(N12453), .ZN(n20811));
    INVX1 U7940 (.I(N12454), .ZN(n20812));
    INVX1 U7941 (.I(N12455), .ZN(n20813));
    INVX1 U7942 (.I(N12456), .ZN(n20814));
    INVX1 U7943 (.I(N12457), .ZN(n20815));
    INVX1 U7944 (.I(N12458), .ZN(N20816));
    INVX1 U7945 (.I(N12459), .ZN(n20817));
    INVX1 U7946 (.I(N12460), .ZN(N20818));
    INVX1 U7947 (.I(N12461), .ZN(n20819));
    INVX1 U7948 (.I(N12462), .ZN(n20820));
    INVX1 U7949 (.I(N12463), .ZN(n20821));
    INVX1 U7950 (.I(N12464), .ZN(n20822));
    INVX1 U7951 (.I(N12465), .ZN(N20823));
    INVX1 U7952 (.I(N12466), .ZN(N20824));
    INVX1 U7953 (.I(N12467), .ZN(n20825));
    INVX1 U7954 (.I(N12468), .ZN(n20826));
    INVX1 U7955 (.I(N12469), .ZN(n20827));
    INVX1 U7956 (.I(N12470), .ZN(n20828));
    INVX1 U7957 (.I(N12471), .ZN(n20829));
    INVX1 U7958 (.I(N12472), .ZN(n20830));
    INVX1 U7959 (.I(N12473), .ZN(n20831));
    INVX1 U7960 (.I(N12474), .ZN(n20832));
    INVX1 U7961 (.I(N12475), .ZN(n20833));
    INVX1 U7962 (.I(N12476), .ZN(n20834));
    INVX1 U7963 (.I(N12477), .ZN(n20835));
    INVX1 U7964 (.I(N12478), .ZN(n20836));
    INVX1 U7965 (.I(N12479), .ZN(n20837));
    INVX1 U7966 (.I(N12480), .ZN(n20838));
    INVX1 U7967 (.I(N12481), .ZN(n20839));
    INVX1 U7968 (.I(N12482), .ZN(n20840));
    INVX1 U7969 (.I(N12483), .ZN(n20841));
    INVX1 U7970 (.I(N12484), .ZN(n20842));
    INVX1 U7971 (.I(N12485), .ZN(N20843));
    INVX1 U7972 (.I(N12486), .ZN(n20844));
    INVX1 U7973 (.I(N12487), .ZN(n20845));
    INVX1 U7974 (.I(N12488), .ZN(n20846));
    INVX1 U7975 (.I(N12489), .ZN(n20847));
    INVX1 U7976 (.I(N12490), .ZN(n20848));
    INVX1 U7977 (.I(N12491), .ZN(n20849));
    INVX1 U7978 (.I(N12492), .ZN(n20850));
    INVX1 U7979 (.I(N12493), .ZN(N20851));
    INVX1 U7980 (.I(N12494), .ZN(n20852));
    INVX1 U7981 (.I(N12495), .ZN(n20853));
    INVX1 U7982 (.I(N12496), .ZN(n20854));
    INVX1 U7983 (.I(N12497), .ZN(n20855));
    INVX1 U7984 (.I(N12498), .ZN(n20856));
    INVX1 U7985 (.I(N12499), .ZN(n20857));
    INVX1 U7986 (.I(N12500), .ZN(n20858));
    INVX1 U7987 (.I(N12501), .ZN(n20859));
    INVX1 U7988 (.I(N12502), .ZN(n20860));
    INVX1 U7989 (.I(N12503), .ZN(n20861));
    INVX1 U7990 (.I(N12504), .ZN(n20862));
    INVX1 U7991 (.I(N12505), .ZN(N20863));
    INVX1 U7992 (.I(N12506), .ZN(N20864));
    INVX1 U7993 (.I(N12507), .ZN(n20865));
    INVX1 U7994 (.I(N12508), .ZN(n20866));
    INVX1 U7995 (.I(N12509), .ZN(n20867));
    INVX1 U7996 (.I(N12510), .ZN(n20868));
    INVX1 U7997 (.I(N12511), .ZN(n20869));
    INVX1 U7998 (.I(N12512), .ZN(N20870));
    INVX1 U7999 (.I(N12513), .ZN(n20871));
    INVX1 U8000 (.I(N12514), .ZN(n20872));
    INVX1 U8001 (.I(N12515), .ZN(N20873));
    INVX1 U8002 (.I(N12516), .ZN(N20874));
    INVX1 U8003 (.I(N12517), .ZN(n20875));
    INVX1 U8004 (.I(N12518), .ZN(n20876));
    INVX1 U8005 (.I(N12519), .ZN(n20877));
    INVX1 U8006 (.I(N12520), .ZN(n20878));
    INVX1 U8007 (.I(N12521), .ZN(n20879));
    INVX1 U8008 (.I(N12522), .ZN(n20880));
    INVX1 U8009 (.I(N12523), .ZN(n20881));
    INVX1 U8010 (.I(N12524), .ZN(n20882));
    INVX1 U8011 (.I(N12525), .ZN(n20883));
    INVX1 U8012 (.I(N12526), .ZN(n20884));
    INVX1 U8013 (.I(N12527), .ZN(n20885));
    INVX1 U8014 (.I(N12528), .ZN(n20886));
    INVX1 U8015 (.I(N12529), .ZN(n20887));
    INVX1 U8016 (.I(N12530), .ZN(N20888));
    INVX1 U8017 (.I(N12531), .ZN(n20889));
    INVX1 U8018 (.I(N12532), .ZN(n20890));
    INVX1 U8019 (.I(N12533), .ZN(n20891));
    INVX1 U8020 (.I(N12534), .ZN(n20892));
    INVX1 U8021 (.I(N12535), .ZN(N20893));
    INVX1 U8022 (.I(N12536), .ZN(n20894));
    INVX1 U8023 (.I(N12537), .ZN(n20895));
    INVX1 U8024 (.I(N12538), .ZN(n20896));
    INVX1 U8025 (.I(N12539), .ZN(n20897));
    INVX1 U8026 (.I(N12540), .ZN(n20898));
    INVX1 U8027 (.I(N12541), .ZN(n20899));
    INVX1 U8028 (.I(N12542), .ZN(N20900));
    INVX1 U8029 (.I(N12543), .ZN(n20901));
    INVX1 U8030 (.I(N12544), .ZN(N20902));
    INVX1 U8031 (.I(N12545), .ZN(n20903));
    INVX1 U8032 (.I(N12546), .ZN(n20904));
    INVX1 U8033 (.I(N12547), .ZN(n20905));
    INVX1 U8034 (.I(N12548), .ZN(N20906));
    INVX1 U8035 (.I(N12549), .ZN(n20907));
    INVX1 U8036 (.I(N12550), .ZN(n20908));
    INVX1 U8037 (.I(N12551), .ZN(n20909));
    INVX1 U8038 (.I(N12552), .ZN(n20910));
    INVX1 U8039 (.I(N12553), .ZN(N20911));
    INVX1 U8040 (.I(N12554), .ZN(n20912));
    INVX1 U8041 (.I(N12555), .ZN(n20913));
    INVX1 U8042 (.I(N12556), .ZN(n20914));
    INVX1 U8043 (.I(N12557), .ZN(n20915));
    INVX1 U8044 (.I(N12558), .ZN(N20916));
    INVX1 U8045 (.I(N12559), .ZN(n20917));
    INVX1 U8046 (.I(N12560), .ZN(n20918));
    INVX1 U8047 (.I(N12561), .ZN(n20919));
    INVX1 U8048 (.I(N12562), .ZN(n20920));
    INVX1 U8049 (.I(N12563), .ZN(N20921));
    INVX1 U8050 (.I(N12564), .ZN(n20922));
    INVX1 U8051 (.I(N12565), .ZN(n20923));
    INVX1 U8052 (.I(N12566), .ZN(N20924));
    INVX1 U8053 (.I(N12567), .ZN(n20925));
    INVX1 U8054 (.I(N12568), .ZN(n20926));
    INVX1 U8055 (.I(N12569), .ZN(n20927));
    INVX1 U8056 (.I(N12570), .ZN(n20928));
    INVX1 U8057 (.I(N12571), .ZN(n20929));
    INVX1 U8058 (.I(N12572), .ZN(n20930));
    INVX1 U8059 (.I(N12573), .ZN(n20931));
    INVX1 U8060 (.I(N12574), .ZN(n20932));
    INVX1 U8061 (.I(N12575), .ZN(N20933));
    INVX1 U8062 (.I(N12576), .ZN(n20934));
    INVX1 U8063 (.I(N12577), .ZN(N20935));
    INVX1 U8064 (.I(N12578), .ZN(n20936));
    INVX1 U8065 (.I(N12579), .ZN(n20937));
    INVX1 U8066 (.I(N12580), .ZN(N20938));
    INVX1 U8067 (.I(N12581), .ZN(n20939));
    INVX1 U8068 (.I(N12582), .ZN(n20940));
    INVX1 U8069 (.I(N12583), .ZN(N20941));
    INVX1 U8070 (.I(N12584), .ZN(n20942));
    INVX1 U8071 (.I(N12585), .ZN(n20943));
    INVX1 U8072 (.I(N12586), .ZN(n20944));
    INVX1 U8073 (.I(N12587), .ZN(n20945));
    INVX1 U8074 (.I(N12588), .ZN(n20946));
    INVX1 U8075 (.I(N12589), .ZN(n20947));
    INVX1 U8076 (.I(N12590), .ZN(n20948));
    INVX1 U8077 (.I(N12591), .ZN(n20949));
    INVX1 U8078 (.I(N12592), .ZN(n20950));
    INVX1 U8079 (.I(N12593), .ZN(n20951));
    INVX1 U8080 (.I(N12594), .ZN(N20952));
    INVX1 U8081 (.I(N12595), .ZN(n20953));
    INVX1 U8082 (.I(N12596), .ZN(n20954));
    INVX1 U8083 (.I(N12597), .ZN(n20955));
    INVX1 U8084 (.I(N12598), .ZN(n20956));
    INVX1 U8085 (.I(N12599), .ZN(n20957));
    INVX1 U8086 (.I(N12600), .ZN(N20958));
    INVX1 U8087 (.I(N12601), .ZN(n20959));
    INVX1 U8088 (.I(N12602), .ZN(n20960));
    INVX1 U8089 (.I(N12603), .ZN(n20961));
    INVX1 U8090 (.I(N12604), .ZN(n20962));
    INVX1 U8091 (.I(N12605), .ZN(N20963));
    INVX1 U8092 (.I(N12606), .ZN(n20964));
    INVX1 U8093 (.I(N12607), .ZN(n20965));
    INVX1 U8094 (.I(N12608), .ZN(n20966));
    INVX1 U8095 (.I(N12609), .ZN(n20967));
    INVX1 U8096 (.I(N12610), .ZN(n20968));
    INVX1 U8097 (.I(N12611), .ZN(n20969));
    INVX1 U8098 (.I(N12612), .ZN(N20970));
    INVX1 U8099 (.I(N12613), .ZN(N20971));
    INVX1 U8100 (.I(N12614), .ZN(n20972));
    INVX1 U8101 (.I(N12615), .ZN(n20973));
    INVX1 U8102 (.I(N12616), .ZN(n20974));
    INVX1 U8103 (.I(N12617), .ZN(n20975));
    INVX1 U8104 (.I(N12618), .ZN(n20976));
    INVX1 U8105 (.I(N12619), .ZN(n20977));
    INVX1 U8106 (.I(N12620), .ZN(n20978));
    INVX1 U8107 (.I(N12621), .ZN(n20979));
    INVX1 U8108 (.I(N12622), .ZN(n20980));
    INVX1 U8109 (.I(N12623), .ZN(n20981));
    INVX1 U8110 (.I(N12624), .ZN(n20982));
    INVX1 U8111 (.I(N12625), .ZN(n20983));
    INVX1 U8112 (.I(N12626), .ZN(n20984));
    INVX1 U8113 (.I(N12627), .ZN(n20985));
    INVX1 U8114 (.I(N12628), .ZN(n20986));
    INVX1 U8115 (.I(N12629), .ZN(n20987));
    INVX1 U8116 (.I(N12630), .ZN(n20988));
    INVX1 U8117 (.I(N12631), .ZN(n20989));
    INVX1 U8118 (.I(N12632), .ZN(n20990));
    INVX1 U8119 (.I(N12633), .ZN(n20991));
    INVX1 U8120 (.I(N12634), .ZN(n20992));
    INVX1 U8121 (.I(N12635), .ZN(n20993));
    INVX1 U8122 (.I(N12636), .ZN(n20994));
    INVX1 U8123 (.I(N12637), .ZN(n20995));
    INVX1 U8124 (.I(N12638), .ZN(n20996));
    INVX1 U8125 (.I(N12639), .ZN(n20997));
    INVX1 U8126 (.I(N12640), .ZN(n20998));
    INVX1 U8127 (.I(N12641), .ZN(n20999));
    INVX1 U8128 (.I(N12642), .ZN(n21000));
    INVX1 U8129 (.I(N12643), .ZN(N21001));
    INVX1 U8130 (.I(N12644), .ZN(n21002));
    INVX1 U8131 (.I(N12645), .ZN(n21003));
    INVX1 U8132 (.I(N12646), .ZN(n21004));
    INVX1 U8133 (.I(N12647), .ZN(n21005));
    INVX1 U8134 (.I(N12648), .ZN(n21006));
    INVX1 U8135 (.I(N12649), .ZN(n21007));
    INVX1 U8136 (.I(N12650), .ZN(n21008));
    INVX1 U8137 (.I(N12651), .ZN(n21009));
    INVX1 U8138 (.I(N12652), .ZN(n21010));
    INVX1 U8139 (.I(N12653), .ZN(n21011));
    INVX1 U8140 (.I(N12654), .ZN(n21012));
    INVX1 U8141 (.I(N12655), .ZN(n21013));
    INVX1 U8142 (.I(N12656), .ZN(n21014));
    INVX1 U8143 (.I(N12657), .ZN(n21015));
    INVX1 U8144 (.I(N12658), .ZN(n21016));
    INVX1 U8145 (.I(N12659), .ZN(n21017));
    INVX1 U8146 (.I(N12660), .ZN(n21018));
    INVX1 U8147 (.I(N12661), .ZN(N21019));
    INVX1 U8148 (.I(N12662), .ZN(n21020));
    INVX1 U8149 (.I(N12663), .ZN(n21021));
    INVX1 U8150 (.I(N12664), .ZN(N21022));
    INVX1 U8151 (.I(N12665), .ZN(N21023));
    INVX1 U8152 (.I(N12666), .ZN(N21024));
    INVX1 U8153 (.I(N12667), .ZN(n21025));
    INVX1 U8154 (.I(N12668), .ZN(n21026));
    INVX1 U8155 (.I(N12669), .ZN(n21027));
    INVX1 U8156 (.I(N12670), .ZN(n21028));
    INVX1 U8157 (.I(N12671), .ZN(n21029));
    INVX1 U8158 (.I(N12672), .ZN(n21030));
    INVX1 U8159 (.I(N12673), .ZN(n21031));
    INVX1 U8160 (.I(N12674), .ZN(n21032));
    INVX1 U8161 (.I(N12675), .ZN(n21033));
    INVX1 U8162 (.I(N12676), .ZN(n21034));
    INVX1 U8163 (.I(N12677), .ZN(n21035));
    INVX1 U8164 (.I(N12678), .ZN(N21036));
    INVX1 U8165 (.I(N12679), .ZN(N21037));
    INVX1 U8166 (.I(N12680), .ZN(N21038));
    INVX1 U8167 (.I(N12681), .ZN(n21039));
    INVX1 U8168 (.I(N12682), .ZN(n21040));
    INVX1 U8169 (.I(N12683), .ZN(N21041));
    INVX1 U8170 (.I(N12684), .ZN(n21042));
    INVX1 U8171 (.I(N12685), .ZN(n21043));
    INVX1 U8172 (.I(N12686), .ZN(n21044));
    INVX1 U8173 (.I(N12687), .ZN(n21045));
    INVX1 U8174 (.I(N12688), .ZN(n21046));
    INVX1 U8175 (.I(N12689), .ZN(n21047));
    INVX1 U8176 (.I(N12690), .ZN(n21048));
    INVX1 U8177 (.I(N12691), .ZN(n21049));
    INVX1 U8178 (.I(N12692), .ZN(N21050));
    INVX1 U8179 (.I(N12693), .ZN(N21051));
    INVX1 U8180 (.I(N12694), .ZN(n21052));
    INVX1 U8181 (.I(N12695), .ZN(n21053));
    INVX1 U8182 (.I(N12696), .ZN(n21054));
    INVX1 U8183 (.I(N12697), .ZN(n21055));
    INVX1 U8184 (.I(N12698), .ZN(n21056));
    INVX1 U8185 (.I(N12699), .ZN(n21057));
    INVX1 U8186 (.I(N12700), .ZN(n21058));
    INVX1 U8187 (.I(N12701), .ZN(n21059));
    INVX1 U8188 (.I(N12702), .ZN(n21060));
    INVX1 U8189 (.I(N12703), .ZN(n21061));
    INVX1 U8190 (.I(N12704), .ZN(n21062));
    INVX1 U8191 (.I(N12705), .ZN(n21063));
    INVX1 U8192 (.I(N12706), .ZN(N21064));
    INVX1 U8193 (.I(N12707), .ZN(N21065));
    INVX1 U8194 (.I(N12708), .ZN(n21066));
    INVX1 U8195 (.I(N12709), .ZN(n21067));
    INVX1 U8196 (.I(N12710), .ZN(n21068));
    INVX1 U8197 (.I(N12711), .ZN(n21069));
    INVX1 U8198 (.I(N12712), .ZN(n21070));
    INVX1 U8199 (.I(N12713), .ZN(n21071));
    INVX1 U8200 (.I(N12714), .ZN(n21072));
    INVX1 U8201 (.I(N12715), .ZN(n21073));
    INVX1 U8202 (.I(N12716), .ZN(N21074));
    INVX1 U8203 (.I(N12717), .ZN(n21075));
    INVX1 U8204 (.I(N12718), .ZN(n21076));
    INVX1 U8205 (.I(N12719), .ZN(n21077));
    INVX1 U8206 (.I(N12720), .ZN(n21078));
    INVX1 U8207 (.I(N12721), .ZN(n21079));
    INVX1 U8208 (.I(N12722), .ZN(n21080));
    INVX1 U8209 (.I(N12723), .ZN(n21081));
    INVX1 U8210 (.I(N12724), .ZN(n21082));
    INVX1 U8211 (.I(N12725), .ZN(n21083));
    INVX1 U8212 (.I(N12726), .ZN(n21084));
    INVX1 U8213 (.I(N12727), .ZN(N21085));
    INVX1 U8214 (.I(N12728), .ZN(N21086));
    INVX1 U8215 (.I(N12729), .ZN(n21087));
    INVX1 U8216 (.I(N12730), .ZN(n21088));
    INVX1 U8217 (.I(N12731), .ZN(n21089));
    INVX1 U8218 (.I(N12732), .ZN(n21090));
    INVX1 U8219 (.I(N12733), .ZN(n21091));
    INVX1 U8220 (.I(N12734), .ZN(n21092));
    INVX1 U8221 (.I(N12735), .ZN(n21093));
    INVX1 U8222 (.I(N12736), .ZN(N21094));
    INVX1 U8223 (.I(N12737), .ZN(N21095));
    INVX1 U8224 (.I(N12738), .ZN(N21096));
    INVX1 U8225 (.I(N12739), .ZN(n21097));
    INVX1 U8226 (.I(N12740), .ZN(n21098));
    INVX1 U8227 (.I(N12741), .ZN(n21099));
    INVX1 U8228 (.I(N12742), .ZN(n21100));
    INVX1 U8229 (.I(N12743), .ZN(n21101));
    INVX1 U8230 (.I(N12744), .ZN(n21102));
    INVX1 U8231 (.I(N12745), .ZN(n21103));
    INVX1 U8232 (.I(N12746), .ZN(n21104));
    INVX1 U8233 (.I(N12747), .ZN(n21105));
    INVX1 U8234 (.I(N12748), .ZN(N21106));
    INVX1 U8235 (.I(N12749), .ZN(n21107));
    INVX1 U8236 (.I(N12750), .ZN(n21108));
    INVX1 U8237 (.I(N12751), .ZN(n21109));
    INVX1 U8238 (.I(N12752), .ZN(n21110));
    INVX1 U8239 (.I(N12753), .ZN(n21111));
    INVX1 U8240 (.I(N12754), .ZN(n21112));
    INVX1 U8241 (.I(N12755), .ZN(n21113));
    INVX1 U8242 (.I(N12756), .ZN(n21114));
    INVX1 U8243 (.I(N12757), .ZN(N21115));
    INVX1 U8244 (.I(N12758), .ZN(N21116));
    INVX1 U8245 (.I(N12759), .ZN(n21117));
    INVX1 U8246 (.I(N12760), .ZN(n21118));
    INVX1 U8247 (.I(N12761), .ZN(N21119));
    INVX1 U8248 (.I(N12762), .ZN(n21120));
    INVX1 U8249 (.I(N12763), .ZN(n21121));
    INVX1 U8250 (.I(N12764), .ZN(N21122));
    INVX1 U8251 (.I(N12765), .ZN(n21123));
    INVX1 U8252 (.I(N12766), .ZN(n21124));
    INVX1 U8253 (.I(N12767), .ZN(n21125));
    INVX1 U8254 (.I(N12768), .ZN(n21126));
    INVX1 U8255 (.I(N12769), .ZN(n21127));
    INVX1 U8256 (.I(N12770), .ZN(n21128));
    INVX1 U8257 (.I(N12771), .ZN(n21129));
    INVX1 U8258 (.I(N12772), .ZN(n21130));
    INVX1 U8259 (.I(N12773), .ZN(n21131));
    INVX1 U8260 (.I(N12774), .ZN(n21132));
    INVX1 U8261 (.I(N12775), .ZN(n21133));
    INVX1 U8262 (.I(N12776), .ZN(N21134));
    INVX1 U8263 (.I(N12777), .ZN(n21135));
    INVX1 U8264 (.I(N12778), .ZN(n21136));
    INVX1 U8265 (.I(N12779), .ZN(n21137));
    INVX1 U8266 (.I(N12780), .ZN(n21138));
    INVX1 U8267 (.I(N12781), .ZN(n21139));
    INVX1 U8268 (.I(N12782), .ZN(N21140));
    INVX1 U8269 (.I(N12783), .ZN(n21141));
    INVX1 U8270 (.I(N12784), .ZN(n21142));
    INVX1 U8271 (.I(N12785), .ZN(n21143));
    INVX1 U8272 (.I(N12786), .ZN(n21144));
    INVX1 U8273 (.I(N12787), .ZN(N21145));
    INVX1 U8274 (.I(N12788), .ZN(n21146));
    INVX1 U8275 (.I(N12789), .ZN(n21147));
    INVX1 U8276 (.I(N12790), .ZN(n21148));
    INVX1 U8277 (.I(N12791), .ZN(n21149));
    INVX1 U8278 (.I(N12792), .ZN(N21150));
    INVX1 U8279 (.I(N12793), .ZN(n21151));
    INVX1 U8280 (.I(N12794), .ZN(n21152));
    INVX1 U8281 (.I(N12795), .ZN(n21153));
    INVX1 U8282 (.I(N12796), .ZN(n21154));
    INVX1 U8283 (.I(N12797), .ZN(n21155));
    INVX1 U8284 (.I(N12798), .ZN(n21156));
    INVX1 U8285 (.I(N12799), .ZN(N21157));
    INVX1 U8286 (.I(N12800), .ZN(n21158));
    INVX1 U8287 (.I(N12801), .ZN(n21159));
    INVX1 U8288 (.I(N12802), .ZN(n21160));
    INVX1 U8289 (.I(N12803), .ZN(N21161));
    INVX1 U8290 (.I(N12804), .ZN(n21162));
    INVX1 U8291 (.I(N12805), .ZN(n21163));
    INVX1 U8292 (.I(N12806), .ZN(n21164));
    INVX1 U8293 (.I(N12807), .ZN(n21165));
    INVX1 U8294 (.I(N12808), .ZN(n21166));
    INVX1 U8295 (.I(N12809), .ZN(n21167));
    INVX1 U8296 (.I(N12810), .ZN(n21168));
    INVX1 U8297 (.I(N12811), .ZN(n21169));
    INVX1 U8298 (.I(N12812), .ZN(N21170));
    INVX1 U8299 (.I(N12813), .ZN(n21171));
    INVX1 U8300 (.I(N12814), .ZN(n21172));
    INVX1 U8301 (.I(N12815), .ZN(n21173));
    INVX1 U8302 (.I(N12816), .ZN(n21174));
    INVX1 U8303 (.I(N12817), .ZN(n21175));
    INVX1 U8304 (.I(N12818), .ZN(n21176));
    INVX1 U8305 (.I(N12819), .ZN(n21177));
    INVX1 U8306 (.I(N12820), .ZN(n21178));
    INVX1 U8307 (.I(N12821), .ZN(n21179));
    INVX1 U8308 (.I(N12822), .ZN(n21180));
    INVX1 U8309 (.I(N12823), .ZN(n21181));
    INVX1 U8310 (.I(N12824), .ZN(n21182));
    INVX1 U8311 (.I(N12825), .ZN(n21183));
    INVX1 U8312 (.I(N12826), .ZN(n21184));
    INVX1 U8313 (.I(N12827), .ZN(n21185));
    INVX1 U8314 (.I(N12828), .ZN(n21186));
    INVX1 U8315 (.I(N12829), .ZN(n21187));
    INVX1 U8316 (.I(N12830), .ZN(n21188));
    INVX1 U8317 (.I(N12831), .ZN(n21189));
    INVX1 U8318 (.I(N12832), .ZN(n21190));
    INVX1 U8319 (.I(N12833), .ZN(N21191));
    INVX1 U8320 (.I(N12834), .ZN(N21192));
    INVX1 U8321 (.I(N12835), .ZN(n21193));
    INVX1 U8322 (.I(N12836), .ZN(n21194));
    INVX1 U8323 (.I(N12837), .ZN(n21195));
    INVX1 U8324 (.I(N12838), .ZN(n21196));
    INVX1 U8325 (.I(N12839), .ZN(n21197));
    INVX1 U8326 (.I(N12840), .ZN(n21198));
    INVX1 U8327 (.I(N12841), .ZN(n21199));
    INVX1 U8328 (.I(N12842), .ZN(n21200));
    INVX1 U8329 (.I(N12843), .ZN(n21201));
    INVX1 U8330 (.I(N12844), .ZN(n21202));
    INVX1 U8331 (.I(N12845), .ZN(N21203));
    INVX1 U8332 (.I(N12846), .ZN(n21204));
    INVX1 U8333 (.I(N12847), .ZN(n21205));
    INVX1 U8334 (.I(N12848), .ZN(N21206));
    INVX1 U8335 (.I(N12849), .ZN(n21207));
    INVX1 U8336 (.I(N12850), .ZN(n21208));
    INVX1 U8337 (.I(N12851), .ZN(n21209));
    INVX1 U8338 (.I(N12852), .ZN(n21210));
    INVX1 U8339 (.I(N12853), .ZN(N21211));
    INVX1 U8340 (.I(N12854), .ZN(n21212));
    INVX1 U8341 (.I(N12855), .ZN(N21213));
    INVX1 U8342 (.I(N12856), .ZN(N21214));
    INVX1 U8343 (.I(N12857), .ZN(n21215));
    INVX1 U8344 (.I(N12858), .ZN(n21216));
    INVX1 U8345 (.I(N12859), .ZN(N21217));
    INVX1 U8346 (.I(N12860), .ZN(n21218));
    INVX1 U8347 (.I(N12861), .ZN(N21219));
    INVX1 U8348 (.I(N12862), .ZN(n21220));
    INVX1 U8349 (.I(N12863), .ZN(n21221));
    INVX1 U8350 (.I(N12864), .ZN(n21222));
    INVX1 U8351 (.I(N12865), .ZN(n21223));
    INVX1 U8352 (.I(N12866), .ZN(n21224));
    INVX1 U8353 (.I(N12867), .ZN(n21225));
    INVX1 U8354 (.I(N12868), .ZN(N21226));
    INVX1 U8355 (.I(N12869), .ZN(N21227));
    INVX1 U8356 (.I(N12870), .ZN(N21228));
    INVX1 U8357 (.I(N12871), .ZN(n21229));
    INVX1 U8358 (.I(N12872), .ZN(n21230));
    NOR2X1 U8359 (.A1(n18639), .A2(n18946), .ZN(N21231));
    NANDX1 U8360 (.A1(N4134), .A2(N3242), .ZN(n21232));
    NOR2X1 U8361 (.A1(N9230), .A2(n18152), .ZN(n21233));
    NANDX1 U8362 (.A1(N8227), .A2(N3680), .ZN(n21234));
    INVX1 U8363 (.I(n18974), .ZN(N21235));
    NOR2X1 U8364 (.A1(n13390), .A2(n16309), .ZN(n21236));
    NOR2X1 U8365 (.A1(n19778), .A2(N11330), .ZN(n21237));
    INVX1 U8366 (.I(N8891), .ZN(N21238));
    NANDX1 U8367 (.A1(n13133), .A2(N5587), .ZN(n21239));
    INVX1 U8368 (.I(n15650), .ZN(n21240));
    INVX1 U8369 (.I(n20334), .ZN(N21241));
    INVX1 U8370 (.I(N549), .ZN(n21242));
    NANDX1 U8371 (.A1(N10008), .A2(n19494), .ZN(n21243));
    NOR2X1 U8372 (.A1(N8684), .A2(n17277), .ZN(n21244));
    NOR2X1 U8373 (.A1(n17913), .A2(n14198), .ZN(n21245));
    INVX1 U8374 (.I(n20681), .ZN(n21246));
    NANDX1 U8375 (.A1(N12195), .A2(n12966), .ZN(n21247));
    NANDX1 U8376 (.A1(n20126), .A2(N2586), .ZN(N21248));
    INVX1 U8377 (.I(n18673), .ZN(n21249));
    NANDX1 U8378 (.A1(N11290), .A2(N875), .ZN(n21250));
    INVX1 U8379 (.I(n18965), .ZN(N21251));
    NANDX1 U8380 (.A1(n18586), .A2(n13384), .ZN(N21252));
    INVX1 U8381 (.I(N12231), .ZN(n21253));
    NANDX1 U8382 (.A1(N12734), .A2(N1995), .ZN(N21254));
    NOR2X1 U8383 (.A1(N10997), .A2(N943), .ZN(n21255));
    NOR2X1 U8384 (.A1(N7043), .A2(N10082), .ZN(n21256));
    NANDX1 U8385 (.A1(n15782), .A2(n14645), .ZN(N21257));
    NOR2X1 U8386 (.A1(N6970), .A2(N151), .ZN(n21258));
    NOR2X1 U8387 (.A1(n13575), .A2(n20276), .ZN(n21259));
    INVX1 U8388 (.I(N1302), .ZN(n21260));
    NOR2X1 U8389 (.A1(N11437), .A2(N7133), .ZN(N21261));
    INVX1 U8390 (.I(n14558), .ZN(n21262));
    NANDX1 U8391 (.A1(N8680), .A2(N6455), .ZN(n21263));
    NOR2X1 U8392 (.A1(n20865), .A2(n18686), .ZN(N21264));
    NOR2X1 U8393 (.A1(N12368), .A2(n15222), .ZN(n21265));
    NANDX1 U8394 (.A1(n17906), .A2(n16165), .ZN(n21266));
    NANDX1 U8395 (.A1(n19490), .A2(n20788), .ZN(n21267));
    INVX1 U8396 (.I(n14041), .ZN(n21268));
    NOR2X1 U8397 (.A1(n14782), .A2(n15552), .ZN(n21269));
    NOR2X1 U8398 (.A1(N9718), .A2(N7897), .ZN(N21270));
    NOR2X1 U8399 (.A1(N7239), .A2(N9198), .ZN(n21271));
    NOR2X1 U8400 (.A1(n13218), .A2(N10872), .ZN(n21272));
    NOR2X1 U8401 (.A1(N6545), .A2(N10281), .ZN(n21273));
    NOR2X1 U8402 (.A1(N7541), .A2(N1842), .ZN(N21274));
    INVX1 U8403 (.I(n20768), .ZN(n21275));
    NOR2X1 U8404 (.A1(N5494), .A2(n14760), .ZN(N21276));
    NANDX1 U8405 (.A1(N2169), .A2(N4236), .ZN(n21277));
    INVX1 U8406 (.I(N428), .ZN(n21278));
    NANDX1 U8407 (.A1(N1349), .A2(N9010), .ZN(n21279));
    NOR2X1 U8408 (.A1(n16130), .A2(N3332), .ZN(n21280));
    NOR2X1 U8409 (.A1(n20389), .A2(N5770), .ZN(n21281));
    NOR2X1 U8410 (.A1(N6398), .A2(N9509), .ZN(n21282));
    NANDX1 U8411 (.A1(n19615), .A2(n20380), .ZN(n21283));
    NOR2X1 U8412 (.A1(n20701), .A2(N9430), .ZN(N21284));
    NOR2X1 U8413 (.A1(N7011), .A2(N5814), .ZN(N21285));
    INVX1 U8414 (.I(N6549), .ZN(n21286));
    NOR2X1 U8415 (.A1(n15578), .A2(n15850), .ZN(N21287));
    NOR2X1 U8416 (.A1(n17747), .A2(n14627), .ZN(n21288));
    NOR2X1 U8417 (.A1(N12716), .A2(n12961), .ZN(n21289));
    NANDX1 U8418 (.A1(n16268), .A2(N4267), .ZN(n21290));
    NOR2X1 U8419 (.A1(n19599), .A2(n14781), .ZN(N21291));
    INVX1 U8420 (.I(n19910), .ZN(N21292));
    NOR2X1 U8421 (.A1(n19339), .A2(N8188), .ZN(n21293));
    NANDX1 U8422 (.A1(N12265), .A2(N1879), .ZN(n21294));
    INVX1 U8423 (.I(N11735), .ZN(n21295));
    INVX1 U8424 (.I(N10411), .ZN(N21296));
    INVX1 U8425 (.I(N11664), .ZN(n21297));
    INVX1 U8426 (.I(n14377), .ZN(n21298));
    NOR2X1 U8427 (.A1(N9385), .A2(N3538), .ZN(n21299));
    NOR2X1 U8428 (.A1(N443), .A2(N12706), .ZN(n21300));
    NOR2X1 U8429 (.A1(N7700), .A2(N4437), .ZN(n21301));
    NANDX1 U8430 (.A1(N2737), .A2(N3245), .ZN(N21302));
    INVX1 U8431 (.I(N1105), .ZN(n21303));
    NANDX1 U8432 (.A1(N11907), .A2(n21014), .ZN(N21304));
    NANDX1 U8433 (.A1(N4557), .A2(N2513), .ZN(n21305));
    INVX1 U8434 (.I(n16821), .ZN(N21306));
    NOR2X1 U8435 (.A1(n20157), .A2(N1867), .ZN(N21307));
    INVX1 U8436 (.I(N3879), .ZN(n21308));
    NOR2X1 U8437 (.A1(N675), .A2(n18916), .ZN(n21309));
    NANDX1 U8438 (.A1(n21162), .A2(N1612), .ZN(n21310));
    NANDX1 U8439 (.A1(N870), .A2(N2054), .ZN(n21311));
    NANDX1 U8440 (.A1(N9028), .A2(N9753), .ZN(n21312));
    INVX1 U8441 (.I(N4525), .ZN(n21313));
    NANDX1 U8442 (.A1(n15850), .A2(n19262), .ZN(n21314));
    NOR2X1 U8443 (.A1(N7186), .A2(N4481), .ZN(n21315));
    INVX1 U8444 (.I(N5067), .ZN(N21316));
    NOR2X1 U8445 (.A1(n20746), .A2(N10540), .ZN(n21317));
    INVX1 U8446 (.I(N3907), .ZN(n21318));
    NOR2X1 U8447 (.A1(N6494), .A2(N8690), .ZN(n21319));
    NANDX1 U8448 (.A1(n16189), .A2(N3906), .ZN(n21320));
    NANDX1 U8449 (.A1(n13573), .A2(N3838), .ZN(n21321));
    INVX1 U8450 (.I(N9036), .ZN(n21322));
    INVX1 U8451 (.I(n14092), .ZN(N21323));
    INVX1 U8452 (.I(N8276), .ZN(n21324));
    NANDX1 U8453 (.A1(N8579), .A2(N12800), .ZN(N21325));
    INVX1 U8454 (.I(n18970), .ZN(n21326));
    INVX1 U8455 (.I(N12323), .ZN(N21327));
    NOR2X1 U8456 (.A1(N9853), .A2(N9326), .ZN(n21328));
    INVX1 U8457 (.I(n18890), .ZN(n21329));
    NOR2X1 U8458 (.A1(n15073), .A2(N2287), .ZN(N21330));
    INVX1 U8459 (.I(n19081), .ZN(N21331));
    NANDX1 U8460 (.A1(N10521), .A2(N279), .ZN(N21332));
    NOR2X1 U8461 (.A1(n14427), .A2(n16164), .ZN(N21333));
    NOR2X1 U8462 (.A1(N12806), .A2(N12430), .ZN(N21334));
    NANDX1 U8463 (.A1(N12054), .A2(N5291), .ZN(n21335));
    NANDX1 U8464 (.A1(n20329), .A2(N2446), .ZN(N21336));
    INVX1 U8465 (.I(N6440), .ZN(n21337));
    INVX1 U8466 (.I(N1346), .ZN(n21338));
    NANDX1 U8467 (.A1(n13497), .A2(N6271), .ZN(n21339));
    NOR2X1 U8468 (.A1(n17364), .A2(n16262), .ZN(n21340));
    INVX1 U8469 (.I(n20746), .ZN(n21341));
    NOR2X1 U8470 (.A1(N10694), .A2(N1347), .ZN(n21342));
    NANDX1 U8471 (.A1(n14015), .A2(N6410), .ZN(n21343));
    NANDX1 U8472 (.A1(N1379), .A2(n20836), .ZN(n21344));
    NANDX1 U8473 (.A1(n18087), .A2(N12411), .ZN(n21345));
    INVX1 U8474 (.I(N1370), .ZN(n21346));
    NOR2X1 U8475 (.A1(N9968), .A2(N1857), .ZN(n21347));
    NANDX1 U8476 (.A1(N12414), .A2(N5463), .ZN(n21348));
    INVX1 U8477 (.I(n13588), .ZN(N21349));
    NANDX1 U8478 (.A1(N9666), .A2(N5854), .ZN(N21350));
    INVX1 U8479 (.I(N10100), .ZN(n21351));
    NOR2X1 U8480 (.A1(n18424), .A2(N2735), .ZN(N21352));
    NANDX1 U8481 (.A1(N1839), .A2(N7970), .ZN(n21353));
    NOR2X1 U8482 (.A1(N4335), .A2(N755), .ZN(N21354));
    INVX1 U8483 (.I(N1650), .ZN(n21355));
    NOR2X1 U8484 (.A1(N3405), .A2(n15129), .ZN(N21356));
    NOR2X1 U8485 (.A1(N10357), .A2(n19806), .ZN(N21357));
    NOR2X1 U8486 (.A1(N8132), .A2(N3086), .ZN(n21358));
    NOR2X1 U8487 (.A1(n20777), .A2(N10041), .ZN(n21359));
    NOR2X1 U8488 (.A1(n18631), .A2(N2398), .ZN(n21360));
    NANDX1 U8489 (.A1(N1608), .A2(N8251), .ZN(n21361));
    NOR2X1 U8490 (.A1(N6250), .A2(N4779), .ZN(N21362));
    NANDX1 U8491 (.A1(N3526), .A2(N822), .ZN(n21363));
    INVX1 U8492 (.I(N11496), .ZN(n21364));
    INVX1 U8493 (.I(n19411), .ZN(n21365));
    NOR2X1 U8494 (.A1(N2011), .A2(n21061), .ZN(n21366));
    NOR2X1 U8495 (.A1(n21187), .A2(N9501), .ZN(n21367));
    NANDX1 U8496 (.A1(N4855), .A2(N8076), .ZN(N21368));
    NANDX1 U8497 (.A1(N7528), .A2(N5703), .ZN(n21369));
    NANDX1 U8498 (.A1(N7074), .A2(n15743), .ZN(n21370));
    INVX1 U8499 (.I(n20246), .ZN(N21371));
    INVX1 U8500 (.I(N9612), .ZN(N21372));
    INVX1 U8501 (.I(n20932), .ZN(n21373));
    NANDX1 U8502 (.A1(N6873), .A2(N4480), .ZN(n21374));
    NOR2X1 U8503 (.A1(N4940), .A2(N5302), .ZN(n21375));
    NANDX1 U8504 (.A1(n16435), .A2(N3513), .ZN(n21376));
    INVX1 U8505 (.I(N1996), .ZN(N21377));
    INVX1 U8506 (.I(n20438), .ZN(n21378));
    INVX1 U8507 (.I(n15794), .ZN(n21379));
    INVX1 U8508 (.I(N2458), .ZN(n21380));
    NOR2X1 U8509 (.A1(N11326), .A2(N10127), .ZN(n21381));
    NANDX1 U8510 (.A1(n17028), .A2(N9095), .ZN(N21382));
    INVX1 U8511 (.I(N6083), .ZN(n21383));
    INVX1 U8512 (.I(N7577), .ZN(n21384));
    NANDX1 U8513 (.A1(N3519), .A2(N2742), .ZN(n21385));
    INVX1 U8514 (.I(n13403), .ZN(N21386));
    INVX1 U8515 (.I(N1715), .ZN(n21387));
    INVX1 U8516 (.I(N9096), .ZN(N21388));
    NANDX1 U8517 (.A1(n16493), .A2(N4300), .ZN(n21389));
    NANDX1 U8518 (.A1(n15870), .A2(N6296), .ZN(n21390));
    NANDX1 U8519 (.A1(N9620), .A2(N11757), .ZN(n21391));
    INVX1 U8520 (.I(N12869), .ZN(n21392));
    NANDX1 U8521 (.A1(N9431), .A2(n18736), .ZN(n21393));
    INVX1 U8522 (.I(n16377), .ZN(n21394));
    NANDX1 U8523 (.A1(n17061), .A2(N3708), .ZN(N21395));
    NOR2X1 U8524 (.A1(n16425), .A2(N5826), .ZN(n21396));
    NANDX1 U8525 (.A1(n19943), .A2(N3110), .ZN(N21397));
    NANDX1 U8526 (.A1(N6658), .A2(N7265), .ZN(n21398));
    NOR2X1 U8527 (.A1(N723), .A2(N10902), .ZN(N21399));
    INVX1 U8528 (.I(N11757), .ZN(n21400));
    NOR2X1 U8529 (.A1(N7352), .A2(N938), .ZN(n21401));
    NOR2X1 U8530 (.A1(N1571), .A2(N10557), .ZN(N21402));
    NOR2X1 U8531 (.A1(N11584), .A2(n17968), .ZN(n21403));
    INVX1 U8532 (.I(n21014), .ZN(N21404));
    INVX1 U8533 (.I(n17828), .ZN(n21405));
    NOR2X1 U8534 (.A1(n19090), .A2(n13658), .ZN(N21406));
    NOR2X1 U8535 (.A1(n13017), .A2(N8853), .ZN(n21407));
    NOR2X1 U8536 (.A1(N4478), .A2(N2107), .ZN(n21408));
    NANDX1 U8537 (.A1(N8945), .A2(N8764), .ZN(n21409));
    NOR2X1 U8538 (.A1(n15127), .A2(N4028), .ZN(n21410));
    NANDX1 U8539 (.A1(n17409), .A2(n15784), .ZN(n21411));
    NANDX1 U8540 (.A1(n19302), .A2(n16722), .ZN(n21412));
    INVX1 U8541 (.I(n15415), .ZN(n21413));
    INVX1 U8542 (.I(N9563), .ZN(n21414));
    INVX1 U8543 (.I(n18557), .ZN(n21415));
    INVX1 U8544 (.I(N93), .ZN(N21416));
    NOR2X1 U8545 (.A1(N5106), .A2(N10795), .ZN(n21417));
    NANDX1 U8546 (.A1(n18763), .A2(n19745), .ZN(n21418));
    INVX1 U8547 (.I(N6385), .ZN(n21419));
    NOR2X1 U8548 (.A1(n17237), .A2(N3034), .ZN(n21420));
    INVX1 U8549 (.I(N4951), .ZN(N21421));
    INVX1 U8550 (.I(n13264), .ZN(n21422));
    INVX1 U8551 (.I(N10367), .ZN(n21423));
    NOR2X1 U8552 (.A1(N10798), .A2(N4920), .ZN(n21424));
    INVX1 U8553 (.I(N8869), .ZN(n21425));
    NOR2X1 U8554 (.A1(N12585), .A2(N3053), .ZN(N21426));
    INVX1 U8555 (.I(n16689), .ZN(n21427));
    NANDX1 U8556 (.A1(n14099), .A2(N3966), .ZN(n21428));
    NOR2X1 U8557 (.A1(N210), .A2(N9071), .ZN(n21429));
    INVX1 U8558 (.I(n21183), .ZN(n21430));
    NANDX1 U8559 (.A1(N1847), .A2(n18170), .ZN(n21431));
    NOR2X1 U8560 (.A1(N4222), .A2(N8718), .ZN(N21432));
    NOR2X1 U8561 (.A1(N3251), .A2(N8210), .ZN(N21433));
    NANDX1 U8562 (.A1(N11056), .A2(N1599), .ZN(n21434));
    INVX1 U8563 (.I(N6994), .ZN(n21435));
    INVX1 U8564 (.I(N5499), .ZN(n21436));
    INVX1 U8565 (.I(n15807), .ZN(n21437));
    NOR2X1 U8566 (.A1(N2476), .A2(n13401), .ZN(N21438));
    INVX1 U8567 (.I(n19164), .ZN(n21439));
    NANDX1 U8568 (.A1(N10092), .A2(N1900), .ZN(n21440));
    NANDX1 U8569 (.A1(N4844), .A2(N10970), .ZN(n21441));
    NOR2X1 U8570 (.A1(N4796), .A2(n17573), .ZN(n21442));
    NOR2X1 U8571 (.A1(n17507), .A2(n19645), .ZN(n21443));
    INVX1 U8572 (.I(N4994), .ZN(n21444));
    NOR2X1 U8573 (.A1(N721), .A2(N7745), .ZN(N21445));
    NANDX1 U8574 (.A1(N11776), .A2(N9344), .ZN(n21446));
    NOR2X1 U8575 (.A1(n13312), .A2(n16281), .ZN(n21447));
    NANDX1 U8576 (.A1(N3203), .A2(N5399), .ZN(n21448));
    INVX1 U8577 (.I(N5679), .ZN(n21449));
    NOR2X1 U8578 (.A1(N1712), .A2(n19384), .ZN(N21450));
    NANDX1 U8579 (.A1(N6345), .A2(n15825), .ZN(n21451));
    NOR2X1 U8580 (.A1(N5730), .A2(N5565), .ZN(N21452));
    NOR2X1 U8581 (.A1(N10525), .A2(n17679), .ZN(n21453));
    NANDX1 U8582 (.A1(N1343), .A2(n16093), .ZN(n21454));
    INVX1 U8583 (.I(N878), .ZN(n21455));
    INVX1 U8584 (.I(N11930), .ZN(n21456));
    NOR2X1 U8585 (.A1(n13343), .A2(n18247), .ZN(N21457));
    NANDX1 U8586 (.A1(n13112), .A2(N10328), .ZN(n21458));
    NOR2X1 U8587 (.A1(n12921), .A2(N8073), .ZN(N21459));
    NOR2X1 U8588 (.A1(n18639), .A2(N8293), .ZN(n21460));
    NANDX1 U8589 (.A1(n14892), .A2(N6446), .ZN(n21461));
    INVX1 U8590 (.I(n15778), .ZN(n21462));
    NANDX1 U8591 (.A1(n16342), .A2(N278), .ZN(n21463));
    NANDX1 U8592 (.A1(N4687), .A2(N5344), .ZN(n21464));
    NANDX1 U8593 (.A1(n18426), .A2(N6687), .ZN(N21465));
    NANDX1 U8594 (.A1(N2947), .A2(N2106), .ZN(N21466));
    NOR2X1 U8595 (.A1(N9418), .A2(N10728), .ZN(N21467));
    NANDX1 U8596 (.A1(N977), .A2(N2005), .ZN(N21468));
    NANDX1 U8597 (.A1(N11304), .A2(N9563), .ZN(N21469));
    NOR2X1 U8598 (.A1(n13918), .A2(n17061), .ZN(N21470));
    NANDX1 U8599 (.A1(N980), .A2(N6356), .ZN(n21471));
    NANDX1 U8600 (.A1(N1968), .A2(n20296), .ZN(n21472));
    NANDX1 U8601 (.A1(n18780), .A2(N9949), .ZN(n21473));
    NOR2X1 U8602 (.A1(n19926), .A2(n14635), .ZN(n21474));
    NANDX1 U8603 (.A1(N12062), .A2(N6372), .ZN(n21475));
    INVX1 U8604 (.I(n14833), .ZN(n21476));
    NANDX1 U8605 (.A1(N7807), .A2(N10527), .ZN(n21477));
    INVX1 U8606 (.I(n13076), .ZN(n21478));
    NOR2X1 U8607 (.A1(N8796), .A2(n15081), .ZN(n21479));
    INVX1 U8608 (.I(n20100), .ZN(n21480));
    NANDX1 U8609 (.A1(n13089), .A2(N7329), .ZN(N21481));
    NANDX1 U8610 (.A1(n18876), .A2(N8309), .ZN(n21482));
    INVX1 U8611 (.I(N12867), .ZN(N21483));
    NANDX1 U8612 (.A1(N9519), .A2(n17177), .ZN(n21484));
    INVX1 U8613 (.I(n14009), .ZN(N21485));
    INVX1 U8614 (.I(n16834), .ZN(n21486));
    NOR2X1 U8615 (.A1(n20778), .A2(N2207), .ZN(n21487));
    NANDX1 U8616 (.A1(N5249), .A2(n17040), .ZN(n21488));
    NOR2X1 U8617 (.A1(n13055), .A2(N878), .ZN(n21489));
    NANDX1 U8618 (.A1(n20672), .A2(N4669), .ZN(n21490));
    NANDX1 U8619 (.A1(n14522), .A2(N3920), .ZN(N21491));
    NANDX1 U8620 (.A1(N7018), .A2(n17008), .ZN(n21492));
    INVX1 U8621 (.I(n16574), .ZN(n21493));
    NANDX1 U8622 (.A1(N5703), .A2(N11255), .ZN(n21494));
    NOR2X1 U8623 (.A1(N5062), .A2(n15315), .ZN(n21495));
    INVX1 U8624 (.I(N7428), .ZN(n21496));
    NANDX1 U8625 (.A1(N7624), .A2(n18803), .ZN(n21497));
    INVX1 U8626 (.I(N7172), .ZN(N21498));
    NOR2X1 U8627 (.A1(n12915), .A2(N6962), .ZN(n21499));
    NANDX1 U8628 (.A1(n19642), .A2(n14558), .ZN(n21500));
    NANDX1 U8629 (.A1(N7501), .A2(n13999), .ZN(n21501));
    INVX1 U8630 (.I(N9614), .ZN(n21502));
    NOR2X1 U8631 (.A1(N9909), .A2(n20909), .ZN(N21503));
    INVX1 U8632 (.I(N5686), .ZN(n21504));
    NANDX1 U8633 (.A1(n19966), .A2(N9423), .ZN(n21505));
    INVX1 U8634 (.I(N9990), .ZN(n21506));
    NOR2X1 U8635 (.A1(N7836), .A2(n19847), .ZN(n21507));
    INVX1 U8636 (.I(N9805), .ZN(n21508));
    NOR2X1 U8637 (.A1(n19509), .A2(N7377), .ZN(N21509));
    INVX1 U8638 (.I(n21222), .ZN(n21510));
    NANDX1 U8639 (.A1(N2982), .A2(N6953), .ZN(n21511));
    INVX1 U8640 (.I(n17165), .ZN(n21512));
    INVX1 U8641 (.I(n19836), .ZN(n21513));
    INVX1 U8642 (.I(N8821), .ZN(n21514));
    INVX1 U8643 (.I(N7591), .ZN(n21515));
    NANDX1 U8644 (.A1(n14504), .A2(N7269), .ZN(N21516));
    NOR2X1 U8645 (.A1(n14732), .A2(N4342), .ZN(n21517));
    NANDX1 U8646 (.A1(N2924), .A2(N1658), .ZN(N21518));
    NOR2X1 U8647 (.A1(N2260), .A2(N9494), .ZN(n21519));
    INVX1 U8648 (.I(n19603), .ZN(n21520));
    NANDX1 U8649 (.A1(N1405), .A2(n17882), .ZN(N21521));
    INVX1 U8650 (.I(N12702), .ZN(n21522));
    NOR2X1 U8651 (.A1(N1684), .A2(N10225), .ZN(N21523));
    INVX1 U8652 (.I(N3824), .ZN(n21524));
    NANDX1 U8653 (.A1(n14189), .A2(n18202), .ZN(n21525));
    NOR2X1 U8654 (.A1(n17551), .A2(N1567), .ZN(n21526));
    NOR2X1 U8655 (.A1(N6973), .A2(N10612), .ZN(N21527));
    NANDX1 U8656 (.A1(n15559), .A2(n19885), .ZN(n21528));
    INVX1 U8657 (.I(N7107), .ZN(n21529));
    INVX1 U8658 (.I(n14078), .ZN(N21530));
    NOR2X1 U8659 (.A1(n19610), .A2(n18113), .ZN(n21531));
    INVX1 U8660 (.I(n17982), .ZN(n21532));
    INVX1 U8661 (.I(n15060), .ZN(n21533));
    NANDX1 U8662 (.A1(N10708), .A2(N1073), .ZN(n21534));
    NANDX1 U8663 (.A1(N6933), .A2(N11298), .ZN(n21535));
    NOR2X1 U8664 (.A1(N10757), .A2(N11999), .ZN(n21536));
    INVX1 U8665 (.I(N7728), .ZN(N21537));
    NANDX1 U8666 (.A1(n19320), .A2(N3836), .ZN(N21538));
    NANDX1 U8667 (.A1(n20834), .A2(n14447), .ZN(n21539));
    INVX1 U8668 (.I(N9704), .ZN(N21540));
    NANDX1 U8669 (.A1(N441), .A2(n16811), .ZN(n21541));
    NANDX1 U8670 (.A1(N9060), .A2(n14539), .ZN(n21542));
    INVX1 U8671 (.I(N5942), .ZN(n21543));
    NOR2X1 U8672 (.A1(n20124), .A2(N11205), .ZN(n21544));
    INVX1 U8673 (.I(N2610), .ZN(n21545));
    INVX1 U8674 (.I(N12179), .ZN(N21546));
    INVX1 U8675 (.I(N2157), .ZN(N21547));
    INVX1 U8676 (.I(N11779), .ZN(n21548));
    NOR2X1 U8677 (.A1(N8786), .A2(N8090), .ZN(n21549));
    NANDX1 U8678 (.A1(N3690), .A2(N6179), .ZN(n21550));
    INVX1 U8679 (.I(N4862), .ZN(n21551));
    INVX1 U8680 (.I(n17090), .ZN(n21552));
    INVX1 U8681 (.I(N10028), .ZN(n21553));
    INVX1 U8682 (.I(N3637), .ZN(n21554));
    INVX1 U8683 (.I(N7265), .ZN(N21555));
    NANDX1 U8684 (.A1(N9230), .A2(n14865), .ZN(n21556));
    NOR2X1 U8685 (.A1(N10735), .A2(N8300), .ZN(n21557));
    INVX1 U8686 (.I(N611), .ZN(n21558));
    NOR2X1 U8687 (.A1(n19607), .A2(N12790), .ZN(n21559));
    INVX1 U8688 (.I(n16306), .ZN(n21560));
    INVX1 U8689 (.I(n14740), .ZN(N21561));
    NANDX1 U8690 (.A1(n18363), .A2(n17371), .ZN(N21562));
    NANDX1 U8691 (.A1(n16594), .A2(n18091), .ZN(n21563));
    NANDX1 U8692 (.A1(n15998), .A2(n18415), .ZN(n21564));
    INVX1 U8693 (.I(N3422), .ZN(n21565));
    NANDX1 U8694 (.A1(N3341), .A2(N7058), .ZN(N21566));
    NANDX1 U8695 (.A1(N10606), .A2(n19753), .ZN(N21567));
    NANDX1 U8696 (.A1(n20012), .A2(N6243), .ZN(n21568));
    NANDX1 U8697 (.A1(N7081), .A2(N3937), .ZN(N21569));
    NANDX1 U8698 (.A1(N12531), .A2(N2314), .ZN(n21570));
    NANDX1 U8699 (.A1(n15492), .A2(n13161), .ZN(N21571));
    INVX1 U8700 (.I(N3544), .ZN(n21572));
    NANDX1 U8701 (.A1(N4371), .A2(n15456), .ZN(n21573));
    NOR2X1 U8702 (.A1(n20964), .A2(N12317), .ZN(n21574));
    NOR2X1 U8703 (.A1(n15731), .A2(N4043), .ZN(n21575));
    NOR2X1 U8704 (.A1(n13694), .A2(N5796), .ZN(n21576));
    INVX1 U8705 (.I(n20751), .ZN(n21577));
    NOR2X1 U8706 (.A1(n18417), .A2(n13815), .ZN(n21578));
    INVX1 U8707 (.I(n17198), .ZN(n21579));
    NOR2X1 U8708 (.A1(N3091), .A2(N3048), .ZN(n21580));
    INVX1 U8709 (.I(n14652), .ZN(n21581));
    NANDX1 U8710 (.A1(n15391), .A2(n17771), .ZN(N21582));
    INVX1 U8711 (.I(N7321), .ZN(n21583));
    INVX1 U8712 (.I(n18239), .ZN(N21584));
    NOR2X1 U8713 (.A1(n13607), .A2(N12464), .ZN(N21585));
    NOR2X1 U8714 (.A1(N7883), .A2(n19322), .ZN(N21586));
    NOR2X1 U8715 (.A1(n18155), .A2(N2134), .ZN(n21587));
    NOR2X1 U8716 (.A1(N10619), .A2(N7929), .ZN(n21588));
    INVX1 U8717 (.I(N10139), .ZN(n21589));
    NANDX1 U8718 (.A1(N5616), .A2(n18496), .ZN(N21590));
    INVX1 U8719 (.I(N1583), .ZN(N21591));
    NOR2X1 U8720 (.A1(N10255), .A2(n20402), .ZN(n21592));
    NOR2X1 U8721 (.A1(n19448), .A2(N3834), .ZN(n21593));
    INVX1 U8722 (.I(n15989), .ZN(n21594));
    NANDX1 U8723 (.A1(N5191), .A2(N3995), .ZN(n21595));
    NANDX1 U8724 (.A1(N11827), .A2(N12144), .ZN(n21596));
    NANDX1 U8725 (.A1(n19115), .A2(n20026), .ZN(N21597));
    NANDX1 U8726 (.A1(n15263), .A2(n16950), .ZN(N21598));
    NOR2X1 U8727 (.A1(n15881), .A2(N6338), .ZN(n21599));
    NOR2X1 U8728 (.A1(n18853), .A2(N11019), .ZN(n21600));
    INVX1 U8729 (.I(N3238), .ZN(n21601));
    INVX1 U8730 (.I(n15881), .ZN(n21602));
    INVX1 U8731 (.I(n14689), .ZN(n21603));
    INVX1 U8732 (.I(N3992), .ZN(n21604));
    INVX1 U8733 (.I(n18895), .ZN(n21605));
    NOR2X1 U8734 (.A1(N5956), .A2(N8195), .ZN(n21606));
    NANDX1 U8735 (.A1(N5689), .A2(N12190), .ZN(N21607));
    INVX1 U8736 (.I(n17515), .ZN(n21608));
    INVX1 U8737 (.I(n16513), .ZN(N21609));
    NOR2X1 U8738 (.A1(n17670), .A2(N10458), .ZN(N21610));
    INVX1 U8739 (.I(N7931), .ZN(N21611));
    INVX1 U8740 (.I(n14395), .ZN(n21612));
    INVX1 U8741 (.I(N10543), .ZN(N21613));
    NANDX1 U8742 (.A1(n14371), .A2(n13802), .ZN(n21614));
    NANDX1 U8743 (.A1(n17196), .A2(N2994), .ZN(n21615));
    NOR2X1 U8744 (.A1(N10654), .A2(n18213), .ZN(n21616));
    INVX1 U8745 (.I(n13281), .ZN(N21617));
    NOR2X1 U8746 (.A1(n20975), .A2(n13779), .ZN(n21618));
    NANDX1 U8747 (.A1(n20639), .A2(n19467), .ZN(n21619));
    INVX1 U8748 (.I(n14610), .ZN(n21620));
    NANDX1 U8749 (.A1(N7217), .A2(N4434), .ZN(n21621));
    NANDX1 U8750 (.A1(n19428), .A2(n14891), .ZN(N21622));
    NANDX1 U8751 (.A1(N671), .A2(N196), .ZN(n21623));
    NANDX1 U8752 (.A1(N9481), .A2(N5281), .ZN(N21624));
    NANDX1 U8753 (.A1(N2621), .A2(n19082), .ZN(n21625));
    INVX1 U8754 (.I(n14358), .ZN(n21626));
    NANDX1 U8755 (.A1(N5880), .A2(N3781), .ZN(n21627));
    INVX1 U8756 (.I(n19029), .ZN(n21628));
    INVX1 U8757 (.I(N8247), .ZN(N21629));
    NOR2X1 U8758 (.A1(n19924), .A2(N5630), .ZN(n21630));
    INVX1 U8759 (.I(N12702), .ZN(N21631));
    NANDX1 U8760 (.A1(N645), .A2(N1764), .ZN(n21632));
    NOR2X1 U8761 (.A1(n20850), .A2(N766), .ZN(n21633));
    NANDX1 U8762 (.A1(N9052), .A2(n19512), .ZN(n21634));
    NOR2X1 U8763 (.A1(N3789), .A2(N10192), .ZN(n21635));
    NANDX1 U8764 (.A1(N9069), .A2(n12889), .ZN(N21636));
    NOR2X1 U8765 (.A1(N6920), .A2(N4152), .ZN(N21637));
    INVX1 U8766 (.I(N2307), .ZN(n21638));
    NANDX1 U8767 (.A1(N3004), .A2(n15906), .ZN(n21639));
    NOR2X1 U8768 (.A1(n14607), .A2(n18694), .ZN(n21640));
    NANDX1 U8769 (.A1(n13300), .A2(n18865), .ZN(N21641));
    NOR2X1 U8770 (.A1(n20543), .A2(N7379), .ZN(n21642));
    NANDX1 U8771 (.A1(N1076), .A2(n18882), .ZN(n21643));
    NOR2X1 U8772 (.A1(n17613), .A2(N1894), .ZN(n21644));
    NANDX1 U8773 (.A1(n15894), .A2(N6806), .ZN(n21645));
    NANDX1 U8774 (.A1(n20628), .A2(n21198), .ZN(n21646));
    NOR2X1 U8775 (.A1(N12286), .A2(N11522), .ZN(n21647));
    INVX1 U8776 (.I(N10980), .ZN(n21648));
    NOR2X1 U8777 (.A1(n16744), .A2(n15552), .ZN(n21649));
    NANDX1 U8778 (.A1(N11419), .A2(N12465), .ZN(n21650));
    NOR2X1 U8779 (.A1(N3424), .A2(N6921), .ZN(n21651));
    NOR2X1 U8780 (.A1(N1058), .A2(N8641), .ZN(n21652));
    INVX1 U8781 (.I(N8437), .ZN(n21653));
    NANDX1 U8782 (.A1(N4438), .A2(N630), .ZN(N21654));
    NANDX1 U8783 (.A1(n16593), .A2(n18295), .ZN(n21655));
    INVX1 U8784 (.I(N5798), .ZN(n21656));
    INVX1 U8785 (.I(n17015), .ZN(n21657));
    INVX1 U8786 (.I(n19609), .ZN(n21658));
    INVX1 U8787 (.I(N12023), .ZN(n21659));
    NOR2X1 U8788 (.A1(n12883), .A2(N1772), .ZN(n21660));
    NANDX1 U8789 (.A1(N8396), .A2(N11865), .ZN(n21661));
    INVX1 U8790 (.I(n14356), .ZN(n21662));
    NOR2X1 U8791 (.A1(N3911), .A2(n17779), .ZN(n21663));
    NANDX1 U8792 (.A1(n13419), .A2(n13379), .ZN(n21664));
    INVX1 U8793 (.I(n16781), .ZN(n21665));
    NOR2X1 U8794 (.A1(n18749), .A2(n21218), .ZN(n21666));
    INVX1 U8795 (.I(n20822), .ZN(n21667));
    NANDX1 U8796 (.A1(n14050), .A2(N1783), .ZN(n21668));
    NANDX1 U8797 (.A1(N12461), .A2(n18797), .ZN(N21669));
    NANDX1 U8798 (.A1(N10839), .A2(N11784), .ZN(n21670));
    INVX1 U8799 (.I(n15280), .ZN(n21671));
    NANDX1 U8800 (.A1(n14677), .A2(N9235), .ZN(N21672));
    NOR2X1 U8801 (.A1(n21084), .A2(N6021), .ZN(n21673));
    NOR2X1 U8802 (.A1(N2953), .A2(N9932), .ZN(n21674));
    INVX1 U8803 (.I(N7514), .ZN(N21675));
    INVX1 U8804 (.I(n14282), .ZN(n21676));
    NOR2X1 U8805 (.A1(n18900), .A2(N9408), .ZN(n21677));
    NANDX1 U8806 (.A1(n13429), .A2(N5163), .ZN(n21678));
    NOR2X1 U8807 (.A1(N8779), .A2(n13754), .ZN(n21679));
    INVX1 U8808 (.I(N4468), .ZN(n21680));
    NOR2X1 U8809 (.A1(N799), .A2(N5351), .ZN(n21681));
    INVX1 U8810 (.I(N7124), .ZN(n21682));
    NANDX1 U8811 (.A1(N4413), .A2(N5102), .ZN(n21683));
    NOR2X1 U8812 (.A1(N8189), .A2(N560), .ZN(N21684));
    NOR2X1 U8813 (.A1(n14210), .A2(N10373), .ZN(N21685));
    NANDX1 U8814 (.A1(n18683), .A2(N5818), .ZN(N21686));
    INVX1 U8815 (.I(n20802), .ZN(N21687));
    NOR2X1 U8816 (.A1(N5132), .A2(n13013), .ZN(N21688));
    NANDX1 U8817 (.A1(N12449), .A2(n20983), .ZN(n21689));
    NOR2X1 U8818 (.A1(n13899), .A2(N3073), .ZN(n21690));
    NANDX1 U8819 (.A1(n17131), .A2(N7540), .ZN(n21691));
    NOR2X1 U8820 (.A1(n17929), .A2(N7433), .ZN(N21692));
    INVX1 U8821 (.I(n19594), .ZN(n21693));
    NOR2X1 U8822 (.A1(N9349), .A2(N3466), .ZN(N21694));
    NANDX1 U8823 (.A1(N12079), .A2(n19797), .ZN(n21695));
    NANDX1 U8824 (.A1(n20830), .A2(N3481), .ZN(n21696));
    INVX1 U8825 (.I(n18282), .ZN(n21697));
    NANDX1 U8826 (.A1(n20581), .A2(N12395), .ZN(N21698));
    INVX1 U8827 (.I(n20254), .ZN(n21699));
    NANDX1 U8828 (.A1(n16444), .A2(N11472), .ZN(n21700));
    NOR2X1 U8829 (.A1(n18967), .A2(n19912), .ZN(n21701));
    NOR2X1 U8830 (.A1(n14013), .A2(n15812), .ZN(n21702));
    NOR2X1 U8831 (.A1(N8585), .A2(N7052), .ZN(n21703));
    NOR2X1 U8832 (.A1(n13521), .A2(N5415), .ZN(n21704));
    NANDX1 U8833 (.A1(n17411), .A2(N3422), .ZN(N21705));
    INVX1 U8834 (.I(N8259), .ZN(n21706));
    INVX1 U8835 (.I(n21186), .ZN(n21707));
    INVX1 U8836 (.I(N10), .ZN(n21708));
    INVX1 U8837 (.I(N4910), .ZN(n21709));
    NANDX1 U8838 (.A1(N3324), .A2(N11847), .ZN(n21710));
    NOR2X1 U8839 (.A1(N2347), .A2(N10565), .ZN(n21711));
    NOR2X1 U8840 (.A1(n13818), .A2(N9036), .ZN(N21712));
    NANDX1 U8841 (.A1(N7041), .A2(N10580), .ZN(n21713));
    INVX1 U8842 (.I(n17394), .ZN(n21714));
    NOR2X1 U8843 (.A1(N874), .A2(n18987), .ZN(N21715));
    NANDX1 U8844 (.A1(n14394), .A2(n18943), .ZN(n21716));
    INVX1 U8845 (.I(N10574), .ZN(N21717));
    NOR2X1 U8846 (.A1(n13016), .A2(n13375), .ZN(n21718));
    NOR2X1 U8847 (.A1(N7514), .A2(n15775), .ZN(N21719));
    INVX1 U8848 (.I(N11487), .ZN(n21720));
    NANDX1 U8849 (.A1(n17295), .A2(n14810), .ZN(N21721));
    INVX1 U8850 (.I(N8080), .ZN(n21722));
    NANDX1 U8851 (.A1(n16407), .A2(N9851), .ZN(n21723));
    NANDX1 U8852 (.A1(N4212), .A2(N3899), .ZN(n21724));
    INVX1 U8853 (.I(N9333), .ZN(n21725));
    NANDX1 U8854 (.A1(N2030), .A2(n18079), .ZN(n21726));
    INVX1 U8855 (.I(n21016), .ZN(N21727));
    NANDX1 U8856 (.A1(N539), .A2(n18728), .ZN(n21728));
    NANDX1 U8857 (.A1(N5655), .A2(n14404), .ZN(n21729));
    INVX1 U8858 (.I(n13571), .ZN(n21730));
    NOR2X1 U8859 (.A1(N2749), .A2(N8115), .ZN(n21731));
    INVX1 U8860 (.I(n14235), .ZN(n21732));
    INVX1 U8861 (.I(n16119), .ZN(n21733));
    NANDX1 U8862 (.A1(N7952), .A2(N2968), .ZN(n21734));
    INVX1 U8863 (.I(N3128), .ZN(n21735));
    NOR2X1 U8864 (.A1(n18337), .A2(N1881), .ZN(n21736));
    INVX1 U8865 (.I(N2973), .ZN(n21737));
    NANDX1 U8866 (.A1(n17760), .A2(N5002), .ZN(n21738));
    INVX1 U8867 (.I(N9363), .ZN(N21739));
    INVX1 U8868 (.I(n19256), .ZN(n21740));
    NOR2X1 U8869 (.A1(n18056), .A2(N6933), .ZN(N21741));
    INVX1 U8870 (.I(N11230), .ZN(N21742));
    NOR2X1 U8871 (.A1(n18210), .A2(n17839), .ZN(n21743));
    INVX1 U8872 (.I(n20866), .ZN(n21744));
    NOR2X1 U8873 (.A1(n13692), .A2(N1745), .ZN(N21745));
    NOR2X1 U8874 (.A1(n16047), .A2(N4238), .ZN(N21746));
    NOR2X1 U8875 (.A1(N8869), .A2(N1907), .ZN(n21747));
    INVX1 U8876 (.I(N517), .ZN(n21748));
    NANDX1 U8877 (.A1(n16762), .A2(n19261), .ZN(n21749));
    NOR2X1 U8878 (.A1(n13291), .A2(n18804), .ZN(n21750));
    INVX1 U8879 (.I(n17196), .ZN(n21751));
    INVX1 U8880 (.I(N10171), .ZN(n21752));
    NANDX1 U8881 (.A1(N9500), .A2(N11646), .ZN(N21753));
    NANDX1 U8882 (.A1(n20729), .A2(n13813), .ZN(n21754));
    INVX1 U8883 (.I(N11879), .ZN(n21755));
    NANDX1 U8884 (.A1(N11976), .A2(N7311), .ZN(n21756));
    NANDX1 U8885 (.A1(N8262), .A2(n13403), .ZN(n21757));
    INVX1 U8886 (.I(N7042), .ZN(N21758));
    NANDX1 U8887 (.A1(N3959), .A2(N8948), .ZN(n21759));
    NOR2X1 U8888 (.A1(n20248), .A2(N12735), .ZN(n21760));
    INVX1 U8889 (.I(n18278), .ZN(n21761));
    INVX1 U8890 (.I(N4641), .ZN(n21762));
    NOR2X1 U8891 (.A1(n13193), .A2(N606), .ZN(n21763));
    INVX1 U8892 (.I(N2133), .ZN(n21764));
    NANDX1 U8893 (.A1(n16794), .A2(N8320), .ZN(n21765));
    INVX1 U8894 (.I(N10834), .ZN(n21766));
    INVX1 U8895 (.I(n17799), .ZN(n21767));
    NOR2X1 U8896 (.A1(n14173), .A2(N3086), .ZN(n21768));
    NOR2X1 U8897 (.A1(n14446), .A2(N5889), .ZN(N21769));
    NANDX1 U8898 (.A1(n14994), .A2(n12930), .ZN(N21770));
    INVX1 U8899 (.I(n13495), .ZN(n21771));
    INVX1 U8900 (.I(N8328), .ZN(N21772));
    NOR2X1 U8901 (.A1(N7924), .A2(n20908), .ZN(N21773));
    NANDX1 U8902 (.A1(N8971), .A2(N4318), .ZN(n21774));
    NANDX1 U8903 (.A1(N933), .A2(n20695), .ZN(n21775));
    INVX1 U8904 (.I(n18837), .ZN(n21776));
    INVX1 U8905 (.I(N11894), .ZN(n21777));
    NOR2X1 U8906 (.A1(N478), .A2(N1498), .ZN(n21778));
    INVX1 U8907 (.I(n18276), .ZN(n21779));
    NANDX1 U8908 (.A1(N10085), .A2(n15903), .ZN(n21780));
    NANDX1 U8909 (.A1(N3300), .A2(N561), .ZN(N21781));
    NOR2X1 U8910 (.A1(N12836), .A2(n13491), .ZN(n21782));
    INVX1 U8911 (.I(n20872), .ZN(n21783));
    NOR2X1 U8912 (.A1(n16595), .A2(N6695), .ZN(n21784));
    INVX1 U8913 (.I(n16272), .ZN(n21785));
    NANDX1 U8914 (.A1(N4343), .A2(n15131), .ZN(N21786));
    NANDX1 U8915 (.A1(n21047), .A2(n14595), .ZN(n21787));
    NANDX1 U8916 (.A1(n13196), .A2(N4156), .ZN(N21788));
    INVX1 U8917 (.I(n13664), .ZN(n21789));
    NOR2X1 U8918 (.A1(N1633), .A2(n15034), .ZN(n21790));
    NANDX1 U8919 (.A1(n14926), .A2(N3888), .ZN(n21791));
    INVX1 U8920 (.I(n15780), .ZN(n21792));
    INVX1 U8921 (.I(N7224), .ZN(n21793));
    NANDX1 U8922 (.A1(n14564), .A2(n15256), .ZN(n21794));
    INVX1 U8923 (.I(N8747), .ZN(N21795));
    NANDX1 U8924 (.A1(N10312), .A2(n15441), .ZN(N21796));
    NOR2X1 U8925 (.A1(N5353), .A2(N5006), .ZN(N21797));
    NOR2X1 U8926 (.A1(n20483), .A2(n19378), .ZN(N21798));
    NOR2X1 U8927 (.A1(N8389), .A2(n13078), .ZN(n21799));
    INVX1 U8928 (.I(N12544), .ZN(n21800));
    NANDX1 U8929 (.A1(n18179), .A2(N6260), .ZN(n21801));
    NANDX1 U8930 (.A1(N6524), .A2(n18251), .ZN(n21802));
    NOR2X1 U8931 (.A1(N4953), .A2(n19456), .ZN(n21803));
    NOR2X1 U8932 (.A1(N6681), .A2(N5449), .ZN(n21804));
    NANDX1 U8933 (.A1(n15787), .A2(n15247), .ZN(n21805));
    NANDX1 U8934 (.A1(N3303), .A2(n17951), .ZN(n21806));
    NOR2X1 U8935 (.A1(n18744), .A2(n16028), .ZN(n21807));
    INVX1 U8936 (.I(n18291), .ZN(n21808));
    NANDX1 U8937 (.A1(N12342), .A2(n16438), .ZN(n21809));
    INVX1 U8938 (.I(n20730), .ZN(n21810));
    NANDX1 U8939 (.A1(N3367), .A2(N6585), .ZN(n21811));
    INVX1 U8940 (.I(n16087), .ZN(n21812));
    NANDX1 U8941 (.A1(n14510), .A2(N1380), .ZN(N21813));
    INVX1 U8942 (.I(N12134), .ZN(n21814));
    INVX1 U8943 (.I(N2631), .ZN(n21815));
    NANDX1 U8944 (.A1(n13012), .A2(N2622), .ZN(n21816));
    NANDX1 U8945 (.A1(N2110), .A2(n17868), .ZN(n21817));
    NOR2X1 U8946 (.A1(N5413), .A2(n14588), .ZN(n21818));
    INVX1 U8947 (.I(n18698), .ZN(n21819));
    INVX1 U8948 (.I(N11100), .ZN(n21820));
    NOR2X1 U8949 (.A1(N11459), .A2(N2212), .ZN(n21821));
    NANDX1 U8950 (.A1(N10310), .A2(N1711), .ZN(n21822));
    INVX1 U8951 (.I(N8218), .ZN(n21823));
    NOR2X1 U8952 (.A1(n13455), .A2(N3074), .ZN(n21824));
    INVX1 U8953 (.I(N6735), .ZN(n21825));
    INVX1 U8954 (.I(n14629), .ZN(n21826));
    NOR2X1 U8955 (.A1(N10784), .A2(n17259), .ZN(n21827));
    NOR2X1 U8956 (.A1(n18337), .A2(n14422), .ZN(n21828));
    INVX1 U8957 (.I(n20447), .ZN(n21829));
    NOR2X1 U8958 (.A1(N10547), .A2(n20401), .ZN(n21830));
    NOR2X1 U8959 (.A1(N3099), .A2(n17868), .ZN(n21831));
    NOR2X1 U8960 (.A1(N8741), .A2(N1479), .ZN(n21832));
    INVX1 U8961 (.I(N10952), .ZN(N21833));
    INVX1 U8962 (.I(n19195), .ZN(n21834));
    INVX1 U8963 (.I(N4401), .ZN(N21835));
    NANDX1 U8964 (.A1(N10041), .A2(N12397), .ZN(n21836));
    NOR2X1 U8965 (.A1(n20264), .A2(n19131), .ZN(n21837));
    INVX1 U8966 (.I(n13662), .ZN(n21838));
    NOR2X1 U8967 (.A1(n19032), .A2(N4232), .ZN(n21839));
    NOR2X1 U8968 (.A1(N10680), .A2(n18654), .ZN(n21840));
    NOR2X1 U8969 (.A1(N9896), .A2(N8482), .ZN(n21841));
    NOR2X1 U8970 (.A1(N3608), .A2(N7440), .ZN(N21842));
    INVX1 U8971 (.I(n16017), .ZN(n21843));
    INVX1 U8972 (.I(N2538), .ZN(n21844));
    INVX1 U8973 (.I(n13752), .ZN(n21845));
    NOR2X1 U8974 (.A1(n19021), .A2(N11716), .ZN(n21846));
    NOR2X1 U8975 (.A1(N2191), .A2(N12439), .ZN(n21847));
    NOR2X1 U8976 (.A1(N9130), .A2(n16235), .ZN(n21848));
    NANDX1 U8977 (.A1(N1572), .A2(N3253), .ZN(n21849));
    NANDX1 U8978 (.A1(n12882), .A2(n16826), .ZN(n21850));
    NANDX1 U8979 (.A1(n15220), .A2(N6276), .ZN(n21851));
    INVX1 U8980 (.I(N830), .ZN(N21852));
    NOR2X1 U8981 (.A1(N10501), .A2(n18217), .ZN(n21853));
    NANDX1 U8982 (.A1(N12482), .A2(N12014), .ZN(n21854));
    INVX1 U8983 (.I(n17349), .ZN(n21855));
    NOR2X1 U8984 (.A1(n21144), .A2(N4412), .ZN(n21856));
    NANDX1 U8985 (.A1(n13476), .A2(n16128), .ZN(N21857));
    INVX1 U8986 (.I(N10209), .ZN(n21858));
    NOR2X1 U8987 (.A1(N9712), .A2(n19338), .ZN(n21859));
    INVX1 U8988 (.I(N7331), .ZN(N21860));
    INVX1 U8989 (.I(n15907), .ZN(n21861));
    INVX1 U8990 (.I(N7103), .ZN(N21862));
    NANDX1 U8991 (.A1(N1977), .A2(n16864), .ZN(n21863));
    INVX1 U8992 (.I(N3995), .ZN(N21864));
    NOR2X1 U8993 (.A1(N12116), .A2(n14495), .ZN(n21865));
    NOR2X1 U8994 (.A1(n20978), .A2(N5747), .ZN(n21866));
    INVX1 U8995 (.I(N3397), .ZN(n21867));
    NOR2X1 U8996 (.A1(N9097), .A2(n19082), .ZN(N21868));
    NANDX1 U8997 (.A1(N4989), .A2(N11327), .ZN(N21869));
    NANDX1 U8998 (.A1(n16114), .A2(n16077), .ZN(n21870));
    NANDX1 U8999 (.A1(n20368), .A2(n14184), .ZN(N21871));
    NANDX1 U9000 (.A1(N6468), .A2(N8405), .ZN(n21872));
    NANDX1 U9001 (.A1(n14163), .A2(n15507), .ZN(n21873));
    NOR2X1 U9002 (.A1(n16139), .A2(N11140), .ZN(n21874));
    INVX1 U9003 (.I(n20133), .ZN(n21875));
    NOR2X1 U9004 (.A1(N8112), .A2(N7940), .ZN(N21876));
    NOR2X1 U9005 (.A1(N7859), .A2(N8228), .ZN(n21877));
    NOR2X1 U9006 (.A1(N5797), .A2(n20406), .ZN(n21878));
    NOR2X1 U9007 (.A1(N3648), .A2(n15765), .ZN(n21879));
    NOR2X1 U9008 (.A1(N9517), .A2(N564), .ZN(n21880));
    NANDX1 U9009 (.A1(N4363), .A2(N8470), .ZN(n21881));
    INVX1 U9010 (.I(n13089), .ZN(N21882));
    INVX1 U9011 (.I(n15026), .ZN(n21883));
    NOR2X1 U9012 (.A1(N12120), .A2(N2500), .ZN(n21884));
    NOR2X1 U9013 (.A1(N1255), .A2(n18638), .ZN(N21885));
    NOR2X1 U9014 (.A1(n18480), .A2(N12083), .ZN(n21886));
    INVX1 U9015 (.I(N5361), .ZN(n21887));
    NOR2X1 U9016 (.A1(n13730), .A2(N7762), .ZN(n21888));
    INVX1 U9017 (.I(N3870), .ZN(N21889));
    INVX1 U9018 (.I(N736), .ZN(n21890));
    INVX1 U9019 (.I(N11748), .ZN(N21891));
    NANDX1 U9020 (.A1(N1871), .A2(n15806), .ZN(n21892));
    NANDX1 U9021 (.A1(n16750), .A2(n14710), .ZN(n21893));
    INVX1 U9022 (.I(N4078), .ZN(n21894));
    NANDX1 U9023 (.A1(N1185), .A2(n13645), .ZN(n21895));
    NANDX1 U9024 (.A1(N7847), .A2(n16145), .ZN(n21896));
    INVX1 U9025 (.I(N9101), .ZN(n21897));
    NANDX1 U9026 (.A1(N6444), .A2(N892), .ZN(N21898));
    INVX1 U9027 (.I(N8808), .ZN(n21899));
    NANDX1 U9028 (.A1(n13509), .A2(N1307), .ZN(n21900));
    NOR2X1 U9029 (.A1(n15069), .A2(N5176), .ZN(n21901));
    INVX1 U9030 (.I(n15804), .ZN(N21902));
    NANDX1 U9031 (.A1(N7172), .A2(N5616), .ZN(n21903));
    NOR2X1 U9032 (.A1(N1747), .A2(N1448), .ZN(n21904));
    NANDX1 U9033 (.A1(N10999), .A2(n16064), .ZN(n21905));
    NOR2X1 U9034 (.A1(n17566), .A2(n17248), .ZN(n21906));
    NOR2X1 U9035 (.A1(n13480), .A2(n19636), .ZN(n21907));
    INVX1 U9036 (.I(N3931), .ZN(N21908));
    INVX1 U9037 (.I(N4567), .ZN(N21909));
    INVX1 U9038 (.I(N8398), .ZN(n21910));
    NANDX1 U9039 (.A1(n13723), .A2(N9192), .ZN(n21911));
    NOR2X1 U9040 (.A1(n15030), .A2(N12289), .ZN(n21912));
    INVX1 U9041 (.I(n14747), .ZN(n21913));
    NANDX1 U9042 (.A1(N10289), .A2(n17569), .ZN(N21914));
    NANDX1 U9043 (.A1(n15904), .A2(N1031), .ZN(n21915));
    INVX1 U9044 (.I(N11893), .ZN(N21916));
    INVX1 U9045 (.I(n16713), .ZN(n21917));
    NANDX1 U9046 (.A1(N10386), .A2(n13049), .ZN(N21918));
    INVX1 U9047 (.I(N11945), .ZN(n21919));
    NANDX1 U9048 (.A1(n16921), .A2(N8417), .ZN(n21920));
    NANDX1 U9049 (.A1(N3197), .A2(n12983), .ZN(n21921));
    INVX1 U9050 (.I(N6136), .ZN(n21922));
    NANDX1 U9051 (.A1(N1178), .A2(N9869), .ZN(n21923));
    NANDX1 U9052 (.A1(n16207), .A2(N927), .ZN(n21924));
    NANDX1 U9053 (.A1(N4266), .A2(N3181), .ZN(n21925));
    INVX1 U9054 (.I(n16376), .ZN(n21926));
    NANDX1 U9055 (.A1(N814), .A2(N11949), .ZN(n21927));
    INVX1 U9056 (.I(N12707), .ZN(n21928));
    NANDX1 U9057 (.A1(n13804), .A2(n19432), .ZN(n21929));
    INVX1 U9058 (.I(N5622), .ZN(N21930));
    INVX1 U9059 (.I(n19146), .ZN(n21931));
    INVX1 U9060 (.I(N6950), .ZN(n21932));
    INVX1 U9061 (.I(N3773), .ZN(n21933));
    NOR2X1 U9062 (.A1(n19315), .A2(N12458), .ZN(n21934));
    NOR2X1 U9063 (.A1(N9121), .A2(n13635), .ZN(N21935));
    NOR2X1 U9064 (.A1(N5031), .A2(N3154), .ZN(n21936));
    INVX1 U9065 (.I(n16655), .ZN(n21937));
    NOR2X1 U9066 (.A1(n13881), .A2(N1566), .ZN(n21938));
    NOR2X1 U9067 (.A1(N5258), .A2(n18151), .ZN(n21939));
    NOR2X1 U9068 (.A1(N2349), .A2(N9627), .ZN(n21940));
    NOR2X1 U9069 (.A1(n16152), .A2(N2371), .ZN(n21941));
    NOR2X1 U9070 (.A1(n16316), .A2(n13629), .ZN(n21942));
    INVX1 U9071 (.I(n16318), .ZN(N21943));
    NANDX1 U9072 (.A1(n17317), .A2(n20090), .ZN(n21944));
    INVX1 U9073 (.I(N9943), .ZN(n21945));
    NOR2X1 U9074 (.A1(N9399), .A2(n13605), .ZN(n21946));
    NOR2X1 U9075 (.A1(n19173), .A2(n13177), .ZN(n21947));
    NANDX1 U9076 (.A1(N8643), .A2(N8602), .ZN(n21948));
    INVX1 U9077 (.I(N1294), .ZN(n21949));
    NANDX1 U9078 (.A1(N10796), .A2(N6551), .ZN(n21950));
    NANDX1 U9079 (.A1(n14392), .A2(N8899), .ZN(n21951));
    NOR2X1 U9080 (.A1(n20261), .A2(n19592), .ZN(n21952));
    NANDX1 U9081 (.A1(N12101), .A2(n14677), .ZN(n21953));
    INVX1 U9082 (.I(n17628), .ZN(N21954));
    NOR2X1 U9083 (.A1(N10228), .A2(N8256), .ZN(n21955));
    INVX1 U9084 (.I(N8804), .ZN(n21956));
    INVX1 U9085 (.I(N3567), .ZN(N21957));
    INVX1 U9086 (.I(N10573), .ZN(N21958));
    INVX1 U9087 (.I(N10687), .ZN(N21959));
    NANDX1 U9088 (.A1(n13560), .A2(n19330), .ZN(n21960));
    NANDX1 U9089 (.A1(N6020), .A2(n20623), .ZN(n21961));
    INVX1 U9090 (.I(n16815), .ZN(n21962));
    NOR2X1 U9091 (.A1(N11999), .A2(N9976), .ZN(n21963));
    NANDX1 U9092 (.A1(n17796), .A2(N3548), .ZN(N21964));
    INVX1 U9093 (.I(N4733), .ZN(n21965));
    NANDX1 U9094 (.A1(N11505), .A2(n15613), .ZN(N21966));
    NOR2X1 U9095 (.A1(n15811), .A2(N4610), .ZN(n21967));
    NANDX1 U9096 (.A1(n13518), .A2(N7955), .ZN(n21968));
    NANDX1 U9097 (.A1(n17084), .A2(n20699), .ZN(n21969));
    NOR2X1 U9098 (.A1(n13455), .A2(N4698), .ZN(n21970));
    NANDX1 U9099 (.A1(N5784), .A2(n18569), .ZN(N21971));
    NOR2X1 U9100 (.A1(N11803), .A2(N12503), .ZN(n21972));
    NOR2X1 U9101 (.A1(N1930), .A2(n12987), .ZN(n21973));
    NANDX1 U9102 (.A1(N11905), .A2(N11453), .ZN(n21974));
    NOR2X1 U9103 (.A1(N9995), .A2(n13738), .ZN(n21975));
    INVX1 U9104 (.I(n20184), .ZN(n21976));
    INVX1 U9105 (.I(N11009), .ZN(n21977));
    NOR2X1 U9106 (.A1(n14364), .A2(N10160), .ZN(N21978));
    INVX1 U9107 (.I(N1194), .ZN(n21979));
    NOR2X1 U9108 (.A1(N5505), .A2(n18277), .ZN(n21980));
    NANDX1 U9109 (.A1(N1199), .A2(N10502), .ZN(n21981));
    NOR2X1 U9110 (.A1(N9727), .A2(N10827), .ZN(N21982));
    INVX1 U9111 (.I(N8144), .ZN(N21983));
    NANDX1 U9112 (.A1(n21204), .A2(N11474), .ZN(n21984));
    NOR2X1 U9113 (.A1(n12960), .A2(N5572), .ZN(n21985));
    NOR2X1 U9114 (.A1(n18954), .A2(n17465), .ZN(n21986));
    NOR2X1 U9115 (.A1(N11461), .A2(N12861), .ZN(N21987));
    NOR2X1 U9116 (.A1(N4557), .A2(n18411), .ZN(n21988));
    NANDX1 U9117 (.A1(n13462), .A2(N7340), .ZN(N21989));
    NOR2X1 U9118 (.A1(n14655), .A2(n19996), .ZN(n21990));
    NANDX1 U9119 (.A1(N11702), .A2(N10890), .ZN(N21991));
    INVX1 U9120 (.I(n16745), .ZN(n21992));
    INVX1 U9121 (.I(N2239), .ZN(n21993));
    NANDX1 U9122 (.A1(N9724), .A2(N4925), .ZN(N21994));
    INVX1 U9123 (.I(N9697), .ZN(N21995));
    NANDX1 U9124 (.A1(n15924), .A2(n17198), .ZN(N21996));
    NANDX1 U9125 (.A1(n20241), .A2(n14921), .ZN(n21997));
    NANDX1 U9126 (.A1(N7863), .A2(n20923), .ZN(N21998));
    INVX1 U9127 (.I(n21127), .ZN(N21999));
    NOR2X1 U9128 (.A1(N1556), .A2(n13243), .ZN(n22000));
    NANDX1 U9129 (.A1(N3438), .A2(N4511), .ZN(n22001));
    NANDX1 U9130 (.A1(N2203), .A2(n17055), .ZN(n22002));
    NOR2X1 U9131 (.A1(N7634), .A2(N9568), .ZN(N22003));
    NANDX1 U9132 (.A1(N3198), .A2(N6348), .ZN(n22004));
    NANDX1 U9133 (.A1(n12921), .A2(N11272), .ZN(n22005));
    NANDX1 U9134 (.A1(n17159), .A2(N981), .ZN(n22006));
    NANDX1 U9135 (.A1(n13126), .A2(n17491), .ZN(n22007));
    NANDX1 U9136 (.A1(N1358), .A2(n14464), .ZN(N22008));
    INVX1 U9137 (.I(N1050), .ZN(n22009));
    NOR2X1 U9138 (.A1(n16917), .A2(n21071), .ZN(n22010));
    NOR2X1 U9139 (.A1(N8929), .A2(N12093), .ZN(n22011));
    NOR2X1 U9140 (.A1(N7982), .A2(N12311), .ZN(n22012));
    NANDX1 U9141 (.A1(N3806), .A2(N3001), .ZN(n22013));
    INVX1 U9142 (.I(N7915), .ZN(N22014));
    NANDX1 U9143 (.A1(n15031), .A2(n14263), .ZN(n22015));
    NOR2X1 U9144 (.A1(N1263), .A2(n20076), .ZN(n22016));
    NANDX1 U9145 (.A1(n18421), .A2(n21057), .ZN(n22017));
    INVX1 U9146 (.I(N4858), .ZN(N22018));
    NOR2X1 U9147 (.A1(N132), .A2(N6215), .ZN(N22019));
    NANDX1 U9148 (.A1(n17151), .A2(N7265), .ZN(n22020));
    NANDX1 U9149 (.A1(N7379), .A2(N1647), .ZN(n22021));
    NANDX1 U9150 (.A1(N10850), .A2(n13739), .ZN(n22022));
    NANDX1 U9151 (.A1(n18831), .A2(N4819), .ZN(N22023));
    INVX1 U9152 (.I(N1406), .ZN(N22024));
    NANDX1 U9153 (.A1(n13836), .A2(N9321), .ZN(n22025));
    INVX1 U9154 (.I(N7637), .ZN(N22026));
    NOR2X1 U9155 (.A1(n20026), .A2(N3441), .ZN(n22027));
    NOR2X1 U9156 (.A1(N853), .A2(N632), .ZN(n22028));
    INVX1 U9157 (.I(N7599), .ZN(N22029));
    INVX1 U9158 (.I(N1967), .ZN(n22030));
    INVX1 U9159 (.I(N6246), .ZN(n22031));
    NOR2X1 U9160 (.A1(n19423), .A2(N8052), .ZN(N22032));
    NOR2X1 U9161 (.A1(N113), .A2(N9698), .ZN(n22033));
    NANDX1 U9162 (.A1(N10962), .A2(n17978), .ZN(n22034));
    NOR2X1 U9163 (.A1(N8562), .A2(N1566), .ZN(n22035));
    NOR2X1 U9164 (.A1(N9968), .A2(n19699), .ZN(n22036));
    NANDX1 U9165 (.A1(n19288), .A2(n16119), .ZN(N22037));
    NANDX1 U9166 (.A1(n16182), .A2(n14914), .ZN(n22038));
    INVX1 U9167 (.I(N6463), .ZN(n22039));
    NOR2X1 U9168 (.A1(n14533), .A2(n17801), .ZN(N22040));
    NANDX1 U9169 (.A1(N9106), .A2(n19767), .ZN(n22041));
    INVX1 U9170 (.I(n15351), .ZN(n22042));
    NOR2X1 U9171 (.A1(n12913), .A2(N2172), .ZN(N22043));
    NANDX1 U9172 (.A1(n13025), .A2(N6411), .ZN(n22044));
    NOR2X1 U9173 (.A1(N2757), .A2(N3158), .ZN(n22045));
    INVX1 U9174 (.I(N11318), .ZN(n22046));
    NANDX1 U9175 (.A1(N12058), .A2(n15827), .ZN(n22047));
    INVX1 U9176 (.I(n20341), .ZN(n22048));
    NOR2X1 U9177 (.A1(n13851), .A2(N9572), .ZN(N22049));
    INVX1 U9178 (.I(N2077), .ZN(n22050));
    NOR2X1 U9179 (.A1(N4382), .A2(N12385), .ZN(n22051));
    INVX1 U9180 (.I(N952), .ZN(N22052));
    NANDX1 U9181 (.A1(N4651), .A2(n20718), .ZN(N22053));
    NOR2X1 U9182 (.A1(n14543), .A2(n15395), .ZN(n22054));
    INVX1 U9183 (.I(N11256), .ZN(n22055));
    INVX1 U9184 (.I(N1800), .ZN(n22056));
    NOR2X1 U9185 (.A1(N7390), .A2(n20328), .ZN(n22057));
    NOR2X1 U9186 (.A1(n19542), .A2(N10415), .ZN(N22058));
    NOR2X1 U9187 (.A1(N4912), .A2(n20784), .ZN(N22059));
    INVX1 U9188 (.I(n19794), .ZN(N22060));
    NOR2X1 U9189 (.A1(N4983), .A2(N8136), .ZN(n22061));
    INVX1 U9190 (.I(N1601), .ZN(n22062));
    INVX1 U9191 (.I(N10279), .ZN(n22063));
    INVX1 U9192 (.I(N466), .ZN(N22064));
    NANDX1 U9193 (.A1(N12129), .A2(n20889), .ZN(n22065));
    INVX1 U9194 (.I(N9222), .ZN(N22066));
    NOR2X1 U9195 (.A1(n15195), .A2(n13768), .ZN(N22067));
    NOR2X1 U9196 (.A1(n18650), .A2(n15567), .ZN(N22068));
    NOR2X1 U9197 (.A1(N4810), .A2(N9206), .ZN(N22069));
    INVX1 U9198 (.I(n18893), .ZN(N22070));
    NANDX1 U9199 (.A1(N9426), .A2(n18346), .ZN(N22071));
    NOR2X1 U9200 (.A1(N557), .A2(n16910), .ZN(n22072));
    NANDX1 U9201 (.A1(N81), .A2(N3815), .ZN(N22073));
    NOR2X1 U9202 (.A1(N1681), .A2(n14193), .ZN(n22074));
    INVX1 U9203 (.I(N10207), .ZN(n22075));
    INVX1 U9204 (.I(N11494), .ZN(N22076));
    INVX1 U9205 (.I(n14316), .ZN(N22077));
    NOR2X1 U9206 (.A1(N4869), .A2(N1829), .ZN(n22078));
    NANDX1 U9207 (.A1(n18636), .A2(N597), .ZN(n22079));
    NANDX1 U9208 (.A1(N7515), .A2(n17030), .ZN(N22080));
    NANDX1 U9209 (.A1(n16720), .A2(N6368), .ZN(N22081));
    NANDX1 U9210 (.A1(N9652), .A2(N10335), .ZN(n22082));
    NANDX1 U9211 (.A1(N2137), .A2(N5434), .ZN(n22083));
    INVX1 U9212 (.I(n18373), .ZN(N22084));
    NANDX1 U9213 (.A1(N6614), .A2(n19275), .ZN(n22085));
    NANDX1 U9214 (.A1(n15348), .A2(N3768), .ZN(n22086));
    NANDX1 U9215 (.A1(N3318), .A2(n15261), .ZN(n22087));
    NANDX1 U9216 (.A1(N12175), .A2(N5325), .ZN(n22088));
    INVX1 U9217 (.I(n14003), .ZN(n22089));
    NOR2X1 U9218 (.A1(n20178), .A2(n14599), .ZN(n22090));
    INVX1 U9219 (.I(N1004), .ZN(n22091));
    INVX1 U9220 (.I(n20145), .ZN(n22092));
    NANDX1 U9221 (.A1(N5850), .A2(n14378), .ZN(n22093));
    INVX1 U9222 (.I(n16185), .ZN(n22094));
    INVX1 U9223 (.I(n18595), .ZN(n22095));
    INVX1 U9224 (.I(N3068), .ZN(n22096));
    NANDX1 U9225 (.A1(N443), .A2(N4223), .ZN(n22097));
    NOR2X1 U9226 (.A1(n17951), .A2(n19571), .ZN(n22098));
    INVX1 U9227 (.I(N3206), .ZN(n22099));
    NOR2X1 U9228 (.A1(N6121), .A2(N5337), .ZN(N22100));
    NANDX1 U9229 (.A1(N5987), .A2(N6879), .ZN(n22101));
    INVX1 U9230 (.I(N11111), .ZN(N22102));
    NOR2X1 U9231 (.A1(N10287), .A2(N7997), .ZN(n22103));
    INVX1 U9232 (.I(N9769), .ZN(N22104));
    NOR2X1 U9233 (.A1(n13635), .A2(n15619), .ZN(N22105));
    NANDX1 U9234 (.A1(N8863), .A2(N5115), .ZN(n22106));
    NOR2X1 U9235 (.A1(N6228), .A2(N44), .ZN(n22107));
    INVX1 U9236 (.I(n16506), .ZN(n22108));
    INVX1 U9237 (.I(N12471), .ZN(n22109));
    NOR2X1 U9238 (.A1(n12979), .A2(N5353), .ZN(n22110));
    INVX1 U9239 (.I(n16184), .ZN(n22111));
    NANDX1 U9240 (.A1(N10894), .A2(n16062), .ZN(n22112));
    INVX1 U9241 (.I(n16880), .ZN(n22113));
    NANDX1 U9242 (.A1(N11071), .A2(N6761), .ZN(n22114));
    INVX1 U9243 (.I(n15900), .ZN(n22115));
    INVX1 U9244 (.I(n19219), .ZN(N22116));
    NOR2X1 U9245 (.A1(n16209), .A2(N11624), .ZN(N22117));
    NANDX1 U9246 (.A1(N10808), .A2(n15028), .ZN(n22118));
    NANDX1 U9247 (.A1(N216), .A2(n15797), .ZN(n22119));
    NANDX1 U9248 (.A1(N8464), .A2(N11073), .ZN(n22120));
    NOR2X1 U9249 (.A1(n15476), .A2(N9213), .ZN(N22121));
    NANDX1 U9250 (.A1(n20828), .A2(n13986), .ZN(n22122));
    NANDX1 U9251 (.A1(N1149), .A2(N3649), .ZN(N22123));
    NOR2X1 U9252 (.A1(N11073), .A2(n20528), .ZN(n22124));
    NOR2X1 U9253 (.A1(N914), .A2(N600), .ZN(n22125));
    INVX1 U9254 (.I(n16813), .ZN(N22126));
    NANDX1 U9255 (.A1(N2946), .A2(n15792), .ZN(n22127));
    NANDX1 U9256 (.A1(N9111), .A2(n14618), .ZN(n22128));
    INVX1 U9257 (.I(N2908), .ZN(n22129));
    NANDX1 U9258 (.A1(N4983), .A2(n18705), .ZN(n22130));
    INVX1 U9259 (.I(N7988), .ZN(n22131));
    NANDX1 U9260 (.A1(n20948), .A2(N2233), .ZN(N22132));
    NOR2X1 U9261 (.A1(N790), .A2(n17602), .ZN(n22133));
    NANDX1 U9262 (.A1(N12587), .A2(n18750), .ZN(n22134));
    NOR2X1 U9263 (.A1(N3443), .A2(N3134), .ZN(n22135));
    NOR2X1 U9264 (.A1(N6323), .A2(N4047), .ZN(n22136));
    NOR2X1 U9265 (.A1(N11280), .A2(n15401), .ZN(n22137));
    NOR2X1 U9266 (.A1(n14225), .A2(N9963), .ZN(n22138));
    INVX1 U9267 (.I(N2105), .ZN(n22139));
    INVX1 U9268 (.I(N11767), .ZN(N22140));
    INVX1 U9269 (.I(N5532), .ZN(n22141));
    NOR2X1 U9270 (.A1(n18258), .A2(N6239), .ZN(N22142));
    NANDX1 U9271 (.A1(n15888), .A2(N498), .ZN(n22143));
    NANDX1 U9272 (.A1(N1501), .A2(n17059), .ZN(n22144));
    NANDX1 U9273 (.A1(N1098), .A2(N8415), .ZN(N22145));
    NANDX1 U9274 (.A1(n20116), .A2(N6400), .ZN(n22146));
    NANDX1 U9275 (.A1(n17201), .A2(N12722), .ZN(N22147));
    NANDX1 U9276 (.A1(N9427), .A2(n18543), .ZN(n22148));
    NANDX1 U9277 (.A1(N11551), .A2(N11537), .ZN(n22149));
    NOR2X1 U9278 (.A1(n13093), .A2(N8183), .ZN(N22150));
    INVX1 U9279 (.I(N3629), .ZN(n22151));
    NOR2X1 U9280 (.A1(n13159), .A2(N9461), .ZN(n22152));
    INVX1 U9281 (.I(n19397), .ZN(n22153));
    NOR2X1 U9282 (.A1(n15194), .A2(n14437), .ZN(n22154));
    INVX1 U9283 (.I(N11236), .ZN(n22155));
    NANDX1 U9284 (.A1(n19607), .A2(N12333), .ZN(n22156));
    INVX1 U9285 (.I(N2860), .ZN(N22157));
    NOR2X1 U9286 (.A1(N3849), .A2(N5018), .ZN(n22158));
    INVX1 U9287 (.I(N11112), .ZN(n22159));
    NANDX1 U9288 (.A1(N5699), .A2(N8425), .ZN(n22160));
    INVX1 U9289 (.I(n17249), .ZN(N22161));
    INVX1 U9290 (.I(n15876), .ZN(n22162));
    NOR2X1 U9291 (.A1(N1456), .A2(N7731), .ZN(n22163));
    INVX1 U9292 (.I(N3734), .ZN(n22164));
    NANDX1 U9293 (.A1(N11283), .A2(n18811), .ZN(n22165));
    NANDX1 U9294 (.A1(n13332), .A2(N7316), .ZN(n22166));
    NANDX1 U9295 (.A1(N4744), .A2(n18551), .ZN(N22167));
    INVX1 U9296 (.I(N3120), .ZN(n22168));
    INVX1 U9297 (.I(n14517), .ZN(n22169));
    INVX1 U9298 (.I(N9955), .ZN(n22170));
    INVX1 U9299 (.I(N81), .ZN(n22171));
    INVX1 U9300 (.I(n18560), .ZN(n22172));
    NOR2X1 U9301 (.A1(N6467), .A2(N5754), .ZN(N22173));
    INVX1 U9302 (.I(n18257), .ZN(n22174));
    NOR2X1 U9303 (.A1(n16945), .A2(N680), .ZN(n22175));
    NANDX1 U9304 (.A1(n19217), .A2(N2502), .ZN(n22176));
    NANDX1 U9305 (.A1(n18875), .A2(N8327), .ZN(N22177));
    NANDX1 U9306 (.A1(N11241), .A2(N428), .ZN(n22178));
    INVX1 U9307 (.I(N12586), .ZN(n22179));
    INVX1 U9308 (.I(n16745), .ZN(n22180));
    NOR2X1 U9309 (.A1(N2833), .A2(n15482), .ZN(n22181));
    INVX1 U9310 (.I(n19126), .ZN(n22182));
    NOR2X1 U9311 (.A1(N3699), .A2(n19206), .ZN(N22183));
    INVX1 U9312 (.I(N1028), .ZN(n22184));
    NOR2X1 U9313 (.A1(N11441), .A2(N1324), .ZN(N22185));
    INVX1 U9314 (.I(N8467), .ZN(N22186));
    NOR2X1 U9315 (.A1(N10917), .A2(N9146), .ZN(n22187));
    INVX1 U9316 (.I(N8903), .ZN(N22188));
    NANDX1 U9317 (.A1(n14757), .A2(N1089), .ZN(n22189));
    INVX1 U9318 (.I(N177), .ZN(n22190));
    NANDX1 U9319 (.A1(N9485), .A2(n14143), .ZN(N22191));
    INVX1 U9320 (.I(N9198), .ZN(n22192));
    NOR2X1 U9321 (.A1(N1190), .A2(N6573), .ZN(n22193));
    NANDX1 U9322 (.A1(n13212), .A2(N4468), .ZN(n22194));
    INVX1 U9323 (.I(n16910), .ZN(n22195));
    NANDX1 U9324 (.A1(N7631), .A2(N12480), .ZN(n22196));
    INVX1 U9325 (.I(n13613), .ZN(N22197));
    NANDX1 U9326 (.A1(N10548), .A2(N850), .ZN(n22198));
    INVX1 U9327 (.I(n16006), .ZN(N22199));
    NOR2X1 U9328 (.A1(n19236), .A2(n19450), .ZN(n22200));
    INVX1 U9329 (.I(N7304), .ZN(n22201));
    NOR2X1 U9330 (.A1(N4011), .A2(N7480), .ZN(n22202));
    NOR2X1 U9331 (.A1(n13496), .A2(N393), .ZN(n22203));
    NOR2X1 U9332 (.A1(N1463), .A2(n20364), .ZN(N22204));
    NANDX1 U9333 (.A1(N2577), .A2(n18814), .ZN(n22205));
    NOR2X1 U9334 (.A1(N7044), .A2(n16013), .ZN(N22206));
    INVX1 U9335 (.I(n19800), .ZN(n22207));
    INVX1 U9336 (.I(N10590), .ZN(n22208));
    INVX1 U9337 (.I(N10568), .ZN(n22209));
    INVX1 U9338 (.I(n20235), .ZN(n22210));
    NANDX1 U9339 (.A1(N11253), .A2(N9553), .ZN(n22211));
    NANDX1 U9340 (.A1(N3800), .A2(N7772), .ZN(n22212));
    INVX1 U9341 (.I(N11103), .ZN(N22213));
    INVX1 U9342 (.I(N9459), .ZN(n22214));
    NOR2X1 U9343 (.A1(N2342), .A2(n17496), .ZN(N22215));
    NOR2X1 U9344 (.A1(n17059), .A2(n18959), .ZN(n22216));
    NANDX1 U9345 (.A1(N11736), .A2(N305), .ZN(N22217));
    NOR2X1 U9346 (.A1(n14167), .A2(N1891), .ZN(N22218));
    NOR2X1 U9347 (.A1(N12277), .A2(n16232), .ZN(n22219));
    NOR2X1 U9348 (.A1(n17408), .A2(N4689), .ZN(n22220));
    INVX1 U9349 (.I(N9653), .ZN(N22221));
    NOR2X1 U9350 (.A1(n13036), .A2(n20905), .ZN(N22222));
    INVX1 U9351 (.I(N7759), .ZN(N22223));
    NOR2X1 U9352 (.A1(N10101), .A2(n13207), .ZN(n22224));
    NOR2X1 U9353 (.A1(N11722), .A2(n17207), .ZN(N22225));
    NOR2X1 U9354 (.A1(n14063), .A2(n13473), .ZN(n22226));
    NOR2X1 U9355 (.A1(N9892), .A2(N5743), .ZN(n22227));
    NANDX1 U9356 (.A1(n16169), .A2(N589), .ZN(n22228));
    NANDX1 U9357 (.A1(N9105), .A2(n18251), .ZN(n22229));
    INVX1 U9358 (.I(n15923), .ZN(n22230));
    NANDX1 U9359 (.A1(N6786), .A2(N12100), .ZN(n22231));
    NANDX1 U9360 (.A1(N8405), .A2(N522), .ZN(n22232));
    INVX1 U9361 (.I(N211), .ZN(n22233));
    NANDX1 U9362 (.A1(n13047), .A2(N7969), .ZN(N22234));
    NANDX1 U9363 (.A1(N1918), .A2(n15717), .ZN(N22235));
    NANDX1 U9364 (.A1(N8181), .A2(N6235), .ZN(n22236));
    NANDX1 U9365 (.A1(N1014), .A2(n19707), .ZN(N22237));
    NANDX1 U9366 (.A1(N5447), .A2(n19991), .ZN(n22238));
    NOR2X1 U9367 (.A1(n16157), .A2(n20580), .ZN(n22239));
    NANDX1 U9368 (.A1(n19804), .A2(N12142), .ZN(N22240));
    NOR2X1 U9369 (.A1(n14496), .A2(N4164), .ZN(N22241));
    NOR2X1 U9370 (.A1(N5366), .A2(n16647), .ZN(n22242));
    NANDX1 U9371 (.A1(N5887), .A2(N676), .ZN(N22243));
    NOR2X1 U9372 (.A1(N625), .A2(N8265), .ZN(N22244));
    NOR2X1 U9373 (.A1(N9149), .A2(N10182), .ZN(n22245));
    INVX1 U9374 (.I(N11019), .ZN(n22246));
    NANDX1 U9375 (.A1(n15056), .A2(n19357), .ZN(n22247));
    NOR2X1 U9376 (.A1(N8075), .A2(n20991), .ZN(N22248));
    INVX1 U9377 (.I(N6835), .ZN(N22249));
    NANDX1 U9378 (.A1(N3374), .A2(N726), .ZN(n22250));
    INVX1 U9379 (.I(N1947), .ZN(N22251));
    NOR2X1 U9380 (.A1(n16604), .A2(N10984), .ZN(n22252));
    NOR2X1 U9381 (.A1(n19814), .A2(n16349), .ZN(n22253));
    NANDX1 U9382 (.A1(n15657), .A2(n16778), .ZN(n22254));
    NANDX1 U9383 (.A1(N6252), .A2(N11944), .ZN(n22255));
    INVX1 U9384 (.I(N4815), .ZN(n22256));
    NOR2X1 U9385 (.A1(n15194), .A2(n13636), .ZN(N22257));
    NANDX1 U9386 (.A1(N6867), .A2(N2004), .ZN(n22258));
    NANDX1 U9387 (.A1(n15326), .A2(N10078), .ZN(n22259));
    INVX1 U9388 (.I(N2542), .ZN(n22260));
    NOR2X1 U9389 (.A1(n20961), .A2(N5915), .ZN(n22261));
    NANDX1 U9390 (.A1(N8992), .A2(N2403), .ZN(N22262));
    NANDX1 U9391 (.A1(N4365), .A2(n13387), .ZN(N22263));
    INVX1 U9392 (.I(n18721), .ZN(n22264));
    NOR2X1 U9393 (.A1(N11462), .A2(n13147), .ZN(n22265));
    INVX1 U9394 (.I(N8210), .ZN(N22266));
    NANDX1 U9395 (.A1(N10537), .A2(n13222), .ZN(n22267));
    NOR2X1 U9396 (.A1(N10399), .A2(N1727), .ZN(n22268));
    NOR2X1 U9397 (.A1(n15820), .A2(N3135), .ZN(n22269));
    NOR2X1 U9398 (.A1(n19368), .A2(n18460), .ZN(n22270));
    NANDX1 U9399 (.A1(n17217), .A2(n15544), .ZN(n22271));
    NANDX1 U9400 (.A1(n16947), .A2(n16000), .ZN(N22272));
    INVX1 U9401 (.I(N4709), .ZN(n22273));
    INVX1 U9402 (.I(N7627), .ZN(n22274));
    INVX1 U9403 (.I(N10559), .ZN(n22275));
    NOR2X1 U9404 (.A1(N1105), .A2(n13605), .ZN(n22276));
    NOR2X1 U9405 (.A1(N8794), .A2(N6741), .ZN(n22277));
    NANDX1 U9406 (.A1(n17276), .A2(n17277), .ZN(n22278));
    NANDX1 U9407 (.A1(N9342), .A2(N987), .ZN(n22279));
    NANDX1 U9408 (.A1(N4128), .A2(n16807), .ZN(n22280));
    NOR2X1 U9409 (.A1(N917), .A2(N9486), .ZN(n22281));
    NANDX1 U9410 (.A1(N7783), .A2(N5472), .ZN(n22282));
    INVX1 U9411 (.I(N10331), .ZN(n22283));
    NOR2X1 U9412 (.A1(N8873), .A2(n14141), .ZN(N22284));
    NANDX1 U9413 (.A1(N6045), .A2(N538), .ZN(n22285));
    NANDX1 U9414 (.A1(N11145), .A2(N12637), .ZN(n22286));
    INVX1 U9415 (.I(n19292), .ZN(N22287));
    NANDX1 U9416 (.A1(n18807), .A2(N4802), .ZN(n22288));
    INVX1 U9417 (.I(n14852), .ZN(n22289));
    NOR2X1 U9418 (.A1(N6204), .A2(n18735), .ZN(n22290));
    NANDX1 U9419 (.A1(n15316), .A2(N1633), .ZN(n22291));
    NOR2X1 U9420 (.A1(N874), .A2(N2549), .ZN(n22292));
    NANDX1 U9421 (.A1(N4892), .A2(N10332), .ZN(n22293));
    INVX1 U9422 (.I(n18995), .ZN(n22294));
    INVX1 U9423 (.I(n12953), .ZN(n22295));
    INVX1 U9424 (.I(N8114), .ZN(n22296));
    INVX1 U9425 (.I(N7224), .ZN(n22297));
    INVX1 U9426 (.I(N6528), .ZN(n22298));
    NOR2X1 U9427 (.A1(n15829), .A2(n16541), .ZN(n22299));
    NANDX1 U9428 (.A1(N9565), .A2(n14117), .ZN(n22300));
    NANDX1 U9429 (.A1(n18696), .A2(N2280), .ZN(n22301));
    INVX1 U9430 (.I(N3669), .ZN(N22302));
    NANDX1 U9431 (.A1(N2080), .A2(n13526), .ZN(N22303));
    INVX1 U9432 (.I(N4346), .ZN(n22304));
    NOR2X1 U9433 (.A1(n19737), .A2(n16097), .ZN(n22305));
    INVX1 U9434 (.I(N3380), .ZN(n22306));
    NOR2X1 U9435 (.A1(N11598), .A2(n13125), .ZN(N22307));
    NANDX1 U9436 (.A1(N12777), .A2(N8), .ZN(n22308));
    INVX1 U9437 (.I(n20000), .ZN(n22309));
    NANDX1 U9438 (.A1(N7356), .A2(n17138), .ZN(n22310));
    INVX1 U9439 (.I(N2666), .ZN(N22311));
    NOR2X1 U9440 (.A1(n17678), .A2(N11324), .ZN(N22312));
    NANDX1 U9441 (.A1(n15143), .A2(n13603), .ZN(n22313));
    INVX1 U9442 (.I(n13354), .ZN(n22314));
    INVX1 U9443 (.I(n19518), .ZN(N22315));
    INVX1 U9444 (.I(N3886), .ZN(n22316));
    INVX1 U9445 (.I(n14590), .ZN(N22317));
    NOR2X1 U9446 (.A1(n13272), .A2(N1735), .ZN(n22318));
    INVX1 U9447 (.I(N4131), .ZN(n22319));
    NANDX1 U9448 (.A1(n13437), .A2(N2485), .ZN(n22320));
    NOR2X1 U9449 (.A1(N7986), .A2(N8771), .ZN(n22321));
    NANDX1 U9450 (.A1(N5728), .A2(n16126), .ZN(n22322));
    NANDX1 U9451 (.A1(n19299), .A2(n13333), .ZN(n22323));
    NANDX1 U9452 (.A1(N10288), .A2(N3426), .ZN(N22324));
    INVX1 U9453 (.I(N4200), .ZN(n22325));
    INVX1 U9454 (.I(N3460), .ZN(n22326));
    INVX1 U9455 (.I(n19497), .ZN(N22327));
    NANDX1 U9456 (.A1(N12286), .A2(N2152), .ZN(n22328));
    NANDX1 U9457 (.A1(N5645), .A2(n20315), .ZN(N22329));
    NANDX1 U9458 (.A1(N7379), .A2(n20627), .ZN(N22330));
    INVX1 U9459 (.I(n15252), .ZN(n22331));
    INVX1 U9460 (.I(n13350), .ZN(N22332));
    NOR2X1 U9461 (.A1(N9903), .A2(N890), .ZN(n22333));
    NOR2X1 U9462 (.A1(N10172), .A2(N11557), .ZN(N22334));
    INVX1 U9463 (.I(N2782), .ZN(n22335));
    NANDX1 U9464 (.A1(N7328), .A2(n13069), .ZN(n22336));
    INVX1 U9465 (.I(N9121), .ZN(n22337));
    NANDX1 U9466 (.A1(n13195), .A2(N12580), .ZN(n22338));
    NANDX1 U9467 (.A1(N11462), .A2(n14327), .ZN(n22339));
    INVX1 U9468 (.I(n13613), .ZN(N22340));
    NANDX1 U9469 (.A1(n20605), .A2(N7240), .ZN(N22341));
    INVX1 U9470 (.I(N1295), .ZN(N22342));
    NOR2X1 U9471 (.A1(n15077), .A2(N11089), .ZN(N22343));
    INVX1 U9472 (.I(N7196), .ZN(N22344));
    NOR2X1 U9473 (.A1(n12997), .A2(N8086), .ZN(n22345));
    NANDX1 U9474 (.A1(N1938), .A2(n14184), .ZN(n22346));
    NOR2X1 U9475 (.A1(N4720), .A2(N12385), .ZN(n22347));
    NANDX1 U9476 (.A1(n17788), .A2(n14010), .ZN(n22348));
    NANDX1 U9477 (.A1(N8368), .A2(N517), .ZN(n22349));
    NOR2X1 U9478 (.A1(N11043), .A2(N11978), .ZN(N22350));
    NANDX1 U9479 (.A1(N10230), .A2(n20132), .ZN(n22351));
    INVX1 U9480 (.I(N4146), .ZN(n22352));
    INVX1 U9481 (.I(N4489), .ZN(n22353));
    NOR2X1 U9482 (.A1(N1861), .A2(n19565), .ZN(N22354));
    NANDX1 U9483 (.A1(N10413), .A2(N5530), .ZN(n22355));
    INVX1 U9484 (.I(n17951), .ZN(n22356));
    NANDX1 U9485 (.A1(N11155), .A2(n19888), .ZN(n22357));
    NOR2X1 U9486 (.A1(N8207), .A2(N3377), .ZN(n22358));
    NANDX1 U9487 (.A1(N7129), .A2(n21165), .ZN(n22359));
    NANDX1 U9488 (.A1(n15172), .A2(N8302), .ZN(n22360));
    NOR2X1 U9489 (.A1(N9106), .A2(n19344), .ZN(n22361));
    NANDX1 U9490 (.A1(n17366), .A2(N2886), .ZN(n22362));
    NOR2X1 U9491 (.A1(n17643), .A2(N1573), .ZN(N22363));
    INVX1 U9492 (.I(n16673), .ZN(n22364));
    NANDX1 U9493 (.A1(N3837), .A2(N9549), .ZN(N22365));
    NOR2X1 U9494 (.A1(N8791), .A2(N9621), .ZN(n22366));
    NANDX1 U9495 (.A1(N5511), .A2(n17777), .ZN(n22367));
    NANDX1 U9496 (.A1(N4169), .A2(N7971), .ZN(N22368));
    NANDX1 U9497 (.A1(N2087), .A2(n16007), .ZN(n22369));
    INVX1 U9498 (.I(N2021), .ZN(n22370));
    INVX1 U9499 (.I(N5592), .ZN(n22371));
    NOR2X1 U9500 (.A1(N7238), .A2(N9239), .ZN(N22372));
    NANDX1 U9501 (.A1(N9631), .A2(N5374), .ZN(n22373));
    INVX1 U9502 (.I(N5467), .ZN(n22374));
    INVX1 U9503 (.I(n17750), .ZN(n22375));
    NOR2X1 U9504 (.A1(n13001), .A2(n19304), .ZN(n22376));
    NOR2X1 U9505 (.A1(N1319), .A2(N5241), .ZN(N22377));
    NOR2X1 U9506 (.A1(N10939), .A2(n17090), .ZN(n22378));
    NOR2X1 U9507 (.A1(N2028), .A2(N3091), .ZN(n22379));
    NANDX1 U9508 (.A1(N9998), .A2(N7612), .ZN(N22380));
    NOR2X1 U9509 (.A1(N4775), .A2(n19262), .ZN(n22381));
    INVX1 U9510 (.I(N10681), .ZN(N22382));
    NANDX1 U9511 (.A1(n16888), .A2(N12460), .ZN(n22383));
    INVX1 U9512 (.I(n14407), .ZN(n22384));
    NOR2X1 U9513 (.A1(N12776), .A2(N3896), .ZN(n22385));
    NANDX1 U9514 (.A1(N9104), .A2(N415), .ZN(n22386));
    NOR2X1 U9515 (.A1(N874), .A2(n14260), .ZN(n22387));
    NANDX1 U9516 (.A1(n17964), .A2(n14042), .ZN(n22388));
    INVX1 U9517 (.I(N7673), .ZN(n22389));
    INVX1 U9518 (.I(n16719), .ZN(n22390));
    INVX1 U9519 (.I(N7533), .ZN(N22391));
    NANDX1 U9520 (.A1(n14239), .A2(N9687), .ZN(n22392));
    NANDX1 U9521 (.A1(n13555), .A2(N7718), .ZN(n22393));
    NOR2X1 U9522 (.A1(n18777), .A2(N5883), .ZN(n22394));
    NOR2X1 U9523 (.A1(N10007), .A2(n13285), .ZN(n22395));
    NANDX1 U9524 (.A1(N10866), .A2(n20603), .ZN(n22396));
    NANDX1 U9525 (.A1(N11734), .A2(N3018), .ZN(N22397));
    NOR2X1 U9526 (.A1(n20044), .A2(N3891), .ZN(N22398));
    INVX1 U9527 (.I(n12945), .ZN(n22399));
    INVX1 U9528 (.I(n14728), .ZN(N22400));
    NOR2X1 U9529 (.A1(n18610), .A2(N3399), .ZN(N22401));
    INVX1 U9530 (.I(N1621), .ZN(n22402));
    NOR2X1 U9531 (.A1(n13892), .A2(n15860), .ZN(n22403));
    NOR2X1 U9532 (.A1(n16985), .A2(N2726), .ZN(n22404));
    INVX1 U9533 (.I(N10871), .ZN(n22405));
    NANDX1 U9534 (.A1(N2071), .A2(n16186), .ZN(n22406));
    INVX1 U9535 (.I(N9897), .ZN(n22407));
    NANDX1 U9536 (.A1(n15686), .A2(N3811), .ZN(n22408));
    INVX1 U9537 (.I(N6189), .ZN(n22409));
    NANDX1 U9538 (.A1(N3491), .A2(n20774), .ZN(n22410));
    NANDX1 U9539 (.A1(N4177), .A2(N12488), .ZN(n22411));
    NOR2X1 U9540 (.A1(n18904), .A2(N799), .ZN(n22412));
    NOR2X1 U9541 (.A1(n16844), .A2(N5828), .ZN(n22413));
    INVX1 U9542 (.I(N1087), .ZN(n22414));
    INVX1 U9543 (.I(N9827), .ZN(n22415));
    NANDX1 U9544 (.A1(n15474), .A2(N7094), .ZN(n22416));
    NANDX1 U9545 (.A1(n20886), .A2(N7366), .ZN(n22417));
    INVX1 U9546 (.I(n15842), .ZN(n22418));
    NANDX1 U9547 (.A1(N8026), .A2(N3831), .ZN(n22419));
    NANDX1 U9548 (.A1(N11836), .A2(N9978), .ZN(N22420));
    NOR2X1 U9549 (.A1(n18664), .A2(n13468), .ZN(n22421));
    NANDX1 U9550 (.A1(n18465), .A2(N12186), .ZN(n22422));
    INVX1 U9551 (.I(n18890), .ZN(n22423));
    NOR2X1 U9552 (.A1(n14743), .A2(N11237), .ZN(N22424));
    INVX1 U9553 (.I(n20570), .ZN(n22425));
    INVX1 U9554 (.I(N1101), .ZN(n22426));
    INVX1 U9555 (.I(n15030), .ZN(n22427));
    NANDX1 U9556 (.A1(N7844), .A2(N893), .ZN(n22428));
    INVX1 U9557 (.I(N7499), .ZN(n22429));
    INVX1 U9558 (.I(n16991), .ZN(N22430));
    NANDX1 U9559 (.A1(n14986), .A2(n19558), .ZN(n22431));
    NANDX1 U9560 (.A1(N397), .A2(N10163), .ZN(N22432));
    INVX1 U9561 (.I(N7769), .ZN(n22433));
    INVX1 U9562 (.I(N2697), .ZN(n22434));
    NANDX1 U9563 (.A1(n15145), .A2(n14883), .ZN(N22435));
    NANDX1 U9564 (.A1(N12804), .A2(n19284), .ZN(n22436));
    NANDX1 U9565 (.A1(n18582), .A2(N3526), .ZN(n22437));
    INVX1 U9566 (.I(N2555), .ZN(n22438));
    NANDX1 U9567 (.A1(N8392), .A2(n17584), .ZN(N22439));
    INVX1 U9568 (.I(n16235), .ZN(N22440));
    NANDX1 U9569 (.A1(n13543), .A2(N2504), .ZN(n22441));
    NOR2X1 U9570 (.A1(N3845), .A2(n20385), .ZN(n22442));
    INVX1 U9571 (.I(N2172), .ZN(n22443));
    INVX1 U9572 (.I(n20285), .ZN(n22444));
    NOR2X1 U9573 (.A1(n15554), .A2(N1365), .ZN(n22445));
    NOR2X1 U9574 (.A1(N12792), .A2(N10590), .ZN(N22446));
    NANDX1 U9575 (.A1(N986), .A2(N12529), .ZN(n22447));
    NANDX1 U9576 (.A1(n20269), .A2(N7981), .ZN(n22448));
    INVX1 U9577 (.I(n18337), .ZN(n22449));
    NANDX1 U9578 (.A1(N4722), .A2(n17505), .ZN(n22450));
    NOR2X1 U9579 (.A1(N1075), .A2(n17644), .ZN(n22451));
    INVX1 U9580 (.I(N8635), .ZN(n22452));
    NANDX1 U9581 (.A1(n18986), .A2(n18995), .ZN(n22453));
    NOR2X1 U9582 (.A1(n18140), .A2(n17653), .ZN(N22454));
    INVX1 U9583 (.I(n17776), .ZN(n22455));
    INVX1 U9584 (.I(N1618), .ZN(n22456));
    INVX1 U9585 (.I(N12613), .ZN(n22457));
    INVX1 U9586 (.I(n13975), .ZN(n22458));
    NANDX1 U9587 (.A1(N2643), .A2(n14960), .ZN(n22459));
    INVX1 U9588 (.I(N7458), .ZN(N22460));
    NOR2X1 U9589 (.A1(n17023), .A2(N9625), .ZN(n22461));
    NANDX1 U9590 (.A1(N8879), .A2(n14346), .ZN(n22462));
    NANDX1 U9591 (.A1(n14584), .A2(N9962), .ZN(n22463));
    NANDX1 U9592 (.A1(N9836), .A2(n13139), .ZN(n22464));
    INVX1 U9593 (.I(N7591), .ZN(n22465));
    NANDX1 U9594 (.A1(N11173), .A2(N4501), .ZN(n22466));
    INVX1 U9595 (.I(N457), .ZN(N22467));
    NANDX1 U9596 (.A1(n13115), .A2(n17846), .ZN(n22468));
    NOR2X1 U9597 (.A1(N4497), .A2(n17561), .ZN(n22469));
    NOR2X1 U9598 (.A1(N1010), .A2(n14746), .ZN(N22470));
    NOR2X1 U9599 (.A1(N10052), .A2(n16745), .ZN(n22471));
    NOR2X1 U9600 (.A1(N386), .A2(N5139), .ZN(N22472));
    INVX1 U9601 (.I(N9264), .ZN(N22473));
    INVX1 U9602 (.I(n15122), .ZN(n22474));
    NOR2X1 U9603 (.A1(n18530), .A2(N2539), .ZN(n22475));
    NOR2X1 U9604 (.A1(N4980), .A2(n15684), .ZN(n22476));
    INVX1 U9605 (.I(N10424), .ZN(n22477));
    NANDX1 U9606 (.A1(n13627), .A2(N12291), .ZN(n22478));
    INVX1 U9607 (.I(N9215), .ZN(n22479));
    NANDX1 U9608 (.A1(n13012), .A2(N5985), .ZN(n22480));
    NOR2X1 U9609 (.A1(N9342), .A2(n16729), .ZN(n22481));
    NOR2X1 U9610 (.A1(n18629), .A2(n15744), .ZN(n22482));
    NOR2X1 U9611 (.A1(n14144), .A2(N7528), .ZN(n22483));
    NANDX1 U9612 (.A1(n13824), .A2(n20729), .ZN(n22484));
    NOR2X1 U9613 (.A1(N1162), .A2(N9163), .ZN(n22485));
    NOR2X1 U9614 (.A1(n19691), .A2(N11701), .ZN(n22486));
    NANDX1 U9615 (.A1(N3440), .A2(N6154), .ZN(n22487));
    NOR2X1 U9616 (.A1(N8405), .A2(N6322), .ZN(N22488));
    INVX1 U9617 (.I(n20695), .ZN(N22489));
    NOR2X1 U9618 (.A1(n16980), .A2(n19412), .ZN(N22490));
    NOR2X1 U9619 (.A1(n17506), .A2(n17167), .ZN(n22491));
    INVX1 U9620 (.I(N7546), .ZN(n22492));
    INVX1 U9621 (.I(n15780), .ZN(n22493));
    INVX1 U9622 (.I(n19289), .ZN(n22494));
    NOR2X1 U9623 (.A1(N9586), .A2(n17573), .ZN(N22495));
    INVX1 U9624 (.I(N9085), .ZN(n22496));
    INVX1 U9625 (.I(N2448), .ZN(n22497));
    INVX1 U9626 (.I(N3139), .ZN(N22498));
    NANDX1 U9627 (.A1(N3259), .A2(N9381), .ZN(n22499));
    INVX1 U9628 (.I(N3955), .ZN(n22500));
    NANDX1 U9629 (.A1(N1835), .A2(N4818), .ZN(n22501));
    NOR2X1 U9630 (.A1(n17072), .A2(N6304), .ZN(n22502));
    INVX1 U9631 (.I(N9795), .ZN(N22503));
    NANDX1 U9632 (.A1(n19080), .A2(N273), .ZN(n22504));
    NANDX1 U9633 (.A1(N5395), .A2(n16203), .ZN(n22505));
    INVX1 U9634 (.I(N7454), .ZN(n22506));
    NANDX1 U9635 (.A1(n15737), .A2(n17039), .ZN(n22507));
    NOR2X1 U9636 (.A1(N11565), .A2(n20665), .ZN(n22508));
    INVX1 U9637 (.I(N8554), .ZN(n22509));
    NOR2X1 U9638 (.A1(N6716), .A2(N4003), .ZN(N22510));
    INVX1 U9639 (.I(n16096), .ZN(N22511));
    NANDX1 U9640 (.A1(n13978), .A2(n19614), .ZN(N22512));
    NANDX1 U9641 (.A1(n18795), .A2(N9668), .ZN(n22513));
    INVX1 U9642 (.I(N3868), .ZN(n22514));
    NOR2X1 U9643 (.A1(n15216), .A2(n19211), .ZN(n22515));
    NANDX1 U9644 (.A1(N10030), .A2(N10475), .ZN(N22516));
    NOR2X1 U9645 (.A1(N5003), .A2(n17519), .ZN(N22517));
    INVX1 U9646 (.I(N8347), .ZN(n22518));
    NOR2X1 U9647 (.A1(N6832), .A2(N8034), .ZN(n22519));
    NOR2X1 U9648 (.A1(N808), .A2(N11611), .ZN(N22520));
    NANDX1 U9649 (.A1(n13031), .A2(n18326), .ZN(N22521));
    NOR2X1 U9650 (.A1(N1824), .A2(N7733), .ZN(n22522));
    INVX1 U9651 (.I(n15801), .ZN(N22523));
    NOR2X1 U9652 (.A1(N5552), .A2(N7907), .ZN(n22524));
    NANDX1 U9653 (.A1(N5516), .A2(N6316), .ZN(n22525));
    NANDX1 U9654 (.A1(n15273), .A2(N4297), .ZN(n22526));
    INVX1 U9655 (.I(N4073), .ZN(n22527));
    NOR2X1 U9656 (.A1(N2082), .A2(N3617), .ZN(N22528));
    NANDX1 U9657 (.A1(n13104), .A2(N11963), .ZN(n22529));
    NANDX1 U9658 (.A1(n19935), .A2(n19997), .ZN(n22530));
    INVX1 U9659 (.I(n15285), .ZN(n22531));
    NOR2X1 U9660 (.A1(n14520), .A2(N7085), .ZN(n22532));
    INVX1 U9661 (.I(n18517), .ZN(n22533));
    INVX1 U9662 (.I(N4289), .ZN(n22534));
    NANDX1 U9663 (.A1(n19250), .A2(n20719), .ZN(n22535));
    NOR2X1 U9664 (.A1(N5926), .A2(N4356), .ZN(n22536));
    INVX1 U9665 (.I(N12241), .ZN(N22537));
    NANDX1 U9666 (.A1(N3223), .A2(N11079), .ZN(n22538));
    NANDX1 U9667 (.A1(N7295), .A2(n20392), .ZN(n22539));
    NANDX1 U9668 (.A1(N10911), .A2(N4762), .ZN(n22540));
    NANDX1 U9669 (.A1(N1644), .A2(n16929), .ZN(N22541));
    NANDX1 U9670 (.A1(n16182), .A2(N4765), .ZN(n22542));
    NOR2X1 U9671 (.A1(N5328), .A2(n13827), .ZN(n22543));
    INVX1 U9672 (.I(N1884), .ZN(n22544));
    NANDX1 U9673 (.A1(N4704), .A2(N715), .ZN(n22545));
    NANDX1 U9674 (.A1(N2723), .A2(N203), .ZN(n22546));
    NANDX1 U9675 (.A1(N3190), .A2(n20331), .ZN(N22547));
    NOR2X1 U9676 (.A1(N9973), .A2(N8649), .ZN(n22548));
    NOR2X1 U9677 (.A1(n15593), .A2(N11250), .ZN(N22549));
    INVX1 U9678 (.I(n14754), .ZN(n22550));
    NANDX1 U9679 (.A1(N1039), .A2(n14058), .ZN(N22551));
    INVX1 U9680 (.I(n18454), .ZN(N22552));
    NANDX1 U9681 (.A1(N1689), .A2(n13405), .ZN(n22553));
    NOR2X1 U9682 (.A1(N1318), .A2(n13275), .ZN(n22554));
    INVX1 U9683 (.I(N2572), .ZN(n22555));
    INVX1 U9684 (.I(n17627), .ZN(n22556));
    NANDX1 U9685 (.A1(N10414), .A2(N165), .ZN(n22557));
    NOR2X1 U9686 (.A1(N10617), .A2(n13056), .ZN(n22558));
    NANDX1 U9687 (.A1(N9717), .A2(n13897), .ZN(n22559));
    NANDX1 U9688 (.A1(n12907), .A2(n17960), .ZN(N22560));
    NOR2X1 U9689 (.A1(n18698), .A2(N8088), .ZN(N22561));
    NANDX1 U9690 (.A1(N7942), .A2(N3669), .ZN(n22562));
    NANDX1 U9691 (.A1(N4056), .A2(N892), .ZN(N22563));
    INVX1 U9692 (.I(N287), .ZN(n22564));
    NANDX1 U9693 (.A1(N5713), .A2(N1604), .ZN(n22565));
    NANDX1 U9694 (.A1(N12227), .A2(n19947), .ZN(n22566));
    NANDX1 U9695 (.A1(N8623), .A2(N5992), .ZN(n22567));
    NANDX1 U9696 (.A1(N8787), .A2(N5074), .ZN(N22568));
    INVX1 U9697 (.I(N612), .ZN(n22569));
    INVX1 U9698 (.I(N9182), .ZN(n22570));
    NANDX1 U9699 (.A1(n14130), .A2(n16630), .ZN(n22571));
    NOR2X1 U9700 (.A1(n15277), .A2(n14097), .ZN(n22572));
    INVX1 U9701 (.I(N4490), .ZN(n22573));
    NANDX1 U9702 (.A1(N12077), .A2(N2302), .ZN(n22574));
    NANDX1 U9703 (.A1(N7510), .A2(n20183), .ZN(n22575));
    INVX1 U9704 (.I(n16348), .ZN(n22576));
    INVX1 U9705 (.I(N11609), .ZN(n22577));
    NOR2X1 U9706 (.A1(N11434), .A2(N10326), .ZN(N22578));
    NANDX1 U9707 (.A1(n14598), .A2(N10859), .ZN(n22579));
    INVX1 U9708 (.I(N2154), .ZN(n22580));
    INVX1 U9709 (.I(N5210), .ZN(n22581));
    NANDX1 U9710 (.A1(N2046), .A2(n14391), .ZN(n22582));
    INVX1 U9711 (.I(N10717), .ZN(n22583));
    INVX1 U9712 (.I(N12134), .ZN(n22584));
    NOR2X1 U9713 (.A1(n18428), .A2(n20542), .ZN(n22585));
    NOR2X1 U9714 (.A1(N8320), .A2(N11388), .ZN(n22586));
    NOR2X1 U9715 (.A1(N2268), .A2(n18898), .ZN(n22587));
    NOR2X1 U9716 (.A1(N12273), .A2(n14015), .ZN(n22588));
    NOR2X1 U9717 (.A1(N2652), .A2(n20329), .ZN(N22589));
    INVX1 U9718 (.I(N7519), .ZN(n22590));
    INVX1 U9719 (.I(n19370), .ZN(n22591));
    NOR2X1 U9720 (.A1(n16280), .A2(n16065), .ZN(n22592));
    INVX1 U9721 (.I(N259), .ZN(n22593));
    NOR2X1 U9722 (.A1(N9666), .A2(N9191), .ZN(n22594));
    NOR2X1 U9723 (.A1(n20383), .A2(n13522), .ZN(N22595));
    NOR2X1 U9724 (.A1(n19688), .A2(N5261), .ZN(n22596));
    INVX1 U9725 (.I(n18024), .ZN(N22597));
    INVX1 U9726 (.I(N10413), .ZN(n22598));
    NOR2X1 U9727 (.A1(N10390), .A2(N8080), .ZN(n22599));
    NOR2X1 U9728 (.A1(N1432), .A2(n16636), .ZN(n22600));
    NANDX1 U9729 (.A1(n19855), .A2(N10276), .ZN(n22601));
    INVX1 U9730 (.I(N6143), .ZN(n22602));
    NANDX1 U9731 (.A1(n13902), .A2(N3290), .ZN(n22603));
    NANDX1 U9732 (.A1(N3279), .A2(N10910), .ZN(n22604));
    NOR2X1 U9733 (.A1(N11191), .A2(n15117), .ZN(n22605));
    NOR2X1 U9734 (.A1(N4229), .A2(N8811), .ZN(N22606));
    NANDX1 U9735 (.A1(N3942), .A2(N7268), .ZN(n22607));
    NOR2X1 U9736 (.A1(N2966), .A2(n19834), .ZN(n22608));
    INVX1 U9737 (.I(N7920), .ZN(n22609));
    INVX1 U9738 (.I(n14683), .ZN(n22610));
    INVX1 U9739 (.I(n19143), .ZN(n22611));
    INVX1 U9740 (.I(N489), .ZN(n22612));
    NOR2X1 U9741 (.A1(n14739), .A2(N10764), .ZN(n22613));
    INVX1 U9742 (.I(n15423), .ZN(n22614));
    NOR2X1 U9743 (.A1(N1564), .A2(n18712), .ZN(n22615));
    NANDX1 U9744 (.A1(N4842), .A2(N2933), .ZN(n22616));
    NANDX1 U9745 (.A1(N10575), .A2(n18050), .ZN(n22617));
    NANDX1 U9746 (.A1(n14803), .A2(N5630), .ZN(N22618));
    INVX1 U9747 (.I(n13286), .ZN(n22619));
    INVX1 U9748 (.I(N6191), .ZN(n22620));
    NANDX1 U9749 (.A1(N6043), .A2(N10484), .ZN(N22621));
    INVX1 U9750 (.I(N12391), .ZN(N22622));
    NOR2X1 U9751 (.A1(N2565), .A2(N4846), .ZN(n22623));
    INVX1 U9752 (.I(N3053), .ZN(n22624));
    INVX1 U9753 (.I(N2641), .ZN(n22625));
    INVX1 U9754 (.I(N1410), .ZN(n22626));
    INVX1 U9755 (.I(n13245), .ZN(n22627));
    NANDX1 U9756 (.A1(N10087), .A2(N7302), .ZN(n22628));
    NOR2X1 U9757 (.A1(n13020), .A2(N12019), .ZN(N22629));
    NANDX1 U9758 (.A1(N4381), .A2(n15356), .ZN(n22630));
    NOR2X1 U9759 (.A1(N4552), .A2(N4145), .ZN(N22631));
    NANDX1 U9760 (.A1(N11991), .A2(N10335), .ZN(n22632));
    INVX1 U9761 (.I(N12575), .ZN(n22633));
    INVX1 U9762 (.I(N11688), .ZN(N22634));
    INVX1 U9763 (.I(n19295), .ZN(n22635));
    INVX1 U9764 (.I(N3123), .ZN(n22636));
    INVX1 U9765 (.I(N11847), .ZN(n22637));
    NANDX1 U9766 (.A1(N9838), .A2(n20205), .ZN(N22638));
    NANDX1 U9767 (.A1(N1213), .A2(N6761), .ZN(n22639));
    INVX1 U9768 (.I(N5841), .ZN(n22640));
    INVX1 U9769 (.I(N7233), .ZN(n22641));
    NOR2X1 U9770 (.A1(n20623), .A2(N9247), .ZN(n22642));
    NOR2X1 U9771 (.A1(n14748), .A2(N4833), .ZN(n22643));
    NANDX1 U9772 (.A1(n18892), .A2(N8246), .ZN(n22644));
    INVX1 U9773 (.I(N2538), .ZN(n22645));
    INVX1 U9774 (.I(n20211), .ZN(n22646));
    INVX1 U9775 (.I(N7451), .ZN(n22647));
    NOR2X1 U9776 (.A1(N10503), .A2(n16245), .ZN(N22648));
    INVX1 U9777 (.I(n17700), .ZN(n22649));
    NANDX1 U9778 (.A1(N11791), .A2(N849), .ZN(N22650));
    NANDX1 U9779 (.A1(N8839), .A2(n17833), .ZN(n22651));
    NANDX1 U9780 (.A1(n13715), .A2(N2443), .ZN(n22652));
    NOR2X1 U9781 (.A1(n20948), .A2(n15845), .ZN(n22653));
    NOR2X1 U9782 (.A1(N8964), .A2(N12396), .ZN(n22654));
    NOR2X1 U9783 (.A1(n13797), .A2(N8041), .ZN(n22655));
    INVX1 U9784 (.I(n16584), .ZN(N22656));
    NOR2X1 U9785 (.A1(n19166), .A2(n17805), .ZN(n22657));
    NANDX1 U9786 (.A1(N10374), .A2(N4026), .ZN(n22658));
    INVX1 U9787 (.I(n20877), .ZN(N22659));
    NANDX1 U9788 (.A1(N1377), .A2(N11888), .ZN(n22660));
    INVX1 U9789 (.I(n13167), .ZN(n22661));
    NOR2X1 U9790 (.A1(n16593), .A2(n16547), .ZN(n22662));
    INVX1 U9791 (.I(n18273), .ZN(n22663));
    NOR2X1 U9792 (.A1(N6322), .A2(N12785), .ZN(N22664));
    NANDX1 U9793 (.A1(n16708), .A2(N1231), .ZN(n22665));
    NANDX1 U9794 (.A1(N2416), .A2(N4425), .ZN(n22666));
    NOR2X1 U9795 (.A1(N10456), .A2(n21053), .ZN(n22667));
    INVX1 U9796 (.I(n20674), .ZN(n22668));
    NOR2X1 U9797 (.A1(N7062), .A2(N8642), .ZN(n22669));
    NANDX1 U9798 (.A1(N5629), .A2(N9639), .ZN(n22670));
    NANDX1 U9799 (.A1(n20440), .A2(N5557), .ZN(n22671));
    NANDX1 U9800 (.A1(n15425), .A2(n13265), .ZN(n22672));
    INVX1 U9801 (.I(N5329), .ZN(n22673));
    INVX1 U9802 (.I(n19904), .ZN(n22674));
    NANDX1 U9803 (.A1(N12154), .A2(n20768), .ZN(n22675));
    NOR2X1 U9804 (.A1(N9985), .A2(N10787), .ZN(N22676));
    NOR2X1 U9805 (.A1(N1008), .A2(n13202), .ZN(N22677));
    NOR2X1 U9806 (.A1(n16141), .A2(n18200), .ZN(n22678));
    INVX1 U9807 (.I(N5398), .ZN(n22679));
    INVX1 U9808 (.I(N2015), .ZN(n22680));
    INVX1 U9809 (.I(n20827), .ZN(n22681));
    INVX1 U9810 (.I(N7171), .ZN(N22682));
    NANDX1 U9811 (.A1(N1548), .A2(N6380), .ZN(N22683));
    INVX1 U9812 (.I(N4837), .ZN(N22684));
    NOR2X1 U9813 (.A1(n17140), .A2(n20862), .ZN(n22685));
    INVX1 U9814 (.I(n20263), .ZN(n22686));
    NANDX1 U9815 (.A1(n18586), .A2(N5728), .ZN(n22687));
    INVX1 U9816 (.I(N1594), .ZN(n22688));
    NOR2X1 U9817 (.A1(n18943), .A2(N12521), .ZN(n22689));
    NANDX1 U9818 (.A1(N10914), .A2(N1184), .ZN(n22690));
    NOR2X1 U9819 (.A1(N2425), .A2(N10899), .ZN(n22691));
    NANDX1 U9820 (.A1(n14610), .A2(n12913), .ZN(n22692));
    NOR2X1 U9821 (.A1(n14206), .A2(N12141), .ZN(N22693));
    NANDX1 U9822 (.A1(N12524), .A2(N8230), .ZN(N22694));
    NANDX1 U9823 (.A1(n16399), .A2(n13067), .ZN(n22695));
    INVX1 U9824 (.I(N6851), .ZN(n22696));
    NOR2X1 U9825 (.A1(N388), .A2(N425), .ZN(n22697));
    NANDX1 U9826 (.A1(n13515), .A2(N6152), .ZN(n22698));
    NOR2X1 U9827 (.A1(n15109), .A2(n16405), .ZN(N22699));
    NOR2X1 U9828 (.A1(N6399), .A2(N6436), .ZN(n22700));
    INVX1 U9829 (.I(N2124), .ZN(n22701));
    NANDX1 U9830 (.A1(n13834), .A2(n13022), .ZN(n22702));
    NOR2X1 U9831 (.A1(N1755), .A2(n20476), .ZN(n22703));
    NOR2X1 U9832 (.A1(n15960), .A2(N5928), .ZN(N22704));
    INVX1 U9833 (.I(N1795), .ZN(N22705));
    INVX1 U9834 (.I(n18731), .ZN(N22706));
    INVX1 U9835 (.I(N536), .ZN(n22707));
    INVX1 U9836 (.I(n14128), .ZN(n22708));
    INVX1 U9837 (.I(n19062), .ZN(N22709));
    NOR2X1 U9838 (.A1(N7860), .A2(N11346), .ZN(n22710));
    NOR2X1 U9839 (.A1(N10643), .A2(n20996), .ZN(n22711));
    NANDX1 U9840 (.A1(n16596), .A2(N706), .ZN(n22712));
    INVX1 U9841 (.I(N1317), .ZN(n22713));
    NOR2X1 U9842 (.A1(n13088), .A2(N9692), .ZN(N22714));
    NOR2X1 U9843 (.A1(N9973), .A2(N11446), .ZN(N22715));
    NANDX1 U9844 (.A1(N9053), .A2(N717), .ZN(n22716));
    NOR2X1 U9845 (.A1(n17498), .A2(n18283), .ZN(n22717));
    INVX1 U9846 (.I(n14998), .ZN(n22718));
    NOR2X1 U9847 (.A1(N3569), .A2(n17900), .ZN(n22719));
    NOR2X1 U9848 (.A1(N11343), .A2(N10273), .ZN(n22720));
    NANDX1 U9849 (.A1(n13744), .A2(N389), .ZN(n22721));
    NANDX1 U9850 (.A1(N3157), .A2(n15926), .ZN(n22722));
    INVX1 U9851 (.I(n14294), .ZN(n22723));
    INVX1 U9852 (.I(N6377), .ZN(N22724));
    NANDX1 U9853 (.A1(n19460), .A2(n14006), .ZN(n22725));
    NOR2X1 U9854 (.A1(N8622), .A2(n18520), .ZN(n22726));
    NANDX1 U9855 (.A1(n18258), .A2(N6343), .ZN(N22727));
    NANDX1 U9856 (.A1(N7134), .A2(N2610), .ZN(n22728));
    NANDX1 U9857 (.A1(N10167), .A2(n17607), .ZN(n22729));
    INVX1 U9858 (.I(n13735), .ZN(N22730));
    INVX1 U9859 (.I(N9383), .ZN(n22731));
    NOR2X1 U9860 (.A1(n19091), .A2(n21160), .ZN(n22732));
    INVX1 U9861 (.I(n14021), .ZN(n22733));
    NOR2X1 U9862 (.A1(N9831), .A2(N8717), .ZN(n22734));
    NOR2X1 U9863 (.A1(N2894), .A2(N4118), .ZN(n22735));
    INVX1 U9864 (.I(n13046), .ZN(n22736));
    NOR2X1 U9865 (.A1(N10167), .A2(N11658), .ZN(N22737));
    NOR2X1 U9866 (.A1(N7456), .A2(n16258), .ZN(n22738));
    NANDX1 U9867 (.A1(n13798), .A2(N343), .ZN(n22739));
    NOR2X1 U9868 (.A1(N10949), .A2(N2711), .ZN(n22740));
    NANDX1 U9869 (.A1(N1868), .A2(N9409), .ZN(n22741));
    INVX1 U9870 (.I(N10686), .ZN(n22742));
    NANDX1 U9871 (.A1(n21045), .A2(N3088), .ZN(n22743));
    NANDX1 U9872 (.A1(N6489), .A2(N11651), .ZN(n22744));
    NANDX1 U9873 (.A1(N10861), .A2(n14909), .ZN(n22745));
    NANDX1 U9874 (.A1(N8296), .A2(n19026), .ZN(n22746));
    NOR2X1 U9875 (.A1(N111), .A2(N10456), .ZN(n22747));
    NOR2X1 U9876 (.A1(N6311), .A2(n15966), .ZN(n22748));
    NOR2X1 U9877 (.A1(N1338), .A2(n18503), .ZN(N22749));
    INVX1 U9878 (.I(n17452), .ZN(n22750));
    NANDX1 U9879 (.A1(n20609), .A2(n14705), .ZN(n22751));
    INVX1 U9880 (.I(N1246), .ZN(n22752));
    NOR2X1 U9881 (.A1(n17290), .A2(N11931), .ZN(n22753));
    NANDX1 U9882 (.A1(n17104), .A2(N9560), .ZN(n22754));
    INVX1 U9883 (.I(n18134), .ZN(n22755));
    INVX1 U9884 (.I(N5999), .ZN(n22756));
    NOR2X1 U9885 (.A1(n14888), .A2(n20224), .ZN(n22757));
    INVX1 U9886 (.I(N7225), .ZN(n22758));
    INVX1 U9887 (.I(N10712), .ZN(n22759));
    INVX1 U9888 (.I(N8703), .ZN(n22760));
    NOR2X1 U9889 (.A1(N12416), .A2(N4565), .ZN(N22761));
    NANDX1 U9890 (.A1(N4230), .A2(n14225), .ZN(n22762));
    NANDX1 U9891 (.A1(N5714), .A2(n13603), .ZN(n22763));
    INVX1 U9892 (.I(n16120), .ZN(N22764));
    INVX1 U9893 (.I(n15792), .ZN(n22765));
    NANDX1 U9894 (.A1(N90), .A2(N10776), .ZN(n22766));
    NANDX1 U9895 (.A1(N4191), .A2(n19022), .ZN(n22767));
    NANDX1 U9896 (.A1(N4171), .A2(N3790), .ZN(n22768));
    INVX1 U9897 (.I(n13600), .ZN(N22769));
    NOR2X1 U9898 (.A1(n17860), .A2(n20825), .ZN(n22770));
    NOR2X1 U9899 (.A1(N7341), .A2(N11817), .ZN(n22771));
    INVX1 U9900 (.I(n18904), .ZN(n22772));
    NANDX1 U9901 (.A1(n14514), .A2(N5116), .ZN(n22773));
    INVX1 U9902 (.I(N7508), .ZN(n22774));
    NOR2X1 U9903 (.A1(N2028), .A2(n15652), .ZN(n22775));
    INVX1 U9904 (.I(n18147), .ZN(n22776));
    INVX1 U9905 (.I(n16251), .ZN(n22777));
    NANDX1 U9906 (.A1(N3900), .A2(N5796), .ZN(n22778));
    INVX1 U9907 (.I(N8091), .ZN(N22779));
    NOR2X1 U9908 (.A1(N11184), .A2(N12261), .ZN(N22780));
    INVX1 U9909 (.I(n18443), .ZN(n22781));
    INVX1 U9910 (.I(n20473), .ZN(N22782));
    NANDX1 U9911 (.A1(n19996), .A2(N489), .ZN(N22783));
    NOR2X1 U9912 (.A1(N5124), .A2(N10438), .ZN(n22784));
    NOR2X1 U9913 (.A1(N2667), .A2(n19494), .ZN(n22785));
    NOR2X1 U9914 (.A1(n20211), .A2(N313), .ZN(n22786));
    NOR2X1 U9915 (.A1(N1009), .A2(n15965), .ZN(n22787));
    INVX1 U9916 (.I(n13697), .ZN(n22788));
    NANDX1 U9917 (.A1(n13086), .A2(N1562), .ZN(n22789));
    NOR2X1 U9918 (.A1(n13423), .A2(N7791), .ZN(N22790));
    NOR2X1 U9919 (.A1(N11552), .A2(n18975), .ZN(n22791));
    INVX1 U9920 (.I(N8011), .ZN(N22792));
    INVX1 U9921 (.I(n16508), .ZN(n22793));
    INVX1 U9922 (.I(n20343), .ZN(N22794));
    NANDX1 U9923 (.A1(N2284), .A2(N10610), .ZN(n22795));
    NANDX1 U9924 (.A1(N7263), .A2(n14322), .ZN(n22796));
    NANDX1 U9925 (.A1(N68), .A2(N1919), .ZN(N22797));
    INVX1 U9926 (.I(N381), .ZN(n22798));
    NOR2X1 U9927 (.A1(N6678), .A2(n16345), .ZN(n22799));
    NOR2X1 U9928 (.A1(n20375), .A2(n14889), .ZN(n22800));
    NANDX1 U9929 (.A1(n16478), .A2(N11875), .ZN(n22801));
    NOR2X1 U9930 (.A1(N3038), .A2(N1179), .ZN(n22802));
    NANDX1 U9931 (.A1(n16554), .A2(n13057), .ZN(n22803));
    NANDX1 U9932 (.A1(N6053), .A2(N2877), .ZN(N22804));
    NANDX1 U9933 (.A1(n20937), .A2(N12692), .ZN(n22805));
    NOR2X1 U9934 (.A1(N4858), .A2(N942), .ZN(N22806));
    INVX1 U9935 (.I(n13721), .ZN(n22807));
    NOR2X1 U9936 (.A1(n15003), .A2(n15640), .ZN(n22808));
    NANDX1 U9937 (.A1(n15383), .A2(n13935), .ZN(N22809));
    INVX1 U9938 (.I(N5039), .ZN(N22810));
    NANDX1 U9939 (.A1(N3350), .A2(n19928), .ZN(n22811));
    NOR2X1 U9940 (.A1(n19827), .A2(N10572), .ZN(n22812));
    NOR2X1 U9941 (.A1(n17407), .A2(N6293), .ZN(n22813));
    NANDX1 U9942 (.A1(N12730), .A2(n19349), .ZN(n22814));
    NOR2X1 U9943 (.A1(n13324), .A2(n16767), .ZN(n22815));
    INVX1 U9944 (.I(N7573), .ZN(n22816));
    INVX1 U9945 (.I(N3241), .ZN(n22817));
    INVX1 U9946 (.I(N3712), .ZN(N22818));
    NANDX1 U9947 (.A1(n20693), .A2(N11342), .ZN(N22819));
    NOR2X1 U9948 (.A1(n15102), .A2(N8870), .ZN(n22820));
    NOR2X1 U9949 (.A1(N2348), .A2(n13076), .ZN(N22821));
    NANDX1 U9950 (.A1(N5954), .A2(N10967), .ZN(N22822));
    NOR2X1 U9951 (.A1(N12317), .A2(N4106), .ZN(N22823));
    NANDX1 U9952 (.A1(N8171), .A2(N282), .ZN(N22824));
    NOR2X1 U9953 (.A1(n20840), .A2(n13011), .ZN(n22825));
    NOR2X1 U9954 (.A1(N5560), .A2(n20877), .ZN(n22826));
    NANDX1 U9955 (.A1(n16900), .A2(N7219), .ZN(N22827));
    NOR2X1 U9956 (.A1(n20140), .A2(n14190), .ZN(n22828));
    NOR2X1 U9957 (.A1(n17085), .A2(n13652), .ZN(N22829));
    NANDX1 U9958 (.A1(N2344), .A2(N2065), .ZN(n22830));
    NOR2X1 U9959 (.A1(N2986), .A2(N4412), .ZN(N22831));
    NOR2X1 U9960 (.A1(N8667), .A2(N10365), .ZN(n22832));
    INVX1 U9961 (.I(N7586), .ZN(n22833));
    NANDX1 U9962 (.A1(n15757), .A2(n17077), .ZN(N22834));
    INVX1 U9963 (.I(n16038), .ZN(n22835));
    NOR2X1 U9964 (.A1(n19545), .A2(N2360), .ZN(n22836));
    NOR2X1 U9965 (.A1(n19647), .A2(n17778), .ZN(n22837));
    INVX1 U9966 (.I(n15316), .ZN(n22838));
    NOR2X1 U9967 (.A1(N3513), .A2(n14225), .ZN(n22839));
    INVX1 U9968 (.I(N3058), .ZN(N22840));
    INVX1 U9969 (.I(N4919), .ZN(n22841));
    NANDX1 U9970 (.A1(N1506), .A2(N1526), .ZN(N22842));
    NANDX1 U9971 (.A1(N4492), .A2(N5937), .ZN(n22843));
    NOR2X1 U9972 (.A1(N7700), .A2(N10844), .ZN(n22844));
    NOR2X1 U9973 (.A1(n15285), .A2(N6836), .ZN(n22845));
    INVX1 U9974 (.I(N5674), .ZN(N22846));
    INVX1 U9975 (.I(N3222), .ZN(n22847));
    INVX1 U9976 (.I(n14170), .ZN(n22848));
    INVX1 U9977 (.I(N4628), .ZN(n22849));
    INVX1 U9978 (.I(n17901), .ZN(N22850));
    INVX1 U9979 (.I(N6671), .ZN(n22851));
    NANDX1 U9980 (.A1(N4904), .A2(n15437), .ZN(n22852));
    NANDX1 U9981 (.A1(N7961), .A2(n14599), .ZN(n22853));
    NOR2X1 U9982 (.A1(n16446), .A2(n16104), .ZN(n22854));
    NOR2X1 U9983 (.A1(N2226), .A2(n15137), .ZN(n22855));
    INVX1 U9984 (.I(N4463), .ZN(n22856));
    NOR2X1 U9985 (.A1(n19782), .A2(N2579), .ZN(n22857));
    NANDX1 U9986 (.A1(n21160), .A2(N10993), .ZN(n22858));
    NOR2X1 U9987 (.A1(N12), .A2(N8756), .ZN(n22859));
    INVX1 U9988 (.I(n14181), .ZN(N22860));
    NOR2X1 U9989 (.A1(n17204), .A2(N5536), .ZN(N22861));
    NANDX1 U9990 (.A1(N2822), .A2(N6748), .ZN(n22862));
    INVX1 U9991 (.I(N2267), .ZN(n22863));
    INVX1 U9992 (.I(n18315), .ZN(n22864));
    NOR2X1 U9993 (.A1(N10094), .A2(n19792), .ZN(n22865));
    NOR2X1 U9994 (.A1(n20740), .A2(N1564), .ZN(n22866));
    NOR2X1 U9995 (.A1(N9188), .A2(N10502), .ZN(n22867));
    INVX1 U9996 (.I(N5336), .ZN(n22868));
    NANDX1 U9997 (.A1(N3793), .A2(N11310), .ZN(n22869));
    INVX1 U9998 (.I(N9327), .ZN(n22870));
    INVX1 U9999 (.I(N8994), .ZN(n22871));
    NOR2X1 U10000 (.A1(N8844), .A2(n17717), .ZN(n22872));
    NOR2X1 U10001 (.A1(n20589), .A2(N2022), .ZN(N22873));
    NANDX1 U10002 (.A1(n17953), .A2(N3312), .ZN(n22874));
    NANDX1 U10003 (.A1(n20219), .A2(N4265), .ZN(n22875));
    NANDX1 U10004 (.A1(N3758), .A2(N8901), .ZN(N22876));
    NANDX1 U10005 (.A1(N3741), .A2(N8410), .ZN(n22877));
    INVX1 U10006 (.I(n16264), .ZN(n22878));
    INVX1 U10007 (.I(N2538), .ZN(n22879));
    NOR2X1 U10008 (.A1(N12016), .A2(N11591), .ZN(N22880));
    NANDX1 U10009 (.A1(N2095), .A2(n15115), .ZN(n22881));
    NANDX1 U10010 (.A1(n14135), .A2(N2878), .ZN(n22882));
    NANDX1 U10011 (.A1(N1749), .A2(n15136), .ZN(n22883));
    NANDX1 U10012 (.A1(N1107), .A2(n17158), .ZN(N22884));
    NOR2X1 U10013 (.A1(n13601), .A2(n20469), .ZN(n22885));
    NOR2X1 U10014 (.A1(N12590), .A2(n19275), .ZN(n22886));
    INVX1 U10015 (.I(n16347), .ZN(n22887));
    NOR2X1 U10016 (.A1(N10150), .A2(n14629), .ZN(N22888));
    INVX1 U10017 (.I(N2185), .ZN(n22889));
    NOR2X1 U10018 (.A1(n16577), .A2(N4722), .ZN(n22890));
    NANDX1 U10019 (.A1(N7362), .A2(N10854), .ZN(n22891));
    INVX1 U10020 (.I(N3999), .ZN(n22892));
    NANDX1 U10021 (.A1(N9254), .A2(n18133), .ZN(N22893));
    NANDX1 U10022 (.A1(N4556), .A2(n14423), .ZN(n22894));
    NANDX1 U10023 (.A1(n15901), .A2(N10072), .ZN(N22895));
    INVX1 U10024 (.I(n16693), .ZN(n22896));
    NOR2X1 U10025 (.A1(N7000), .A2(N1998), .ZN(n22897));
    INVX1 U10026 (.I(n20817), .ZN(n22898));
    INVX1 U10027 (.I(N4689), .ZN(n22899));
    NANDX1 U10028 (.A1(N10593), .A2(n13860), .ZN(N22900));
    NOR2X1 U10029 (.A1(N12778), .A2(n18064), .ZN(N22901));
    INVX1 U10030 (.I(N12041), .ZN(N22902));
    INVX1 U10031 (.I(N2760), .ZN(n22903));
    NOR2X1 U10032 (.A1(n18403), .A2(N6758), .ZN(n22904));
    INVX1 U10033 (.I(N6426), .ZN(n22905));
    NANDX1 U10034 (.A1(N8559), .A2(N5523), .ZN(n22906));
    INVX1 U10035 (.I(N4622), .ZN(n22907));
    INVX1 U10036 (.I(N1466), .ZN(n22908));
    NANDX1 U10037 (.A1(N11428), .A2(N3908), .ZN(n22909));
    INVX1 U10038 (.I(n13425), .ZN(n22910));
    NOR2X1 U10039 (.A1(n13511), .A2(N8410), .ZN(N22911));
    NANDX1 U10040 (.A1(n14583), .A2(n13545), .ZN(n22912));
    NANDX1 U10041 (.A1(n20093), .A2(N5092), .ZN(n22913));
    INVX1 U10042 (.I(n15491), .ZN(N22914));
    INVX1 U10043 (.I(N9771), .ZN(n22915));
    INVX1 U10044 (.I(n13338), .ZN(N22916));
    NANDX1 U10045 (.A1(n19550), .A2(n14282), .ZN(n22917));
    NOR2X1 U10046 (.A1(n17752), .A2(N1610), .ZN(N22918));
    NOR2X1 U10047 (.A1(N9147), .A2(N773), .ZN(n22919));
    NOR2X1 U10048 (.A1(N10612), .A2(n13156), .ZN(N22920));
    NOR2X1 U10049 (.A1(N9061), .A2(N392), .ZN(n22921));
    NOR2X1 U10050 (.A1(N1311), .A2(n13902), .ZN(N22922));
    INVX1 U10051 (.I(n14021), .ZN(n22923));
    NOR2X1 U10052 (.A1(N1596), .A2(n19360), .ZN(n22924));
    INVX1 U10053 (.I(N1229), .ZN(n22925));
    INVX1 U10054 (.I(N10691), .ZN(n22926));
    NANDX1 U10055 (.A1(n20386), .A2(N2253), .ZN(n22927));
    INVX1 U10056 (.I(N640), .ZN(n22928));
    NANDX1 U10057 (.A1(n13833), .A2(N8549), .ZN(n22929));
    INVX1 U10058 (.I(n15443), .ZN(n22930));
    NANDX1 U10059 (.A1(N782), .A2(N10757), .ZN(n22931));
    INVX1 U10060 (.I(N5936), .ZN(n22932));
    INVX1 U10061 (.I(N1824), .ZN(n22933));
    INVX1 U10062 (.I(n18845), .ZN(N22934));
    INVX1 U10063 (.I(N10848), .ZN(n22935));
    NOR2X1 U10064 (.A1(N11978), .A2(n19410), .ZN(n22936));
    INVX1 U10065 (.I(n13573), .ZN(n22937));
    NANDX1 U10066 (.A1(N8512), .A2(n14802), .ZN(n22938));
    NOR2X1 U10067 (.A1(n19202), .A2(N6474), .ZN(n22939));
    NANDX1 U10068 (.A1(n15997), .A2(N6025), .ZN(n22940));
    NANDX1 U10069 (.A1(N11111), .A2(n19858), .ZN(N22941));
    NOR2X1 U10070 (.A1(N2746), .A2(N8612), .ZN(N22942));
    INVX1 U10071 (.I(n19300), .ZN(n22943));
    INVX1 U10072 (.I(N8561), .ZN(n22944));
    NANDX1 U10073 (.A1(N11134), .A2(N4926), .ZN(n22945));
    NOR2X1 U10074 (.A1(N8748), .A2(N7622), .ZN(n22946));
    NANDX1 U10075 (.A1(n20264), .A2(n19599), .ZN(N22947));
    NOR2X1 U10076 (.A1(N6887), .A2(N11941), .ZN(n22948));
    NOR2X1 U10077 (.A1(n15398), .A2(N54), .ZN(n22949));
    NOR2X1 U10078 (.A1(N7911), .A2(N1069), .ZN(n22950));
    NOR2X1 U10079 (.A1(N2677), .A2(N7094), .ZN(N22951));
    NANDX1 U10080 (.A1(N8329), .A2(N263), .ZN(n22952));
    INVX1 U10081 (.I(N5617), .ZN(n22953));
    INVX1 U10082 (.I(N4384), .ZN(n22954));
    INVX1 U10083 (.I(N1553), .ZN(N22955));
    NOR2X1 U10084 (.A1(N2232), .A2(N12686), .ZN(n22956));
    NOR2X1 U10085 (.A1(N10315), .A2(n15976), .ZN(n22957));
    NANDX1 U10086 (.A1(N2558), .A2(N9551), .ZN(n22958));
    NANDX1 U10087 (.A1(n14211), .A2(n16437), .ZN(N22959));
    NOR2X1 U10088 (.A1(n16714), .A2(N5146), .ZN(n22960));
    INVX1 U10089 (.I(N4910), .ZN(n22961));
    NANDX1 U10090 (.A1(n15089), .A2(N9499), .ZN(n22962));
    NANDX1 U10091 (.A1(n16724), .A2(N4432), .ZN(n22963));
    NOR2X1 U10092 (.A1(n16986), .A2(N9172), .ZN(n22964));
    NOR2X1 U10093 (.A1(n20401), .A2(n13555), .ZN(n22965));
    NOR2X1 U10094 (.A1(n16495), .A2(n15582), .ZN(n22966));
    NANDX1 U10095 (.A1(N7951), .A2(N6763), .ZN(n22967));
    INVX1 U10096 (.I(n18468), .ZN(N22968));
    NOR2X1 U10097 (.A1(N5403), .A2(N6788), .ZN(n22969));
    NANDX1 U10098 (.A1(n19613), .A2(N1994), .ZN(n22970));
    INVX1 U10099 (.I(n15096), .ZN(n22971));
    NANDX1 U10100 (.A1(N8887), .A2(n14548), .ZN(n22972));
    INVX1 U10101 (.I(n18517), .ZN(n22973));
    NOR2X1 U10102 (.A1(n19552), .A2(n14010), .ZN(n22974));
    INVX1 U10103 (.I(N11467), .ZN(n22975));
    NOR2X1 U10104 (.A1(N5503), .A2(N8997), .ZN(n22976));
    NOR2X1 U10105 (.A1(n13599), .A2(N4755), .ZN(n22977));
    NOR2X1 U10106 (.A1(N7951), .A2(N2743), .ZN(N22978));
    INVX1 U10107 (.I(N9255), .ZN(n22979));
    NANDX1 U10108 (.A1(n19701), .A2(N3902), .ZN(N22980));
    NANDX1 U10109 (.A1(n21030), .A2(N6033), .ZN(n22981));
    NANDX1 U10110 (.A1(N1793), .A2(N900), .ZN(n22982));
    NOR2X1 U10111 (.A1(N3473), .A2(N4329), .ZN(n22983));
    INVX1 U10112 (.I(n18208), .ZN(N22984));
    NOR2X1 U10113 (.A1(N9083), .A2(n16530), .ZN(n22985));
    NOR2X1 U10114 (.A1(N5414), .A2(N1308), .ZN(n22986));
    NANDX1 U10115 (.A1(N10916), .A2(N10304), .ZN(n22987));
    NOR2X1 U10116 (.A1(N3284), .A2(N9600), .ZN(n22988));
    NOR2X1 U10117 (.A1(N11234), .A2(N6885), .ZN(n22989));
    INVX1 U10118 (.I(n20488), .ZN(n22990));
    NANDX1 U10119 (.A1(N20), .A2(n18932), .ZN(N22991));
    INVX1 U10120 (.I(n21049), .ZN(n22992));
    INVX1 U10121 (.I(N5545), .ZN(n22993));
    NANDX1 U10122 (.A1(n20406), .A2(N8181), .ZN(N22994));
    NOR2X1 U10123 (.A1(N3504), .A2(n19906), .ZN(n22995));
    NOR2X1 U10124 (.A1(n20890), .A2(N7758), .ZN(n22996));
    INVX1 U10125 (.I(N9826), .ZN(N22997));
    NOR2X1 U10126 (.A1(N8980), .A2(N8527), .ZN(N22998));
    NOR2X1 U10127 (.A1(n13826), .A2(n21018), .ZN(n22999));
    INVX1 U10128 (.I(N2195), .ZN(N23000));
    NOR2X1 U10129 (.A1(N6457), .A2(N9079), .ZN(N23001));
    INVX1 U10130 (.I(N257), .ZN(n23002));
    NANDX1 U10131 (.A1(N12588), .A2(n19188), .ZN(n23003));
    NANDX1 U10132 (.A1(N12406), .A2(n17463), .ZN(n23004));
    NANDX1 U10133 (.A1(N8558), .A2(n16638), .ZN(n23005));
    INVX1 U10134 (.I(N8182), .ZN(n23006));
    INVX1 U10135 (.I(n19205), .ZN(N23007));
    NANDX1 U10136 (.A1(n14343), .A2(N275), .ZN(N23008));
    INVX1 U10137 (.I(n18710), .ZN(N23009));
    NOR2X1 U10138 (.A1(N10519), .A2(N6006), .ZN(n23010));
    NOR2X1 U10139 (.A1(n18886), .A2(N335), .ZN(n23011));
    INVX1 U10140 (.I(n15623), .ZN(n23012));
    NOR2X1 U10141 (.A1(N12522), .A2(n19243), .ZN(n23013));
    NOR2X1 U10142 (.A1(N12778), .A2(N8647), .ZN(n23014));
    NOR2X1 U10143 (.A1(N5277), .A2(N5139), .ZN(n23015));
    INVX1 U10144 (.I(N1510), .ZN(n23016));
    NANDX1 U10145 (.A1(N4095), .A2(N12689), .ZN(n23017));
    INVX1 U10146 (.I(N6818), .ZN(N23018));
    NANDX1 U10147 (.A1(n20220), .A2(N6143), .ZN(N23019));
    INVX1 U10148 (.I(n15036), .ZN(n23020));
    INVX1 U10149 (.I(N7047), .ZN(n23021));
    NOR2X1 U10150 (.A1(N12742), .A2(n13053), .ZN(n23022));
    NOR2X1 U10151 (.A1(N4940), .A2(N7929), .ZN(n23023));
    NOR2X1 U10152 (.A1(n20562), .A2(n13825), .ZN(n23024));
    INVX1 U10153 (.I(n13116), .ZN(n23025));
    INVX1 U10154 (.I(n17311), .ZN(N23026));
    NOR2X1 U10155 (.A1(n15421), .A2(n17129), .ZN(n23027));
    NOR2X1 U10156 (.A1(N10958), .A2(n18638), .ZN(N23028));
    NANDX1 U10157 (.A1(N9595), .A2(N10097), .ZN(N23029));
    NANDX1 U10158 (.A1(N10954), .A2(N10780), .ZN(n23030));
    NANDX1 U10159 (.A1(N11638), .A2(n20347), .ZN(n23031));
    INVX1 U10160 (.I(n19319), .ZN(N23032));
    NANDX1 U10161 (.A1(n13302), .A2(N5373), .ZN(n23033));
    INVX1 U10162 (.I(n20478), .ZN(n23034));
    NANDX1 U10163 (.A1(N456), .A2(n17947), .ZN(n23035));
    NANDX1 U10164 (.A1(N8822), .A2(n17022), .ZN(n23036));
    NANDX1 U10165 (.A1(n19879), .A2(N7644), .ZN(n23037));
    INVX1 U10166 (.I(n14069), .ZN(N23038));
    NANDX1 U10167 (.A1(N12586), .A2(N3797), .ZN(n23039));
    NOR2X1 U10168 (.A1(N9056), .A2(N7933), .ZN(n23040));
    INVX1 U10169 (.I(N6540), .ZN(n23041));
    NOR2X1 U10170 (.A1(N10909), .A2(N3014), .ZN(n23042));
    NOR2X1 U10171 (.A1(N4567), .A2(N9066), .ZN(n23043));
    NOR2X1 U10172 (.A1(N5271), .A2(n16909), .ZN(n23044));
    NOR2X1 U10173 (.A1(n19028), .A2(n16157), .ZN(n23045));
    INVX1 U10174 (.I(n14025), .ZN(n23046));
    NANDX1 U10175 (.A1(N5417), .A2(N1616), .ZN(n23047));
    INVX1 U10176 (.I(N11801), .ZN(n23048));
    NOR2X1 U10177 (.A1(N5391), .A2(n18716), .ZN(n23049));
    NOR2X1 U10178 (.A1(N8933), .A2(N10072), .ZN(n23050));
    NANDX1 U10179 (.A1(N9882), .A2(n19127), .ZN(n23051));
    INVX1 U10180 (.I(N10011), .ZN(n23052));
    NOR2X1 U10181 (.A1(N7342), .A2(n20919), .ZN(n23053));
    NANDX1 U10182 (.A1(N11177), .A2(n20027), .ZN(N23054));
    NANDX1 U10183 (.A1(n13101), .A2(N4067), .ZN(n23055));
    NOR2X1 U10184 (.A1(N9480), .A2(n17636), .ZN(N23056));
    NANDX1 U10185 (.A1(n16171), .A2(N10430), .ZN(N23057));
    NANDX1 U10186 (.A1(n16129), .A2(N6587), .ZN(N23058));
    NANDX1 U10187 (.A1(N1241), .A2(n17165), .ZN(N23059));
    INVX1 U10188 (.I(n19957), .ZN(n23060));
    INVX1 U10189 (.I(n20544), .ZN(n23061));
    NOR2X1 U10190 (.A1(N6563), .A2(N3737), .ZN(n23062));
    INVX1 U10191 (.I(N10791), .ZN(n23063));
    NANDX1 U10192 (.A1(n15985), .A2(n18132), .ZN(N23064));
    NANDX1 U10193 (.A1(n17976), .A2(N2621), .ZN(n23065));
    INVX1 U10194 (.I(n18116), .ZN(n23066));
    NOR2X1 U10195 (.A1(N5381), .A2(N8477), .ZN(n23067));
    NANDX1 U10196 (.A1(N1787), .A2(n14993), .ZN(N23068));
    NOR2X1 U10197 (.A1(N6758), .A2(N2236), .ZN(n23069));
    INVX1 U10198 (.I(N7887), .ZN(n23070));
    INVX1 U10199 (.I(N5363), .ZN(n23071));
    NANDX1 U10200 (.A1(n14610), .A2(n19861), .ZN(N23072));
    NOR2X1 U10201 (.A1(N8465), .A2(N1970), .ZN(n23073));
    NANDX1 U10202 (.A1(N12201), .A2(n18977), .ZN(n23074));
    NANDX1 U10203 (.A1(n20489), .A2(n13732), .ZN(n23075));
    NANDX1 U10204 (.A1(n17549), .A2(N5019), .ZN(N23076));
    NANDX1 U10205 (.A1(n18863), .A2(n17677), .ZN(n23077));
    NANDX1 U10206 (.A1(N3013), .A2(N4923), .ZN(n23078));
    NANDX1 U10207 (.A1(n20571), .A2(n14457), .ZN(n23079));
    INVX1 U10208 (.I(N641), .ZN(n23080));
    INVX1 U10209 (.I(n15475), .ZN(N23081));
    INVX1 U10210 (.I(n19691), .ZN(n23082));
    NANDX1 U10211 (.A1(N12347), .A2(N7612), .ZN(n23083));
    NANDX1 U10212 (.A1(n15517), .A2(n16076), .ZN(n23084));
    NANDX1 U10213 (.A1(n19791), .A2(N1588), .ZN(n23085));
    NANDX1 U10214 (.A1(n13625), .A2(n16618), .ZN(N23086));
    NANDX1 U10215 (.A1(N4360), .A2(n12936), .ZN(N23087));
    NOR2X1 U10216 (.A1(n13488), .A2(N10568), .ZN(n23088));
    INVX1 U10217 (.I(n17105), .ZN(n23089));
    NOR2X1 U10218 (.A1(N1698), .A2(n19234), .ZN(N23090));
    INVX1 U10219 (.I(N10696), .ZN(n23091));
    INVX1 U10220 (.I(N8103), .ZN(N23092));
    INVX1 U10221 (.I(n19373), .ZN(N23093));
    NANDX1 U10222 (.A1(n14932), .A2(n13522), .ZN(n23094));
    NOR2X1 U10223 (.A1(N1313), .A2(N6302), .ZN(n23095));
    INVX1 U10224 (.I(n17388), .ZN(n23096));
    NANDX1 U10225 (.A1(N10905), .A2(n18975), .ZN(n23097));
    NOR2X1 U10226 (.A1(N3299), .A2(n14362), .ZN(n23098));
    NANDX1 U10227 (.A1(N2200), .A2(N609), .ZN(n23099));
    NANDX1 U10228 (.A1(n15687), .A2(N11176), .ZN(n23100));
    NANDX1 U10229 (.A1(N6104), .A2(n19298), .ZN(N23101));
    NANDX1 U10230 (.A1(N4107), .A2(N72), .ZN(N23102));
    INVX1 U10231 (.I(N8005), .ZN(n23103));
    NOR2X1 U10232 (.A1(N3909), .A2(N6148), .ZN(n23104));
    INVX1 U10233 (.I(n18840), .ZN(n23105));
    INVX1 U10234 (.I(n16172), .ZN(n23106));
    INVX1 U10235 (.I(n20512), .ZN(n23107));
    NOR2X1 U10236 (.A1(N5394), .A2(n16104), .ZN(n23108));
    NOR2X1 U10237 (.A1(N3139), .A2(n19964), .ZN(n23109));
    NOR2X1 U10238 (.A1(N12042), .A2(n19134), .ZN(N23110));
    NOR2X1 U10239 (.A1(N12651), .A2(n18633), .ZN(N23111));
    INVX1 U10240 (.I(n18368), .ZN(N23112));
    INVX1 U10241 (.I(n13331), .ZN(n23113));
    NOR2X1 U10242 (.A1(N1962), .A2(N11979), .ZN(N23114));
    NANDX1 U10243 (.A1(n20942), .A2(n19984), .ZN(n23115));
    INVX1 U10244 (.I(n19392), .ZN(N23116));
    INVX1 U10245 (.I(N6418), .ZN(N23117));
    NANDX1 U10246 (.A1(n19111), .A2(n17131), .ZN(n23118));
    NOR2X1 U10247 (.A1(n12935), .A2(n18958), .ZN(n23119));
    NANDX1 U10248 (.A1(N7808), .A2(N10459), .ZN(n23120));
    NANDX1 U10249 (.A1(N1083), .A2(n21030), .ZN(N23121));
    NOR2X1 U10250 (.A1(n14758), .A2(N12571), .ZN(n23122));
    NANDX1 U10251 (.A1(N12160), .A2(n19798), .ZN(n23123));
    NANDX1 U10252 (.A1(n16150), .A2(N6440), .ZN(n23124));
    NOR2X1 U10253 (.A1(n18111), .A2(n18418), .ZN(n23125));
    INVX1 U10254 (.I(N12365), .ZN(N23126));
    INVX1 U10255 (.I(N6863), .ZN(n23127));
    NOR2X1 U10256 (.A1(N11155), .A2(N7822), .ZN(n23128));
    NANDX1 U10257 (.A1(N3578), .A2(N3723), .ZN(N23129));
    INVX1 U10258 (.I(n16512), .ZN(n23130));
    NOR2X1 U10259 (.A1(n16247), .A2(n18861), .ZN(n23131));
    INVX1 U10260 (.I(N3097), .ZN(n23132));
    NOR2X1 U10261 (.A1(n16564), .A2(n17761), .ZN(N23133));
    NOR2X1 U10262 (.A1(N7904), .A2(n18387), .ZN(n23134));
    NOR2X1 U10263 (.A1(N1013), .A2(n16151), .ZN(N23135));
    NANDX1 U10264 (.A1(N7452), .A2(N3661), .ZN(n23136));
    INVX1 U10265 (.I(n20412), .ZN(N23137));
    INVX1 U10266 (.I(n18879), .ZN(n23138));
    NOR2X1 U10267 (.A1(N3622), .A2(N8174), .ZN(n23139));
    NANDX1 U10268 (.A1(N11444), .A2(N9013), .ZN(n23140));
    INVX1 U10269 (.I(N9708), .ZN(N23141));
    NOR2X1 U10270 (.A1(n15449), .A2(N241), .ZN(N23142));
    NANDX1 U10271 (.A1(n13079), .A2(N1233), .ZN(n23143));
    INVX1 U10272 (.I(N6334), .ZN(n23144));
    NANDX1 U10273 (.A1(N4043), .A2(n19805), .ZN(n23145));
    NOR2X1 U10274 (.A1(N1200), .A2(n13289), .ZN(n23146));
    NANDX1 U10275 (.A1(n17350), .A2(N7150), .ZN(N23147));
    NOR2X1 U10276 (.A1(n15552), .A2(n13664), .ZN(N23148));
    NANDX1 U10277 (.A1(N12311), .A2(N11312), .ZN(n23149));
    NOR2X1 U10278 (.A1(n15933), .A2(n14028), .ZN(n23150));
    INVX1 U10279 (.I(N6146), .ZN(n23151));
    INVX1 U10280 (.I(N932), .ZN(n23152));
    NOR2X1 U10281 (.A1(N11209), .A2(N10922), .ZN(n23153));
    NOR2X1 U10282 (.A1(n15625), .A2(n18542), .ZN(n23154));
    NANDX1 U10283 (.A1(N1907), .A2(N3646), .ZN(n23155));
    INVX1 U10284 (.I(N491), .ZN(n23156));
    NOR2X1 U10285 (.A1(N1987), .A2(N1690), .ZN(N23157));
    NOR2X1 U10286 (.A1(N2011), .A2(n13581), .ZN(n23158));
    INVX1 U10287 (.I(n19801), .ZN(N23159));
    NOR2X1 U10288 (.A1(N4175), .A2(n20999), .ZN(n23160));
    INVX1 U10289 (.I(N10028), .ZN(n23161));
    NANDX1 U10290 (.A1(N9457), .A2(N2825), .ZN(n23162));
    NOR2X1 U10291 (.A1(n15602), .A2(n20406), .ZN(n23163));
    NOR2X1 U10292 (.A1(N4766), .A2(N4927), .ZN(n23164));
    NOR2X1 U10293 (.A1(n15400), .A2(n20551), .ZN(N23165));
    INVX1 U10294 (.I(N579), .ZN(n23166));
    NOR2X1 U10295 (.A1(N10290), .A2(N3554), .ZN(n23167));
    INVX1 U10296 (.I(N1593), .ZN(n23168));
    INVX1 U10297 (.I(n13721), .ZN(n23169));
    INVX1 U10298 (.I(N2093), .ZN(N23170));
    NANDX1 U10299 (.A1(N2152), .A2(N663), .ZN(n23171));
    NOR2X1 U10300 (.A1(N868), .A2(N432), .ZN(n23172));
    INVX1 U10301 (.I(N10896), .ZN(n23173));
    NANDX1 U10302 (.A1(N6037), .A2(n13720), .ZN(n23174));
    NANDX1 U10303 (.A1(N408), .A2(N7438), .ZN(n23175));
    NANDX1 U10304 (.A1(n20945), .A2(N12364), .ZN(n23176));
    NANDX1 U10305 (.A1(N9656), .A2(N11684), .ZN(n23177));
    NANDX1 U10306 (.A1(N10235), .A2(N1994), .ZN(N23178));
    INVX1 U10307 (.I(n13788), .ZN(n23179));
    NOR2X1 U10308 (.A1(N3896), .A2(n19328), .ZN(n23180));
    INVX1 U10309 (.I(N10079), .ZN(n23181));
    NANDX1 U10310 (.A1(N1669), .A2(N6772), .ZN(n23182));
    INVX1 U10311 (.I(N4725), .ZN(n23183));
    NANDX1 U10312 (.A1(n17056), .A2(n17077), .ZN(n23184));
    NANDX1 U10313 (.A1(n12974), .A2(N1883), .ZN(n23185));
    INVX1 U10314 (.I(n17288), .ZN(N23186));
    NOR2X1 U10315 (.A1(n13003), .A2(n14555), .ZN(n23187));
    NANDX1 U10316 (.A1(n19908), .A2(N5383), .ZN(N23188));
    NOR2X1 U10317 (.A1(N4903), .A2(N2855), .ZN(n23189));
    NANDX1 U10318 (.A1(N6896), .A2(n20930), .ZN(n23190));
    NOR2X1 U10319 (.A1(n15462), .A2(n19367), .ZN(n23191));
    NANDX1 U10320 (.A1(n16517), .A2(N8215), .ZN(n23192));
    INVX1 U10321 (.I(n18185), .ZN(n23193));
    INVX1 U10322 (.I(n12989), .ZN(N23194));
    NOR2X1 U10323 (.A1(n17168), .A2(N3356), .ZN(n23195));
    NANDX1 U10324 (.A1(n14472), .A2(n16329), .ZN(N23196));
    INVX1 U10325 (.I(n14579), .ZN(N23197));
    NOR2X1 U10326 (.A1(N6552), .A2(N894), .ZN(N23198));
    INVX1 U10327 (.I(n18869), .ZN(N23199));
    NOR2X1 U10328 (.A1(N5635), .A2(N3840), .ZN(n23200));
    NOR2X1 U10329 (.A1(N3032), .A2(n14816), .ZN(N23201));
    INVX1 U10330 (.I(N2731), .ZN(n23202));
    INVX1 U10331 (.I(N142), .ZN(n23203));
    NOR2X1 U10332 (.A1(N9066), .A2(n16659), .ZN(n23204));
    NANDX1 U10333 (.A1(N5429), .A2(N8155), .ZN(n23205));
    NOR2X1 U10334 (.A1(n12959), .A2(n20148), .ZN(n23206));
    NANDX1 U10335 (.A1(n16315), .A2(N6756), .ZN(n23207));
    NOR2X1 U10336 (.A1(N11413), .A2(n16477), .ZN(n23208));
    NANDX1 U10337 (.A1(n18341), .A2(n17570), .ZN(n23209));
    INVX1 U10338 (.I(n18593), .ZN(n23210));
    NANDX1 U10339 (.A1(N6456), .A2(n18769), .ZN(n23211));
    INVX1 U10340 (.I(N5471), .ZN(n23212));
    NOR2X1 U10341 (.A1(N1717), .A2(N11382), .ZN(n23213));
    INVX1 U10342 (.I(n14609), .ZN(N23214));
    INVX1 U10343 (.I(n14482), .ZN(n23215));
    NOR2X1 U10344 (.A1(n17265), .A2(n18105), .ZN(n23216));
    INVX1 U10345 (.I(N4190), .ZN(N23217));
    NANDX1 U10346 (.A1(n15373), .A2(n18879), .ZN(N23218));
    INVX1 U10347 (.I(N4999), .ZN(n23219));
    NANDX1 U10348 (.A1(N10529), .A2(N10953), .ZN(n23220));
    NANDX1 U10349 (.A1(n16521), .A2(N8063), .ZN(N23221));
    NANDX1 U10350 (.A1(N2176), .A2(n21197), .ZN(N23222));
    NOR2X1 U10351 (.A1(N8631), .A2(n13278), .ZN(N23223));
    INVX1 U10352 (.I(n14102), .ZN(N23224));
    INVX1 U10353 (.I(n15587), .ZN(N23225));
    INVX1 U10354 (.I(N11689), .ZN(n23226));
    INVX1 U10355 (.I(n20631), .ZN(n23227));
    INVX1 U10356 (.I(N5950), .ZN(N23228));
    INVX1 U10357 (.I(n17587), .ZN(n23229));
    NOR2X1 U10358 (.A1(n15397), .A2(N925), .ZN(n23230));
    INVX1 U10359 (.I(n13045), .ZN(N23231));
    NOR2X1 U10360 (.A1(n17818), .A2(N11990), .ZN(N23232));
    INVX1 U10361 (.I(N7540), .ZN(n23233));
    NOR2X1 U10362 (.A1(n14941), .A2(N10145), .ZN(n23234));
    INVX1 U10363 (.I(n17116), .ZN(n23235));
    NOR2X1 U10364 (.A1(n18224), .A2(n20289), .ZN(n23236));
    INVX1 U10365 (.I(N10864), .ZN(n23237));
    INVX1 U10366 (.I(N10547), .ZN(n23238));
    NOR2X1 U10367 (.A1(N1038), .A2(n16777), .ZN(n23239));
    NANDX1 U10368 (.A1(N438), .A2(n16259), .ZN(n23240));
    NANDX1 U10369 (.A1(N11645), .A2(N12615), .ZN(N23241));
    INVX1 U10370 (.I(N5811), .ZN(n23242));
    NANDX1 U10371 (.A1(N3712), .A2(n13397), .ZN(n23243));
    INVX1 U10372 (.I(N299), .ZN(N23244));
    NOR2X1 U10373 (.A1(n21082), .A2(N2381), .ZN(N23245));
    NANDX1 U10374 (.A1(N9334), .A2(N12525), .ZN(N23246));
    NOR2X1 U10375 (.A1(n20992), .A2(N11719), .ZN(N23247));
    INVX1 U10376 (.I(n20050), .ZN(n23248));
    NANDX1 U10377 (.A1(n14304), .A2(N6521), .ZN(n23249));
    INVX1 U10378 (.I(n14065), .ZN(n23250));
    NOR2X1 U10379 (.A1(N9053), .A2(n17333), .ZN(N23251));
    NANDX1 U10380 (.A1(n19853), .A2(N5321), .ZN(n23252));
    NOR2X1 U10381 (.A1(N5779), .A2(N11985), .ZN(n23253));
    NANDX1 U10382 (.A1(n13859), .A2(N10239), .ZN(n23254));
    INVX1 U10383 (.I(n15290), .ZN(n23255));
    INVX1 U10384 (.I(n21171), .ZN(n23256));
    NANDX1 U10385 (.A1(N7459), .A2(n20592), .ZN(n23257));
    INVX1 U10386 (.I(n14525), .ZN(n23258));
    INVX1 U10387 (.I(n13319), .ZN(N23259));
    NANDX1 U10388 (.A1(n20165), .A2(N6680), .ZN(n23260));
    NOR2X1 U10389 (.A1(n13238), .A2(N7742), .ZN(N23261));
    NOR2X1 U10390 (.A1(N6072), .A2(N9841), .ZN(N23262));
    NOR2X1 U10391 (.A1(N2175), .A2(N12378), .ZN(n23263));
    NOR2X1 U10392 (.A1(N2037), .A2(n21101), .ZN(n23264));
    NOR2X1 U10393 (.A1(N8563), .A2(N8946), .ZN(n23265));
    NANDX1 U10394 (.A1(n18801), .A2(N4730), .ZN(n23266));
    INVX1 U10395 (.I(N2650), .ZN(n23267));
    NANDX1 U10396 (.A1(n20387), .A2(N10108), .ZN(n23268));
    INVX1 U10397 (.I(N12714), .ZN(N23269));
    NANDX1 U10398 (.A1(n15297), .A2(n20575), .ZN(n23270));
    NOR2X1 U10399 (.A1(N8773), .A2(N6024), .ZN(n23271));
    NOR2X1 U10400 (.A1(N780), .A2(n13766), .ZN(n23272));
    NOR2X1 U10401 (.A1(N6852), .A2(n18148), .ZN(n23273));
    NOR2X1 U10402 (.A1(N3568), .A2(N9295), .ZN(n23274));
    NANDX1 U10403 (.A1(N5604), .A2(N3707), .ZN(n23275));
    NANDX1 U10404 (.A1(n14166), .A2(N7195), .ZN(n23276));
    NOR2X1 U10405 (.A1(N6279), .A2(N11924), .ZN(N23277));
    INVX1 U10406 (.I(N8928), .ZN(n23278));
    INVX1 U10407 (.I(n15237), .ZN(n23279));
    NOR2X1 U10408 (.A1(N9708), .A2(N1262), .ZN(N23280));
    NANDX1 U10409 (.A1(N3775), .A2(N606), .ZN(n23281));
    NANDX1 U10410 (.A1(N7089), .A2(N1172), .ZN(n23282));
    INVX1 U10411 (.I(N7869), .ZN(N23283));
    NOR2X1 U10412 (.A1(N5043), .A2(n14720), .ZN(n23284));
    NOR2X1 U10413 (.A1(N4294), .A2(n18287), .ZN(n23285));
    INVX1 U10414 (.I(N552), .ZN(n23286));
    NOR2X1 U10415 (.A1(N8481), .A2(N10513), .ZN(N23287));
    INVX1 U10416 (.I(n15675), .ZN(n23288));
    INVX1 U10417 (.I(N12187), .ZN(N23289));
    NANDX1 U10418 (.A1(N10739), .A2(n21114), .ZN(n23290));
    NOR2X1 U10419 (.A1(N4745), .A2(n13461), .ZN(n23291));
    INVX1 U10420 (.I(N6007), .ZN(n23292));
    NOR2X1 U10421 (.A1(N4297), .A2(N1154), .ZN(n23293));
    NANDX1 U10422 (.A1(N11386), .A2(N2325), .ZN(n23294));
    NOR2X1 U10423 (.A1(n19254), .A2(N11803), .ZN(n23295));
    INVX1 U10424 (.I(N7285), .ZN(n23296));
    NOR2X1 U10425 (.A1(N198), .A2(n20113), .ZN(N23297));
    NOR2X1 U10426 (.A1(N749), .A2(N11856), .ZN(n23298));
    NOR2X1 U10427 (.A1(N5804), .A2(n17764), .ZN(n23299));
    NOR2X1 U10428 (.A1(N462), .A2(N3263), .ZN(N23300));
    NANDX1 U10429 (.A1(N11201), .A2(n18918), .ZN(n23301));
    INVX1 U10430 (.I(N10487), .ZN(n23302));
    INVX1 U10431 (.I(N2373), .ZN(n23303));
    NOR2X1 U10432 (.A1(n20357), .A2(N6670), .ZN(n23304));
    INVX1 U10433 (.I(N1583), .ZN(n23305));
    INVX1 U10434 (.I(n14513), .ZN(n23306));
    NOR2X1 U10435 (.A1(N10620), .A2(n20858), .ZN(n23307));
    NOR2X1 U10436 (.A1(N12446), .A2(N12368), .ZN(n23308));
    NANDX1 U10437 (.A1(N11328), .A2(N8652), .ZN(n23309));
    INVX1 U10438 (.I(N1953), .ZN(n23310));
    NANDX1 U10439 (.A1(N10869), .A2(n14258), .ZN(n23311));
    NANDX1 U10440 (.A1(N5872), .A2(n17520), .ZN(N23312));
    NOR2X1 U10441 (.A1(N11614), .A2(n15208), .ZN(n23313));
    INVX1 U10442 (.I(N871), .ZN(n23314));
    INVX1 U10443 (.I(n16967), .ZN(N23315));
    NOR2X1 U10444 (.A1(n14565), .A2(N2406), .ZN(N23316));
    NOR2X1 U10445 (.A1(n16147), .A2(N9544), .ZN(n23317));
    NANDX1 U10446 (.A1(N8591), .A2(n14705), .ZN(n23318));
    NANDX1 U10447 (.A1(n18168), .A2(N5920), .ZN(n23319));
    NANDX1 U10448 (.A1(N1255), .A2(N11789), .ZN(N23320));
    INVX1 U10449 (.I(N6320), .ZN(n23321));
    INVX1 U10450 (.I(N8976), .ZN(n23322));
    NOR2X1 U10451 (.A1(N1310), .A2(N371), .ZN(n23323));
    NANDX1 U10452 (.A1(n13372), .A2(n18572), .ZN(N23324));
    NANDX1 U10453 (.A1(N1891), .A2(N11936), .ZN(n23325));
    INVX1 U10454 (.I(N1557), .ZN(n23326));
    INVX1 U10455 (.I(n20759), .ZN(n23327));
    NOR2X1 U10456 (.A1(N4619), .A2(N2392), .ZN(n23328));
    INVX1 U10457 (.I(n14162), .ZN(n23329));
    NANDX1 U10458 (.A1(N8712), .A2(N7636), .ZN(n23330));
    INVX1 U10459 (.I(N5650), .ZN(N23331));
    NOR2X1 U10460 (.A1(N12762), .A2(N6904), .ZN(n23332));
    INVX1 U10461 (.I(N2864), .ZN(n23333));
    INVX1 U10462 (.I(N6937), .ZN(n23334));
    INVX1 U10463 (.I(N3722), .ZN(n23335));
    INVX1 U10464 (.I(N6751), .ZN(N23336));
    NANDX1 U10465 (.A1(n16159), .A2(N4093), .ZN(n23337));
    NOR2X1 U10466 (.A1(n18049), .A2(N10570), .ZN(n23338));
    NOR2X1 U10467 (.A1(n14148), .A2(n18241), .ZN(n23339));
    INVX1 U10468 (.I(N9039), .ZN(n23340));
    NOR2X1 U10469 (.A1(n13392), .A2(N9160), .ZN(n23341));
    NOR2X1 U10470 (.A1(N6470), .A2(n17872), .ZN(n23342));
    NOR2X1 U10471 (.A1(n16550), .A2(n18063), .ZN(n23343));
    NANDX1 U10472 (.A1(N8081), .A2(n19508), .ZN(n23344));
    NANDX1 U10473 (.A1(N10944), .A2(N6042), .ZN(n23345));
    NOR2X1 U10474 (.A1(n17324), .A2(N4305), .ZN(n23346));
    INVX1 U10475 (.I(n18617), .ZN(n23347));
    INVX1 U10476 (.I(N2681), .ZN(n23348));
    NOR2X1 U10477 (.A1(N7014), .A2(n20729), .ZN(N23349));
    INVX1 U10478 (.I(n18485), .ZN(n23350));
    INVX1 U10479 (.I(N3600), .ZN(N23351));
    NANDX1 U10480 (.A1(n17226), .A2(n15542), .ZN(n23352));
    NOR2X1 U10481 (.A1(n20928), .A2(N4643), .ZN(n23353));
    NANDX1 U10482 (.A1(n17569), .A2(N11693), .ZN(n23354));
    INVX1 U10483 (.I(N8943), .ZN(n23355));
    NANDX1 U10484 (.A1(N4826), .A2(N1762), .ZN(n23356));
    INVX1 U10485 (.I(N10311), .ZN(n23357));
    NANDX1 U10486 (.A1(N8601), .A2(N6405), .ZN(n23358));
    INVX1 U10487 (.I(n16352), .ZN(N23359));
    INVX1 U10488 (.I(N5586), .ZN(n23360));
    NANDX1 U10489 (.A1(n15583), .A2(N12599), .ZN(n23361));
    INVX1 U10490 (.I(N942), .ZN(n23362));
    NOR2X1 U10491 (.A1(N30), .A2(n20313), .ZN(n23363));
    INVX1 U10492 (.I(n17256), .ZN(n23364));
    NOR2X1 U10493 (.A1(N7608), .A2(N11495), .ZN(N23365));
    INVX1 U10494 (.I(N9034), .ZN(N23366));
    NANDX1 U10495 (.A1(N4270), .A2(N322), .ZN(N23367));
    NOR2X1 U10496 (.A1(n15336), .A2(n20919), .ZN(n23368));
    NANDX1 U10497 (.A1(n18972), .A2(N10000), .ZN(N23369));
    NOR2X1 U10498 (.A1(N884), .A2(N10946), .ZN(N23370));
    INVX1 U10499 (.I(N11777), .ZN(n23371));
    INVX1 U10500 (.I(n16739), .ZN(n23372));
    NANDX1 U10501 (.A1(N3630), .A2(N2650), .ZN(n23373));
    NANDX1 U10502 (.A1(n20343), .A2(N1587), .ZN(N23374));
    INVX1 U10503 (.I(n19425), .ZN(n23375));
    NOR2X1 U10504 (.A1(N2331), .A2(N7360), .ZN(N23376));
    INVX1 U10505 (.I(n13825), .ZN(n23377));
    INVX1 U10506 (.I(N4189), .ZN(N23378));
    INVX1 U10507 (.I(N4206), .ZN(n23379));
    INVX1 U10508 (.I(N827), .ZN(n23380));
    NOR2X1 U10509 (.A1(n19970), .A2(N8446), .ZN(n23381));
    NANDX1 U10510 (.A1(N8739), .A2(n18409), .ZN(n23382));
    INVX1 U10511 (.I(n14226), .ZN(n23383));
    NANDX1 U10512 (.A1(n13567), .A2(n18045), .ZN(n23384));
    NANDX1 U10513 (.A1(N12229), .A2(N444), .ZN(n23385));
    NANDX1 U10514 (.A1(N8191), .A2(n15328), .ZN(n23386));
    INVX1 U10515 (.I(n14497), .ZN(n23387));
    INVX1 U10516 (.I(N5937), .ZN(n23388));
    INVX1 U10517 (.I(n20881), .ZN(n23389));
    INVX1 U10518 (.I(N9422), .ZN(N23390));
    NANDX1 U10519 (.A1(n21052), .A2(n20162), .ZN(N23391));
    NOR2X1 U10520 (.A1(n14645), .A2(n20989), .ZN(N23392));
    NOR2X1 U10521 (.A1(n13384), .A2(N8204), .ZN(n23393));
    INVX1 U10522 (.I(n16665), .ZN(n23394));
    NOR2X1 U10523 (.A1(N4197), .A2(N9660), .ZN(N23395));
    INVX1 U10524 (.I(N12306), .ZN(n23396));
    NOR2X1 U10525 (.A1(N11494), .A2(N3304), .ZN(N23397));
    INVX1 U10526 (.I(N1609), .ZN(n23398));
    NANDX1 U10527 (.A1(n16788), .A2(n14540), .ZN(n23399));
    NANDX1 U10528 (.A1(N3621), .A2(n15019), .ZN(n23400));
    NOR2X1 U10529 (.A1(n19044), .A2(N10652), .ZN(n23401));
    NOR2X1 U10530 (.A1(n13172), .A2(N10473), .ZN(n23402));
    NOR2X1 U10531 (.A1(N6048), .A2(N3887), .ZN(n23403));
    NANDX1 U10532 (.A1(N7547), .A2(N11812), .ZN(n23404));
    NOR2X1 U10533 (.A1(N9954), .A2(N7246), .ZN(n23405));
    NANDX1 U10534 (.A1(n14150), .A2(N11448), .ZN(N23406));
    INVX1 U10535 (.I(n20997), .ZN(n23407));
    NOR2X1 U10536 (.A1(N3596), .A2(N3071), .ZN(n23408));
    NOR2X1 U10537 (.A1(N5205), .A2(N9107), .ZN(n23409));
    NANDX1 U10538 (.A1(n14286), .A2(N2951), .ZN(n23410));
    NANDX1 U10539 (.A1(N8074), .A2(n13621), .ZN(n23411));
    NOR2X1 U10540 (.A1(n18725), .A2(N7025), .ZN(n23412));
    NOR2X1 U10541 (.A1(N7967), .A2(n20590), .ZN(N23413));
    NANDX1 U10542 (.A1(N6395), .A2(N12683), .ZN(n23414));
    NANDX1 U10543 (.A1(n18207), .A2(N7521), .ZN(N23415));
    NANDX1 U10544 (.A1(n19994), .A2(n18056), .ZN(n23416));
    INVX1 U10545 (.I(N10211), .ZN(n23417));
    NOR2X1 U10546 (.A1(n18486), .A2(N1444), .ZN(n23418));
    NANDX1 U10547 (.A1(n16098), .A2(N9909), .ZN(n23419));
    NOR2X1 U10548 (.A1(N3974), .A2(n13930), .ZN(N23420));
    NANDX1 U10549 (.A1(N6924), .A2(n16114), .ZN(n23421));
    INVX1 U10550 (.I(n15086), .ZN(n23422));
    NOR2X1 U10551 (.A1(N6665), .A2(N880), .ZN(n23423));
    NOR2X1 U10552 (.A1(N9173), .A2(N239), .ZN(n23424));
    NANDX1 U10553 (.A1(N10110), .A2(N7463), .ZN(n23425));
    NOR2X1 U10554 (.A1(N1628), .A2(N9526), .ZN(n23426));
    NANDX1 U10555 (.A1(N391), .A2(N6351), .ZN(n23427));
    INVX1 U10556 (.I(N5144), .ZN(n23428));
    NOR2X1 U10557 (.A1(N10278), .A2(N1129), .ZN(n23429));
    NANDX1 U10558 (.A1(N5145), .A2(N11037), .ZN(n23430));
    NANDX1 U10559 (.A1(N3660), .A2(n19509), .ZN(n23431));
    NOR2X1 U10560 (.A1(N5125), .A2(N8934), .ZN(n23432));
    NOR2X1 U10561 (.A1(n20210), .A2(n19587), .ZN(N23433));
    NOR2X1 U10562 (.A1(n21090), .A2(N6406), .ZN(n23434));
    NANDX1 U10563 (.A1(n15870), .A2(N1524), .ZN(n23435));
    NANDX1 U10564 (.A1(N2103), .A2(N2175), .ZN(n23436));
    NANDX1 U10565 (.A1(N11628), .A2(N1936), .ZN(n23437));
    NOR2X1 U10566 (.A1(N12520), .A2(n20416), .ZN(n23438));
    NANDX1 U10567 (.A1(n18111), .A2(N9463), .ZN(N23439));
    NOR2X1 U10568 (.A1(N10766), .A2(N9149), .ZN(n23440));
    NOR2X1 U10569 (.A1(N11462), .A2(N12808), .ZN(n23441));
    NANDX1 U10570 (.A1(N7796), .A2(n17932), .ZN(n23442));
    INVX1 U10571 (.I(n13300), .ZN(n23443));
    NOR2X1 U10572 (.A1(N7823), .A2(N4237), .ZN(n23444));
    INVX1 U10573 (.I(N8770), .ZN(n23445));
    NANDX1 U10574 (.A1(N5952), .A2(N4835), .ZN(n23446));
    INVX1 U10575 (.I(N2596), .ZN(N23447));
    INVX1 U10576 (.I(N4580), .ZN(n23448));
    NANDX1 U10577 (.A1(N3487), .A2(N443), .ZN(n23449));
    NOR2X1 U10578 (.A1(n18444), .A2(N1448), .ZN(n23450));
    INVX1 U10579 (.I(N1219), .ZN(n23451));
    INVX1 U10580 (.I(N2242), .ZN(n23452));
    NOR2X1 U10581 (.A1(N5837), .A2(n13703), .ZN(n23453));
    NANDX1 U10582 (.A1(N911), .A2(n16041), .ZN(n23454));
    INVX1 U10583 (.I(N10377), .ZN(N23455));
    NANDX1 U10584 (.A1(N4641), .A2(N12741), .ZN(N23456));
    NOR2X1 U10585 (.A1(N10495), .A2(n16052), .ZN(N23457));
    NOR2X1 U10586 (.A1(N10989), .A2(n20887), .ZN(N23458));
    NOR2X1 U10587 (.A1(n13584), .A2(N1207), .ZN(N23459));
    NOR2X1 U10588 (.A1(N1119), .A2(n20465), .ZN(n23460));
    NANDX1 U10589 (.A1(n16944), .A2(n17679), .ZN(n23461));
    NOR2X1 U10590 (.A1(N8420), .A2(n18897), .ZN(n23462));
    INVX1 U10591 (.I(N10661), .ZN(n23463));
    NOR2X1 U10592 (.A1(n13795), .A2(n18905), .ZN(n23464));
    NANDX1 U10593 (.A1(n14705), .A2(n13715), .ZN(n23465));
    INVX1 U10594 (.I(n19624), .ZN(n23466));
    NOR2X1 U10595 (.A1(n18119), .A2(N5676), .ZN(n23467));
    INVX1 U10596 (.I(N7384), .ZN(N23468));
    INVX1 U10597 (.I(N2342), .ZN(n23469));
    NANDX1 U10598 (.A1(n15926), .A2(N851), .ZN(n23470));
    NANDX1 U10599 (.A1(N11674), .A2(n19712), .ZN(n23471));
    NANDX1 U10600 (.A1(N10909), .A2(N12327), .ZN(n23472));
    NOR2X1 U10601 (.A1(N1899), .A2(N932), .ZN(n23473));
    INVX1 U10602 (.I(n20795), .ZN(n23474));
    INVX1 U10603 (.I(N10262), .ZN(N23475));
    NOR2X1 U10604 (.A1(N1454), .A2(N7936), .ZN(n23476));
    NOR2X1 U10605 (.A1(n16158), .A2(N421), .ZN(n23477));
    NOR2X1 U10606 (.A1(n14551), .A2(n16786), .ZN(N23478));
    NOR2X1 U10607 (.A1(n14769), .A2(n18809), .ZN(n23479));
    INVX1 U10608 (.I(n15266), .ZN(n23480));
    NOR2X1 U10609 (.A1(n20946), .A2(N4503), .ZN(N23481));
    NANDX1 U10610 (.A1(n20755), .A2(n16176), .ZN(N23482));
    NOR2X1 U10611 (.A1(n16223), .A2(N396), .ZN(n23483));
    INVX1 U10612 (.I(N7405), .ZN(n23484));
    NOR2X1 U10613 (.A1(n17366), .A2(N7006), .ZN(n23485));
    NOR2X1 U10614 (.A1(N5025), .A2(n17267), .ZN(N23486));
    INVX1 U10615 (.I(N6478), .ZN(n23487));
    INVX1 U10616 (.I(n15510), .ZN(n23488));
    NOR2X1 U10617 (.A1(n14707), .A2(N3499), .ZN(N23489));
    NANDX1 U10618 (.A1(N4804), .A2(N9606), .ZN(n23490));
    NANDX1 U10619 (.A1(n18155), .A2(N12181), .ZN(n23491));
    NOR2X1 U10620 (.A1(N12616), .A2(N11896), .ZN(N23492));
    INVX1 U10621 (.I(N7928), .ZN(N23493));
    INVX1 U10622 (.I(N2374), .ZN(N23494));
    NOR2X1 U10623 (.A1(N955), .A2(N2770), .ZN(n23495));
    NOR2X1 U10624 (.A1(N8359), .A2(n20835), .ZN(n23496));
    NOR2X1 U10625 (.A1(N9907), .A2(N11777), .ZN(n23497));
    NANDX1 U10626 (.A1(N485), .A2(N4857), .ZN(n23498));
    NANDX1 U10627 (.A1(n20229), .A2(n20366), .ZN(n23499));
    NANDX1 U10628 (.A1(N8247), .A2(n18406), .ZN(n23500));
    INVX1 U10629 (.I(n13051), .ZN(n23501));
    NANDX1 U10630 (.A1(N8980), .A2(N9975), .ZN(n23502));
    NOR2X1 U10631 (.A1(n17364), .A2(N1360), .ZN(n23503));
    NANDX1 U10632 (.A1(N9020), .A2(N3830), .ZN(n23504));
    NOR2X1 U10633 (.A1(N11394), .A2(N10407), .ZN(n23505));
    INVX1 U10634 (.I(N8705), .ZN(N23506));
    NOR2X1 U10635 (.A1(N8527), .A2(N2851), .ZN(n23507));
    NOR2X1 U10636 (.A1(n18433), .A2(n14627), .ZN(N23508));
    INVX1 U10637 (.I(n13459), .ZN(n23509));
    INVX1 U10638 (.I(N1231), .ZN(n23510));
    INVX1 U10639 (.I(n13160), .ZN(n23511));
    INVX1 U10640 (.I(n15246), .ZN(n23512));
    NANDX1 U10641 (.A1(n16997), .A2(N1608), .ZN(n23513));
    NANDX1 U10642 (.A1(N4746), .A2(N11582), .ZN(n23514));
    INVX1 U10643 (.I(N880), .ZN(N23515));
    INVX1 U10644 (.I(N2640), .ZN(n23516));
    INVX1 U10645 (.I(N5855), .ZN(N23517));
    NOR2X1 U10646 (.A1(N10376), .A2(N10803), .ZN(n23518));
    INVX1 U10647 (.I(n13622), .ZN(n23519));
    NANDX1 U10648 (.A1(N10547), .A2(n16473), .ZN(n23520));
    NANDX1 U10649 (.A1(N2291), .A2(N9869), .ZN(N23521));
    NOR2X1 U10650 (.A1(n15750), .A2(N2664), .ZN(N23522));
    NANDX1 U10651 (.A1(N1519), .A2(N10365), .ZN(n23523));
    NANDX1 U10652 (.A1(n16764), .A2(n20700), .ZN(n23524));
    INVX1 U10653 (.I(n12914), .ZN(n23525));
    NANDX1 U10654 (.A1(N6553), .A2(n19037), .ZN(n23526));
    NOR2X1 U10655 (.A1(N1974), .A2(N5290), .ZN(n23527));
    INVX1 U10656 (.I(N6414), .ZN(N23528));
    NOR2X1 U10657 (.A1(N3175), .A2(N11332), .ZN(n23529));
    NANDX1 U10658 (.A1(N10653), .A2(N3723), .ZN(n23530));
    INVX1 U10659 (.I(n15742), .ZN(n23531));
    INVX1 U10660 (.I(N8879), .ZN(n23532));
    INVX1 U10661 (.I(N3376), .ZN(n23533));
    NANDX1 U10662 (.A1(N12551), .A2(N581), .ZN(n23534));
    NOR2X1 U10663 (.A1(n14069), .A2(N10945), .ZN(N23535));
    NOR2X1 U10664 (.A1(N4145), .A2(N4956), .ZN(n23536));
    INVX1 U10665 (.I(n17058), .ZN(N23537));
    NANDX1 U10666 (.A1(N5772), .A2(n14864), .ZN(n23538));
    NOR2X1 U10667 (.A1(N2287), .A2(n14696), .ZN(n23539));
    NOR2X1 U10668 (.A1(N3243), .A2(n14923), .ZN(N23540));
    INVX1 U10669 (.I(n14574), .ZN(n23541));
    INVX1 U10670 (.I(n13537), .ZN(n23542));
    NANDX1 U10671 (.A1(n17511), .A2(N8048), .ZN(n23543));
    INVX1 U10672 (.I(N5160), .ZN(n23544));
    NANDX1 U10673 (.A1(N9720), .A2(n17713), .ZN(n23545));
    NANDX1 U10674 (.A1(N10300), .A2(n19400), .ZN(n23546));
    INVX1 U10675 (.I(N14), .ZN(N23547));
    NANDX1 U10676 (.A1(N8925), .A2(N4970), .ZN(n23548));
    NANDX1 U10677 (.A1(n20524), .A2(N10135), .ZN(n23549));
    NOR2X1 U10678 (.A1(N8699), .A2(n13982), .ZN(n23550));
    NOR2X1 U10679 (.A1(n17936), .A2(n19150), .ZN(n23551));
    NANDX1 U10680 (.A1(N11629), .A2(N6262), .ZN(n23552));
    NOR2X1 U10681 (.A1(N10893), .A2(n19799), .ZN(n23553));
    NOR2X1 U10682 (.A1(N7173), .A2(N6616), .ZN(N23554));
    NOR2X1 U10683 (.A1(N6874), .A2(N11465), .ZN(n23555));
    NANDX1 U10684 (.A1(N3357), .A2(N2177), .ZN(n23556));
    NANDX1 U10685 (.A1(N1526), .A2(N6957), .ZN(n23557));
    INVX1 U10686 (.I(N7422), .ZN(N23558));
    INVX1 U10687 (.I(N6023), .ZN(N23559));
    INVX1 U10688 (.I(N9716), .ZN(N23560));
    NOR2X1 U10689 (.A1(N7652), .A2(n12956), .ZN(n23561));
    NANDX1 U10690 (.A1(n15368), .A2(N9662), .ZN(n23562));
    NOR2X1 U10691 (.A1(N10553), .A2(n15832), .ZN(N23563));
    NANDX1 U10692 (.A1(n14854), .A2(N5494), .ZN(n23564));
    NOR2X1 U10693 (.A1(n16220), .A2(N7208), .ZN(n23565));
    NOR2X1 U10694 (.A1(N2700), .A2(n14082), .ZN(n23566));
    NANDX1 U10695 (.A1(n20129), .A2(N11980), .ZN(N23567));
    INVX1 U10696 (.I(N5397), .ZN(n23568));
    INVX1 U10697 (.I(n17038), .ZN(n23569));
    NOR2X1 U10698 (.A1(n15468), .A2(N6230), .ZN(n23570));
    NANDX1 U10699 (.A1(N6774), .A2(N10487), .ZN(n23571));
    NANDX1 U10700 (.A1(N8968), .A2(N2213), .ZN(n23572));
    INVX1 U10701 (.I(N3105), .ZN(n23573));
    NANDX1 U10702 (.A1(N11618), .A2(N8199), .ZN(n23574));
    NANDX1 U10703 (.A1(n13792), .A2(N1822), .ZN(N23575));
    NANDX1 U10704 (.A1(N9075), .A2(N12583), .ZN(n23576));
    NOR2X1 U10705 (.A1(N10974), .A2(N9824), .ZN(n23577));
    NOR2X1 U10706 (.A1(n18880), .A2(N8722), .ZN(n23578));
    NANDX1 U10707 (.A1(N7731), .A2(n14118), .ZN(N23579));
    NOR2X1 U10708 (.A1(N3539), .A2(n20568), .ZN(n23580));
    NANDX1 U10709 (.A1(N4310), .A2(N6352), .ZN(n23581));
    INVX1 U10710 (.I(n14797), .ZN(n23582));
    NANDX1 U10711 (.A1(N9281), .A2(N11551), .ZN(n23583));
    NOR2X1 U10712 (.A1(N12385), .A2(N12508), .ZN(n23584));
    NOR2X1 U10713 (.A1(n20583), .A2(N8066), .ZN(n23585));
    NANDX1 U10714 (.A1(n16947), .A2(N3659), .ZN(n23586));
    NOR2X1 U10715 (.A1(N2841), .A2(N1001), .ZN(N23587));
    INVX1 U10716 (.I(N12665), .ZN(N23588));
    INVX1 U10717 (.I(N2812), .ZN(n23589));
    NANDX1 U10718 (.A1(N9139), .A2(N10542), .ZN(N23590));
    INVX1 U10719 (.I(n13900), .ZN(n23591));
    NOR2X1 U10720 (.A1(N2695), .A2(N7439), .ZN(N23592));
    INVX1 U10721 (.I(N3588), .ZN(n23593));
    NANDX1 U10722 (.A1(N1040), .A2(N6422), .ZN(N23594));
    INVX1 U10723 (.I(N7132), .ZN(n23595));
    INVX1 U10724 (.I(N2728), .ZN(n23596));
    NANDX1 U10725 (.A1(n17514), .A2(n17853), .ZN(N23597));
    INVX1 U10726 (.I(N8086), .ZN(n23598));
    INVX1 U10727 (.I(N4674), .ZN(n23599));
    NANDX1 U10728 (.A1(N10951), .A2(N216), .ZN(N23600));
    NOR2X1 U10729 (.A1(N2385), .A2(N12640), .ZN(n23601));
    NANDX1 U10730 (.A1(n18313), .A2(n16321), .ZN(N23602));
    INVX1 U10731 (.I(N440), .ZN(n23603));
    NANDX1 U10732 (.A1(N8181), .A2(n18906), .ZN(n23604));
    INVX1 U10733 (.I(n21112), .ZN(n23605));
    INVX1 U10734 (.I(n13264), .ZN(n23606));
    INVX1 U10735 (.I(N2226), .ZN(N23607));
    INVX1 U10736 (.I(N2594), .ZN(n23608));
    INVX1 U10737 (.I(N877), .ZN(n23609));
    NOR2X1 U10738 (.A1(N12554), .A2(n18729), .ZN(N23610));
    NOR2X1 U10739 (.A1(n15181), .A2(N5609), .ZN(N23611));
    INVX1 U10740 (.I(n17455), .ZN(n23612));
    INVX1 U10741 (.I(N1447), .ZN(N23613));
    NOR2X1 U10742 (.A1(N8028), .A2(N8629), .ZN(n23614));
    INVX1 U10743 (.I(n20882), .ZN(n23615));
    INVX1 U10744 (.I(n13467), .ZN(n23616));
    NOR2X1 U10745 (.A1(N7250), .A2(n16189), .ZN(n23617));
    INVX1 U10746 (.I(N12761), .ZN(n23618));
    INVX1 U10747 (.I(n14800), .ZN(n23619));
    INVX1 U10748 (.I(N6074), .ZN(n23620));
    INVX1 U10749 (.I(N2943), .ZN(n23621));
    NANDX1 U10750 (.A1(N6606), .A2(n19591), .ZN(N23622));
    INVX1 U10751 (.I(n13701), .ZN(n23623));
    NOR2X1 U10752 (.A1(N6226), .A2(N7652), .ZN(n23624));
    NOR2X1 U10753 (.A1(N1999), .A2(n19648), .ZN(n23625));
    NOR2X1 U10754 (.A1(n19217), .A2(N2079), .ZN(n23626));
    NANDX1 U10755 (.A1(N1157), .A2(n15986), .ZN(n23627));
    NANDX1 U10756 (.A1(N4875), .A2(N2764), .ZN(n23628));
    INVX1 U10757 (.I(N6666), .ZN(n23629));
    NANDX1 U10758 (.A1(n17498), .A2(n19427), .ZN(N23630));
    NANDX1 U10759 (.A1(N5609), .A2(n18762), .ZN(n23631));
    NANDX1 U10760 (.A1(n17175), .A2(N474), .ZN(n23632));
    NOR2X1 U10761 (.A1(n18323), .A2(n20064), .ZN(n23633));
    INVX1 U10762 (.I(N5335), .ZN(N23634));
    NANDX1 U10763 (.A1(N6818), .A2(N7528), .ZN(n23635));
    NANDX1 U10764 (.A1(N3358), .A2(N5946), .ZN(N23636));
    NOR2X1 U10765 (.A1(n17117), .A2(N8024), .ZN(n23637));
    NANDX1 U10766 (.A1(n18273), .A2(n18551), .ZN(n23638));
    INVX1 U10767 (.I(n17690), .ZN(n23639));
    NANDX1 U10768 (.A1(N4401), .A2(N3125), .ZN(n23640));
    NOR2X1 U10769 (.A1(N669), .A2(N1321), .ZN(N23641));
    NANDX1 U10770 (.A1(N6277), .A2(n20083), .ZN(n23642));
    INVX1 U10771 (.I(n17994), .ZN(n23643));
    NANDX1 U10772 (.A1(n16928), .A2(n15086), .ZN(n23644));
    NANDX1 U10773 (.A1(n17520), .A2(n20420), .ZN(n23645));
    INVX1 U10774 (.I(n18880), .ZN(N23646));
    NOR2X1 U10775 (.A1(n14493), .A2(N1007), .ZN(n23647));
    NOR2X1 U10776 (.A1(n17157), .A2(n18123), .ZN(n23648));
    INVX1 U10777 (.I(N2810), .ZN(n23649));
    NOR2X1 U10778 (.A1(N12548), .A2(N3250), .ZN(n23650));
    NANDX1 U10779 (.A1(N12632), .A2(N7651), .ZN(n23651));
    INVX1 U10780 (.I(N4980), .ZN(n23652));
    NOR2X1 U10781 (.A1(N10612), .A2(N11118), .ZN(n23653));
    NOR2X1 U10782 (.A1(N4006), .A2(n20745), .ZN(n23654));
    NOR2X1 U10783 (.A1(n19103), .A2(N10984), .ZN(N23655));
    INVX1 U10784 (.I(N888), .ZN(N23656));
    NOR2X1 U10785 (.A1(n14717), .A2(n14367), .ZN(n23657));
    INVX1 U10786 (.I(N204), .ZN(n23658));
    INVX1 U10787 (.I(N471), .ZN(n23659));
    INVX1 U10788 (.I(n19327), .ZN(N23660));
    INVX1 U10789 (.I(N1405), .ZN(N23661));
    NOR2X1 U10790 (.A1(N7071), .A2(n13952), .ZN(n23662));
    NANDX1 U10791 (.A1(n13237), .A2(n21126), .ZN(n23663));
    INVX1 U10792 (.I(N1297), .ZN(n23664));
    NOR2X1 U10793 (.A1(N9208), .A2(N6450), .ZN(n23665));
    NANDX1 U10794 (.A1(n12886), .A2(N10455), .ZN(n23666));
    INVX1 U10795 (.I(n13328), .ZN(N23667));
    NOR2X1 U10796 (.A1(n21032), .A2(n13082), .ZN(n23668));
    NOR2X1 U10797 (.A1(N1617), .A2(N1110), .ZN(n23669));
    NANDX1 U10798 (.A1(N6539), .A2(n17085), .ZN(n23670));
    NOR2X1 U10799 (.A1(N7009), .A2(N3262), .ZN(N23671));
    NOR2X1 U10800 (.A1(n20144), .A2(n20438), .ZN(n23672));
    INVX1 U10801 (.I(N5984), .ZN(n23673));
    NANDX1 U10802 (.A1(N1618), .A2(n13762), .ZN(n23674));
    NANDX1 U10803 (.A1(N2507), .A2(n15059), .ZN(N23675));
    INVX1 U10804 (.I(N6256), .ZN(n23676));
    NANDX1 U10805 (.A1(n17546), .A2(n19141), .ZN(n23677));
    NANDX1 U10806 (.A1(N6363), .A2(N11238), .ZN(n23678));
    NANDX1 U10807 (.A1(N706), .A2(n18862), .ZN(n23679));
    NANDX1 U10808 (.A1(N2322), .A2(n14513), .ZN(N23680));
    NANDX1 U10809 (.A1(N3402), .A2(N10368), .ZN(n23681));
    INVX1 U10810 (.I(N4953), .ZN(n23682));
    NOR2X1 U10811 (.A1(N9268), .A2(N3866), .ZN(n23683));
    NOR2X1 U10812 (.A1(N12188), .A2(N4392), .ZN(n23684));
    NANDX1 U10813 (.A1(n13805), .A2(N12695), .ZN(N23685));
    INVX1 U10814 (.I(N10853), .ZN(n23686));
    NOR2X1 U10815 (.A1(N8458), .A2(n17108), .ZN(n23687));
    NANDX1 U10816 (.A1(N4773), .A2(N9560), .ZN(n23688));
    INVX1 U10817 (.I(N5677), .ZN(n23689));
    NOR2X1 U10818 (.A1(n19616), .A2(N6383), .ZN(n23690));
    INVX1 U10819 (.I(n15141), .ZN(n23691));
    NOR2X1 U10820 (.A1(N6253), .A2(N2101), .ZN(n23692));
    NOR2X1 U10821 (.A1(N11162), .A2(N3896), .ZN(N23693));
    NOR2X1 U10822 (.A1(N3561), .A2(N7705), .ZN(n23694));
    NANDX1 U10823 (.A1(N10939), .A2(n14434), .ZN(n23695));
    NOR2X1 U10824 (.A1(N10246), .A2(N1550), .ZN(n23696));
    NANDX1 U10825 (.A1(N6233), .A2(N12402), .ZN(n23697));
    INVX1 U10826 (.I(n14690), .ZN(n23698));
    NOR2X1 U10827 (.A1(n13125), .A2(n19462), .ZN(N23699));
    NOR2X1 U10828 (.A1(N8825), .A2(n19680), .ZN(N23700));
    NANDX1 U10829 (.A1(N1752), .A2(N4832), .ZN(N23701));
    NOR2X1 U10830 (.A1(N11435), .A2(N2620), .ZN(N23702));
    NOR2X1 U10831 (.A1(n13535), .A2(N3809), .ZN(n23703));
    INVX1 U10832 (.I(N11972), .ZN(n23704));
    NANDX1 U10833 (.A1(N8287), .A2(n14218), .ZN(N23705));
    NOR2X1 U10834 (.A1(n19225), .A2(N7421), .ZN(n23706));
    INVX1 U10835 (.I(N2782), .ZN(n23707));
    NOR2X1 U10836 (.A1(N7468), .A2(N9014), .ZN(N23708));
    INVX1 U10837 (.I(N3478), .ZN(n23709));
    NOR2X1 U10838 (.A1(N2961), .A2(n16603), .ZN(n23710));
    INVX1 U10839 (.I(n15341), .ZN(n23711));
    NOR2X1 U10840 (.A1(n14926), .A2(n16371), .ZN(N23712));
    NANDX1 U10841 (.A1(n14299), .A2(N9142), .ZN(n23713));
    INVX1 U10842 (.I(N11460), .ZN(n23714));
    NOR2X1 U10843 (.A1(n14543), .A2(N9810), .ZN(n23715));
    INVX1 U10844 (.I(n21057), .ZN(n23716));
    NOR2X1 U10845 (.A1(n15720), .A2(n14044), .ZN(n23717));
    NOR2X1 U10846 (.A1(N8256), .A2(N235), .ZN(n23718));
    INVX1 U10847 (.I(N5580), .ZN(n23719));
    INVX1 U10848 (.I(n16641), .ZN(n23720));
    NANDX1 U10849 (.A1(N3887), .A2(n20118), .ZN(n23721));
    NANDX1 U10850 (.A1(N1389), .A2(N10032), .ZN(n23722));
    NOR2X1 U10851 (.A1(n16729), .A2(N3313), .ZN(n23723));
    INVX1 U10852 (.I(N6412), .ZN(n23724));
    NOR2X1 U10853 (.A1(n14245), .A2(n15553), .ZN(n23725));
    INVX1 U10854 (.I(N4474), .ZN(n23726));
    NOR2X1 U10855 (.A1(n13895), .A2(N8826), .ZN(n23727));
    NOR2X1 U10856 (.A1(n13721), .A2(N1896), .ZN(n23728));
    INVX1 U10857 (.I(N1077), .ZN(n23729));
    NOR2X1 U10858 (.A1(N1748), .A2(N1311), .ZN(n23730));
    NOR2X1 U10859 (.A1(N1869), .A2(N5056), .ZN(n23731));
    NANDX1 U10860 (.A1(N11003), .A2(N3484), .ZN(N23732));
    NOR2X1 U10861 (.A1(N11694), .A2(N4873), .ZN(n23733));
    NOR2X1 U10862 (.A1(N7631), .A2(n16143), .ZN(n23734));
    NANDX1 U10863 (.A1(N7576), .A2(N1324), .ZN(n23735));
    NANDX1 U10864 (.A1(N590), .A2(N11418), .ZN(n23736));
    NANDX1 U10865 (.A1(n20836), .A2(N8446), .ZN(n23737));
    NANDX1 U10866 (.A1(N8431), .A2(n12907), .ZN(N23738));
    INVX1 U10867 (.I(N4868), .ZN(N23739));
    NANDX1 U10868 (.A1(N9001), .A2(n19188), .ZN(n23740));
    INVX1 U10869 (.I(N4853), .ZN(n23741));
    NANDX1 U10870 (.A1(n20327), .A2(N4451), .ZN(n23742));
    INVX1 U10871 (.I(N10100), .ZN(n23743));
    INVX1 U10872 (.I(n15683), .ZN(n23744));
    NANDX1 U10873 (.A1(N7348), .A2(N11358), .ZN(n23745));
    NANDX1 U10874 (.A1(n18033), .A2(N4888), .ZN(N23746));
    NANDX1 U10875 (.A1(n13898), .A2(n17991), .ZN(n23747));
    INVX1 U10876 (.I(N4086), .ZN(n23748));
    INVX1 U10877 (.I(n20819), .ZN(N23749));
    INVX1 U10878 (.I(n19193), .ZN(n23750));
    NANDX1 U10879 (.A1(n19979), .A2(N5887), .ZN(n23751));
    INVX1 U10880 (.I(n20919), .ZN(n23752));
    NANDX1 U10881 (.A1(N5386), .A2(n18147), .ZN(n23753));
    INVX1 U10882 (.I(N5605), .ZN(n23754));
    INVX1 U10883 (.I(n18732), .ZN(N23755));
    NOR2X1 U10884 (.A1(N655), .A2(n21208), .ZN(n23756));
    NOR2X1 U10885 (.A1(n16989), .A2(N1867), .ZN(n23757));
    INVX1 U10886 (.I(n14266), .ZN(N23758));
    NOR2X1 U10887 (.A1(N3278), .A2(n19118), .ZN(N23759));
    NANDX1 U10888 (.A1(n15810), .A2(n19101), .ZN(N23760));
    NANDX1 U10889 (.A1(n14110), .A2(n18690), .ZN(n23761));
    NOR2X1 U10890 (.A1(N12072), .A2(N20), .ZN(n23762));
    NANDX1 U10891 (.A1(n17959), .A2(N1990), .ZN(n23763));
    NANDX1 U10892 (.A1(N6158), .A2(N1917), .ZN(n23764));
    INVX1 U10893 (.I(n20439), .ZN(n23765));
    INVX1 U10894 (.I(N9632), .ZN(n23766));
    NANDX1 U10895 (.A1(N5560), .A2(N4828), .ZN(n23767));
    INVX1 U10896 (.I(n19281), .ZN(n23768));
    NOR2X1 U10897 (.A1(n14326), .A2(N12213), .ZN(N23769));
    NANDX1 U10898 (.A1(N7537), .A2(N10032), .ZN(N23770));
    NANDX1 U10899 (.A1(n20103), .A2(N4611), .ZN(N23771));
    NOR2X1 U10900 (.A1(N10066), .A2(n13263), .ZN(N23772));
    NANDX1 U10901 (.A1(N12559), .A2(N4104), .ZN(n23773));
    NOR2X1 U10902 (.A1(n13801), .A2(n16604), .ZN(N23774));
    NOR2X1 U10903 (.A1(N9273), .A2(N1531), .ZN(n23775));
    INVX1 U10904 (.I(n17434), .ZN(n23776));
    NANDX1 U10905 (.A1(N3141), .A2(N377), .ZN(n23777));
    NOR2X1 U10906 (.A1(N3242), .A2(N5205), .ZN(N23778));
    INVX1 U10907 (.I(n17064), .ZN(n23779));
    NANDX1 U10908 (.A1(N2402), .A2(N8046), .ZN(n23780));
    INVX1 U10909 (.I(N9938), .ZN(n23781));
    INVX1 U10910 (.I(N1234), .ZN(n23782));
    NOR2X1 U10911 (.A1(n17230), .A2(N6384), .ZN(N23783));
    INVX1 U10912 (.I(N9262), .ZN(n23784));
    NANDX1 U10913 (.A1(n20518), .A2(n13365), .ZN(n23785));
    INVX1 U10914 (.I(N7630), .ZN(n23786));
    NANDX1 U10915 (.A1(n21097), .A2(N11445), .ZN(n23787));
    NOR2X1 U10916 (.A1(n16716), .A2(N7648), .ZN(n23788));
    INVX1 U10917 (.I(n14398), .ZN(n23789));
    NOR2X1 U10918 (.A1(N2397), .A2(n17640), .ZN(n23790));
    NANDX1 U10919 (.A1(N11703), .A2(n13473), .ZN(N23791));
    INVX1 U10920 (.I(N8647), .ZN(n23792));
    NOR2X1 U10921 (.A1(N2055), .A2(n13126), .ZN(n23793));
    NOR2X1 U10922 (.A1(n19060), .A2(n16478), .ZN(n23794));
    NOR2X1 U10923 (.A1(N4214), .A2(n18978), .ZN(N23795));
    NANDX1 U10924 (.A1(N7749), .A2(n18265), .ZN(n23796));
    NOR2X1 U10925 (.A1(N8455), .A2(N4665), .ZN(n23797));
    INVX1 U10926 (.I(N8321), .ZN(n23798));
    INVX1 U10927 (.I(N7476), .ZN(n23799));
    INVX1 U10928 (.I(n18298), .ZN(N23800));
    NOR2X1 U10929 (.A1(n18204), .A2(N5091), .ZN(n23801));
    INVX1 U10930 (.I(N9155), .ZN(n23802));
    INVX1 U10931 (.I(N10751), .ZN(N23803));
    NANDX1 U10932 (.A1(n20962), .A2(n19397), .ZN(n23804));
    NANDX1 U10933 (.A1(N1787), .A2(N11292), .ZN(N23805));
    INVX1 U10934 (.I(n15388), .ZN(n23806));
    NOR2X1 U10935 (.A1(N7124), .A2(n19601), .ZN(n23807));
    NOR2X1 U10936 (.A1(n14374), .A2(N6119), .ZN(n23808));
    NOR2X1 U10937 (.A1(n13759), .A2(N9115), .ZN(n23809));
    NANDX1 U10938 (.A1(n16424), .A2(n17436), .ZN(n23810));
    NANDX1 U10939 (.A1(N2670), .A2(n15784), .ZN(n23811));
    INVX1 U10940 (.I(N4779), .ZN(n23812));
    NANDX1 U10941 (.A1(N2419), .A2(n19598), .ZN(n23813));
    INVX1 U10942 (.I(N9821), .ZN(n23814));
    NOR2X1 U10943 (.A1(n17851), .A2(N9552), .ZN(N23815));
    NOR2X1 U10944 (.A1(N3162), .A2(N5880), .ZN(n23816));
    NANDX1 U10945 (.A1(N6837), .A2(N38), .ZN(N23817));
    INVX1 U10946 (.I(N8502), .ZN(n23818));
    NOR2X1 U10947 (.A1(N2110), .A2(n17418), .ZN(N23819));
    NANDX1 U10948 (.A1(n13745), .A2(N9946), .ZN(n23820));
    INVX1 U10949 (.I(N3355), .ZN(n23821));
    INVX1 U10950 (.I(n20160), .ZN(n23822));
    NANDX1 U10951 (.A1(N2351), .A2(n14713), .ZN(n23823));
    NANDX1 U10952 (.A1(N1671), .A2(N782), .ZN(N23824));
    INVX1 U10953 (.I(N38), .ZN(n23825));
    INVX1 U10954 (.I(N7723), .ZN(n23826));
    NOR2X1 U10955 (.A1(N8397), .A2(N11817), .ZN(n23827));
    NANDX1 U10956 (.A1(N6100), .A2(N12238), .ZN(n23828));
    NOR2X1 U10957 (.A1(n12936), .A2(N12275), .ZN(n23829));
    NANDX1 U10958 (.A1(n15980), .A2(N5225), .ZN(N23830));
    NOR2X1 U10959 (.A1(N12167), .A2(n20065), .ZN(N23831));
    INVX1 U10960 (.I(n16654), .ZN(N23832));
    INVX1 U10961 (.I(N3526), .ZN(n23833));
    NANDX1 U10962 (.A1(n16261), .A2(N1683), .ZN(n23834));
    NOR2X1 U10963 (.A1(N4285), .A2(n18397), .ZN(n23835));
    NANDX1 U10964 (.A1(n20838), .A2(N10842), .ZN(n23836));
    INVX1 U10965 (.I(N11384), .ZN(n23837));
    NANDX1 U10966 (.A1(n18632), .A2(n14322), .ZN(n23838));
    INVX1 U10967 (.I(n18696), .ZN(n23839));
    NOR2X1 U10968 (.A1(n15930), .A2(N10648), .ZN(n23840));
    NANDX1 U10969 (.A1(N6974), .A2(N423), .ZN(n23841));
    NOR2X1 U10970 (.A1(N6740), .A2(n13537), .ZN(n23842));
    NOR2X1 U10971 (.A1(N116), .A2(n13708), .ZN(N23843));
    NOR2X1 U10972 (.A1(n17447), .A2(N11775), .ZN(N23844));
    NANDX1 U10973 (.A1(N7019), .A2(N7999), .ZN(N23845));
    NANDX1 U10974 (.A1(N11303), .A2(N5165), .ZN(N23846));
    INVX1 U10975 (.I(N5453), .ZN(N23847));
    NANDX1 U10976 (.A1(n15023), .A2(n16836), .ZN(N23848));
    NANDX1 U10977 (.A1(N6966), .A2(N4470), .ZN(n23849));
    NANDX1 U10978 (.A1(N4431), .A2(N3660), .ZN(n23850));
    NOR2X1 U10979 (.A1(N9620), .A2(N4870), .ZN(n23851));
    INVX1 U10980 (.I(N4584), .ZN(N23852));
    NOR2X1 U10981 (.A1(N9069), .A2(n18121), .ZN(N23853));
    NANDX1 U10982 (.A1(N9185), .A2(N5140), .ZN(n23854));
    NANDX1 U10983 (.A1(n21173), .A2(n16914), .ZN(n23855));
    INVX1 U10984 (.I(N6961), .ZN(n23856));
    NOR2X1 U10985 (.A1(N11517), .A2(N12805), .ZN(n23857));
    NANDX1 U10986 (.A1(N11605), .A2(n18257), .ZN(N23858));
    NANDX1 U10987 (.A1(n21169), .A2(N8405), .ZN(n23859));
    INVX1 U10988 (.I(N6904), .ZN(n23860));
    NANDX1 U10989 (.A1(N6701), .A2(N5877), .ZN(N23861));
    INVX1 U10990 (.I(N7515), .ZN(n23862));
    NANDX1 U10991 (.A1(n15945), .A2(N9844), .ZN(n23863));
    INVX1 U10992 (.I(n16773), .ZN(n23864));
    NOR2X1 U10993 (.A1(N6054), .A2(n14811), .ZN(n23865));
    NANDX1 U10994 (.A1(N11193), .A2(N10939), .ZN(n23866));
    NOR2X1 U10995 (.A1(N1418), .A2(N262), .ZN(n23867));
    NOR2X1 U10996 (.A1(n20871), .A2(N11778), .ZN(n23868));
    INVX1 U10997 (.I(n18800), .ZN(N23869));
    NOR2X1 U10998 (.A1(N12683), .A2(N11505), .ZN(N23870));
    NOR2X1 U10999 (.A1(n21087), .A2(N6633), .ZN(n23871));
    NANDX1 U11000 (.A1(N7272), .A2(N7876), .ZN(N23872));
    NOR2X1 U11001 (.A1(n18347), .A2(N9932), .ZN(n23873));
    NANDX1 U11002 (.A1(N7603), .A2(n19775), .ZN(N23874));
    NANDX1 U11003 (.A1(N3145), .A2(n17456), .ZN(n23875));
    INVX1 U11004 (.I(N12497), .ZN(n23876));
    NOR2X1 U11005 (.A1(N8254), .A2(N2205), .ZN(n23877));
    NANDX1 U11006 (.A1(N9671), .A2(n18238), .ZN(N23878));
    NOR2X1 U11007 (.A1(N3853), .A2(N3328), .ZN(n23879));
    INVX1 U11008 (.I(N1423), .ZN(n23880));
    INVX1 U11009 (.I(N3485), .ZN(n23881));
    NOR2X1 U11010 (.A1(N12426), .A2(n19114), .ZN(n23882));
    NANDX1 U11011 (.A1(N5046), .A2(N5155), .ZN(n23883));
    NANDX1 U11012 (.A1(N3542), .A2(n18043), .ZN(n23884));
    NOR2X1 U11013 (.A1(N6618), .A2(N4415), .ZN(n23885));
    NOR2X1 U11014 (.A1(n18856), .A2(N2102), .ZN(n23886));
    NOR2X1 U11015 (.A1(n15918), .A2(N9140), .ZN(n23887));
    NANDX1 U11016 (.A1(N2941), .A2(N11345), .ZN(n23888));
    NANDX1 U11017 (.A1(N7154), .A2(N8352), .ZN(N23889));
    INVX1 U11018 (.I(N11006), .ZN(n23890));
    NANDX1 U11019 (.A1(n20183), .A2(N6970), .ZN(N23891));
    NOR2X1 U11020 (.A1(N2437), .A2(n14439), .ZN(n23892));
    INVX1 U11021 (.I(n16092), .ZN(n23893));
    INVX1 U11022 (.I(N2483), .ZN(N23894));
    NOR2X1 U11023 (.A1(n12912), .A2(N567), .ZN(n23895));
    NOR2X1 U11024 (.A1(N12673), .A2(N1726), .ZN(N23896));
    NANDX1 U11025 (.A1(N10978), .A2(n20581), .ZN(N23897));
    NOR2X1 U11026 (.A1(n15822), .A2(N9810), .ZN(n23898));
    NOR2X1 U11027 (.A1(n18300), .A2(N7293), .ZN(n23899));
    NOR2X1 U11028 (.A1(N8844), .A2(n14446), .ZN(n23900));
    INVX1 U11029 (.I(n16994), .ZN(n23901));
    INVX1 U11030 (.I(n16568), .ZN(n23902));
    NANDX1 U11031 (.A1(N5733), .A2(N1580), .ZN(n23903));
    NANDX1 U11032 (.A1(n14713), .A2(n20247), .ZN(n23904));
    NANDX1 U11033 (.A1(n16564), .A2(n17271), .ZN(N23905));
    NANDX1 U11034 (.A1(N8245), .A2(n17837), .ZN(n23906));
    NANDX1 U11035 (.A1(n20917), .A2(n19562), .ZN(n23907));
    INVX1 U11036 (.I(N5206), .ZN(N23908));
    NOR2X1 U11037 (.A1(N2555), .A2(n21027), .ZN(n23909));
    INVX1 U11038 (.I(n14437), .ZN(n23910));
    NANDX1 U11039 (.A1(N9326), .A2(n16432), .ZN(n23911));
    NOR2X1 U11040 (.A1(n18313), .A2(N5549), .ZN(n23912));
    INVX1 U11041 (.I(N11618), .ZN(n23913));
    NOR2X1 U11042 (.A1(n16815), .A2(N11892), .ZN(n23914));
    NOR2X1 U11043 (.A1(N3051), .A2(N5374), .ZN(n23915));
    NANDX1 U11044 (.A1(N5378), .A2(N707), .ZN(n23916));
    INVX1 U11045 (.I(N7721), .ZN(n23917));
    INVX1 U11046 (.I(N4443), .ZN(n23918));
    INVX1 U11047 (.I(N3179), .ZN(n23919));
    NOR2X1 U11048 (.A1(N6103), .A2(N2926), .ZN(n23920));
    NANDX1 U11049 (.A1(N3199), .A2(N2722), .ZN(n23921));
    INVX1 U11050 (.I(n17635), .ZN(N23922));
    INVX1 U11051 (.I(n16671), .ZN(n23923));
    NOR2X1 U11052 (.A1(N4694), .A2(N8296), .ZN(n23924));
    NANDX1 U11053 (.A1(N11022), .A2(n19913), .ZN(N23925));
    NANDX1 U11054 (.A1(N6606), .A2(N10574), .ZN(N23926));
    INVX1 U11055 (.I(N9656), .ZN(n23927));
    NANDX1 U11056 (.A1(n17157), .A2(N9575), .ZN(n23928));
    NOR2X1 U11057 (.A1(N3763), .A2(N11837), .ZN(n23929));
    NOR2X1 U11058 (.A1(N8205), .A2(N2355), .ZN(n23930));
    INVX1 U11059 (.I(N5520), .ZN(n23931));
    NOR2X1 U11060 (.A1(n15332), .A2(N10832), .ZN(n23932));
    INVX1 U11061 (.I(N12595), .ZN(n23933));
    INVX1 U11062 (.I(n18374), .ZN(n23934));
    INVX1 U11063 (.I(N8159), .ZN(n23935));
    NOR2X1 U11064 (.A1(N5960), .A2(N10996), .ZN(n23936));
    NANDX1 U11065 (.A1(N11523), .A2(N9678), .ZN(n23937));
    NANDX1 U11066 (.A1(N12670), .A2(n14793), .ZN(n23938));
    NOR2X1 U11067 (.A1(n16868), .A2(N4051), .ZN(n23939));
    NOR2X1 U11068 (.A1(N5212), .A2(n15245), .ZN(n23940));
    NANDX1 U11069 (.A1(n17049), .A2(N3243), .ZN(n23941));
    NOR2X1 U11070 (.A1(n19403), .A2(n15649), .ZN(N23942));
    INVX1 U11071 (.I(N1171), .ZN(n23943));
    NOR2X1 U11072 (.A1(N1429), .A2(N1909), .ZN(N23944));
    INVX1 U11073 (.I(n19605), .ZN(n23945));
    NANDX1 U11074 (.A1(N12694), .A2(N1076), .ZN(n23946));
    NANDX1 U11075 (.A1(n18653), .A2(N12071), .ZN(N23947));
    INVX1 U11076 (.I(N3487), .ZN(n23948));
    INVX1 U11077 (.I(N3761), .ZN(n23949));
    NANDX1 U11078 (.A1(N4395), .A2(n18550), .ZN(n23950));
    NOR2X1 U11079 (.A1(N8446), .A2(N2578), .ZN(N23951));
    INVX1 U11080 (.I(N2460), .ZN(n23952));
    NANDX1 U11081 (.A1(N12823), .A2(N245), .ZN(n23953));
    INVX1 U11082 (.I(N5537), .ZN(N23954));
    NOR2X1 U11083 (.A1(n19420), .A2(N1249), .ZN(n23955));
    INVX1 U11084 (.I(n20848), .ZN(n23956));
    INVX1 U11085 (.I(N10383), .ZN(n23957));
    INVX1 U11086 (.I(n17981), .ZN(n23958));
    NOR2X1 U11087 (.A1(N9382), .A2(n16096), .ZN(n23959));
    NOR2X1 U11088 (.A1(n15994), .A2(N4970), .ZN(n23960));
    NOR2X1 U11089 (.A1(N5596), .A2(N3272), .ZN(n23961));
    INVX1 U11090 (.I(N9991), .ZN(n23962));
    INVX1 U11091 (.I(n19788), .ZN(N23963));
    INVX1 U11092 (.I(N3169), .ZN(n23964));
    NANDX1 U11093 (.A1(n15437), .A2(N9308), .ZN(n23965));
    NOR2X1 U11094 (.A1(n15681), .A2(N11442), .ZN(n23966));
    NANDX1 U11095 (.A1(N4886), .A2(N9631), .ZN(N23967));
    NOR2X1 U11096 (.A1(n19612), .A2(N3790), .ZN(n23968));
    INVX1 U11097 (.I(N3306), .ZN(n23969));
    INVX1 U11098 (.I(n18704), .ZN(n23970));
    NANDX1 U11099 (.A1(n16019), .A2(N8111), .ZN(n23971));
    NANDX1 U11100 (.A1(N10783), .A2(n13080), .ZN(n23972));
    NANDX1 U11101 (.A1(n16378), .A2(N10893), .ZN(n23973));
    NANDX1 U11102 (.A1(n20910), .A2(N6025), .ZN(n23974));
    NOR2X1 U11103 (.A1(n18115), .A2(N9193), .ZN(N23975));
    INVX1 U11104 (.I(N6864), .ZN(n23976));
    NOR2X1 U11105 (.A1(N3092), .A2(N1314), .ZN(n23977));
    NANDX1 U11106 (.A1(N4867), .A2(N741), .ZN(N23978));
    NOR2X1 U11107 (.A1(N7891), .A2(n14894), .ZN(n23979));
    NOR2X1 U11108 (.A1(N8613), .A2(N12741), .ZN(n23980));
    NANDX1 U11109 (.A1(N628), .A2(N12434), .ZN(N23981));
    NANDX1 U11110 (.A1(N8738), .A2(n16250), .ZN(n23982));
    NANDX1 U11111 (.A1(n16359), .A2(N6447), .ZN(N23983));
    INVX1 U11112 (.I(N6021), .ZN(n23984));
    NOR2X1 U11113 (.A1(N12792), .A2(N12046), .ZN(n23985));
    NOR2X1 U11114 (.A1(N4219), .A2(n15780), .ZN(n23986));
    NOR2X1 U11115 (.A1(N11082), .A2(N7592), .ZN(n23987));
    NOR2X1 U11116 (.A1(N6937), .A2(N10845), .ZN(N23988));
    NANDX1 U11117 (.A1(N7678), .A2(n18270), .ZN(n23989));
    INVX1 U11118 (.I(N1341), .ZN(n23990));
    NANDX1 U11119 (.A1(N6013), .A2(n14082), .ZN(N23991));
    NOR2X1 U11120 (.A1(N6641), .A2(n21057), .ZN(n23992));
    INVX1 U11121 (.I(n15378), .ZN(n23993));
    NOR2X1 U11122 (.A1(n14252), .A2(N10507), .ZN(N23994));
    NANDX1 U11123 (.A1(N676), .A2(N11069), .ZN(n23995));
    INVX1 U11124 (.I(N8009), .ZN(n23996));
    INVX1 U11125 (.I(n17632), .ZN(n23997));
    NANDX1 U11126 (.A1(n17664), .A2(N4642), .ZN(n23998));
    NOR2X1 U11127 (.A1(n19797), .A2(N10515), .ZN(n23999));
    INVX1 U11128 (.I(N9412), .ZN(n24000));
    INVX1 U11129 (.I(N11234), .ZN(n24001));
    INVX1 U11130 (.I(N2883), .ZN(n24002));
    INVX1 U11131 (.I(N9247), .ZN(n24003));
    INVX1 U11132 (.I(n15739), .ZN(n24004));
    NOR2X1 U11133 (.A1(N10078), .A2(N10107), .ZN(n24005));
    NANDX1 U11134 (.A1(n19997), .A2(n15267), .ZN(n24006));
    NANDX1 U11135 (.A1(N3815), .A2(N5643), .ZN(n24007));
    INVX1 U11136 (.I(n14884), .ZN(n24008));
    INVX1 U11137 (.I(n16970), .ZN(n24009));
    NOR2X1 U11138 (.A1(N2516), .A2(N7967), .ZN(N24010));
    NOR2X1 U11139 (.A1(N1699), .A2(N4586), .ZN(n24011));
    INVX1 U11140 (.I(N12213), .ZN(n24012));
    NOR2X1 U11141 (.A1(N10262), .A2(N12238), .ZN(n24013));
    NOR2X1 U11142 (.A1(n16712), .A2(N9662), .ZN(n24014));
    NANDX1 U11143 (.A1(n20501), .A2(n13099), .ZN(n24015));
    NANDX1 U11144 (.A1(N7935), .A2(n17718), .ZN(n24016));
    NANDX1 U11145 (.A1(N7428), .A2(n16485), .ZN(n24017));
    INVX1 U11146 (.I(n15714), .ZN(n24018));
    NOR2X1 U11147 (.A1(n14410), .A2(N3445), .ZN(n24019));
    NANDX1 U11148 (.A1(n15066), .A2(n20415), .ZN(n24020));
    NOR2X1 U11149 (.A1(N12123), .A2(N1693), .ZN(n24021));
    NOR2X1 U11150 (.A1(n13821), .A2(N6278), .ZN(n24022));
    NOR2X1 U11151 (.A1(n20575), .A2(N8962), .ZN(N24023));
    INVX1 U11152 (.I(N11582), .ZN(N24024));
    INVX1 U11153 (.I(N1991), .ZN(n24025));
    NANDX1 U11154 (.A1(N11764), .A2(N1261), .ZN(n24026));
    INVX1 U11155 (.I(n16389), .ZN(N24027));
    INVX1 U11156 (.I(n19914), .ZN(N24028));
    INVX1 U11157 (.I(N11165), .ZN(n24029));
    NANDX1 U11158 (.A1(n18657), .A2(N190), .ZN(n24030));
    INVX1 U11159 (.I(N11836), .ZN(n24031));
    NOR2X1 U11160 (.A1(N6356), .A2(N213), .ZN(n24032));
    NANDX1 U11161 (.A1(N4928), .A2(N12335), .ZN(N24033));
    NOR2X1 U11162 (.A1(N325), .A2(n20697), .ZN(n24034));
    NOR2X1 U11163 (.A1(N2031), .A2(n20041), .ZN(n24035));
    NANDX1 U11164 (.A1(n13997), .A2(N4935), .ZN(n24036));
    INVX1 U11165 (.I(n15987), .ZN(n24037));
    INVX1 U11166 (.I(n16786), .ZN(n24038));
    NOR2X1 U11167 (.A1(N1685), .A2(N11944), .ZN(n24039));
    NANDX1 U11168 (.A1(n16140), .A2(N603), .ZN(n24040));
    NOR2X1 U11169 (.A1(N4619), .A2(n13801), .ZN(N24041));
    INVX1 U11170 (.I(N7939), .ZN(n24042));
    INVX1 U11171 (.I(N9283), .ZN(N24043));
    NOR2X1 U11172 (.A1(n20390), .A2(N1185), .ZN(n24044));
    NOR2X1 U11173 (.A1(N11494), .A2(N237), .ZN(n24045));
    NANDX1 U11174 (.A1(N10960), .A2(N109), .ZN(n24046));
    NANDX1 U11175 (.A1(N4313), .A2(N8941), .ZN(N24047));
    NOR2X1 U11176 (.A1(N3789), .A2(N8505), .ZN(n24048));
    NOR2X1 U11177 (.A1(n19050), .A2(N4061), .ZN(n24049));
    NOR2X1 U11178 (.A1(n20734), .A2(N10546), .ZN(n24050));
    NANDX1 U11179 (.A1(N10186), .A2(N5691), .ZN(n24051));
    INVX1 U11180 (.I(n14804), .ZN(N24052));
    NANDX1 U11181 (.A1(N9915), .A2(n17284), .ZN(N24053));
    NOR2X1 U11182 (.A1(n13740), .A2(N4889), .ZN(n24054));
    NANDX1 U11183 (.A1(n14924), .A2(n13193), .ZN(n24055));
    INVX1 U11184 (.I(n15161), .ZN(n24056));
    INVX1 U11185 (.I(N7905), .ZN(n24057));
    INVX1 U11186 (.I(N5792), .ZN(n24058));
    NOR2X1 U11187 (.A1(n13293), .A2(N3759), .ZN(n24059));
    INVX1 U11188 (.I(N568), .ZN(n24060));
    NANDX1 U11189 (.A1(N8366), .A2(n20400), .ZN(N24061));
    NANDX1 U11190 (.A1(N2412), .A2(N9715), .ZN(N24062));
    NOR2X1 U11191 (.A1(N12597), .A2(N9947), .ZN(n24063));
    INVX1 U11192 (.I(N6170), .ZN(n24064));
    INVX1 U11193 (.I(n19440), .ZN(N24065));
    INVX1 U11194 (.I(n21188), .ZN(N24066));
    INVX1 U11195 (.I(N1654), .ZN(n24067));
    NOR2X1 U11196 (.A1(N5643), .A2(N9389), .ZN(N24068));
    NOR2X1 U11197 (.A1(n15345), .A2(N4522), .ZN(N24069));
    INVX1 U11198 (.I(n19697), .ZN(n24070));
    NANDX1 U11199 (.A1(N2475), .A2(N11759), .ZN(n24071));
    NANDX1 U11200 (.A1(n13022), .A2(N6868), .ZN(n24072));
    NOR2X1 U11201 (.A1(N157), .A2(N6037), .ZN(n24073));
    INVX1 U11202 (.I(n18340), .ZN(n24074));
    NOR2X1 U11203 (.A1(N11349), .A2(N9706), .ZN(n24075));
    INVX1 U11204 (.I(n15416), .ZN(n24076));
    NOR2X1 U11205 (.A1(N1759), .A2(n13625), .ZN(n24077));
    NOR2X1 U11206 (.A1(N1716), .A2(N4344), .ZN(n24078));
    NANDX1 U11207 (.A1(N8355), .A2(N4528), .ZN(N24079));
    NANDX1 U11208 (.A1(n17396), .A2(n14414), .ZN(N24080));
    NOR2X1 U11209 (.A1(n13112), .A2(n12880), .ZN(N24081));
    NOR2X1 U11210 (.A1(n15587), .A2(N3408), .ZN(n24082));
    INVX1 U11211 (.I(N7378), .ZN(n24083));
    NOR2X1 U11212 (.A1(N3704), .A2(N2076), .ZN(N24084));
    NOR2X1 U11213 (.A1(N9793), .A2(n20416), .ZN(n24085));
    NANDX1 U11214 (.A1(n15683), .A2(N3433), .ZN(n24086));
    INVX1 U11215 (.I(N9868), .ZN(n24087));
    INVX1 U11216 (.I(N10999), .ZN(n24088));
    NANDX1 U11217 (.A1(n15574), .A2(N12715), .ZN(n24089));
    NANDX1 U11218 (.A1(n13494), .A2(n15611), .ZN(n24090));
    INVX1 U11219 (.I(n20801), .ZN(n24091));
    INVX1 U11220 (.I(n14629), .ZN(N24092));
    NANDX1 U11221 (.A1(N3658), .A2(N6278), .ZN(n24093));
    NANDX1 U11222 (.A1(n19244), .A2(N9686), .ZN(n24094));
    NANDX1 U11223 (.A1(n21163), .A2(n14503), .ZN(n24095));
    NANDX1 U11224 (.A1(N2008), .A2(n19898), .ZN(n24096));
    NOR2X1 U11225 (.A1(n16965), .A2(n19815), .ZN(N24097));
    NOR2X1 U11226 (.A1(n20398), .A2(N7825), .ZN(N24098));
    INVX1 U11227 (.I(N7559), .ZN(n24099));
    INVX1 U11228 (.I(N9162), .ZN(n24100));
    NANDX1 U11229 (.A1(N4849), .A2(N4851), .ZN(n24101));
    NANDX1 U11230 (.A1(n20459), .A2(N5066), .ZN(n24102));
    NOR2X1 U11231 (.A1(N5547), .A2(n19695), .ZN(n24103));
    NANDX1 U11232 (.A1(N9204), .A2(N4742), .ZN(N24104));
    NOR2X1 U11233 (.A1(N1759), .A2(N8969), .ZN(n24105));
    NANDX1 U11234 (.A1(n17463), .A2(N2241), .ZN(n24106));
    INVX1 U11235 (.I(n19470), .ZN(n24107));
    INVX1 U11236 (.I(N7359), .ZN(n24108));
    NANDX1 U11237 (.A1(n15265), .A2(N9850), .ZN(n24109));
    NOR2X1 U11238 (.A1(n17631), .A2(n16750), .ZN(n24110));
    NOR2X1 U11239 (.A1(n15223), .A2(N4682), .ZN(n24111));
    NANDX1 U11240 (.A1(n14614), .A2(N9532), .ZN(n24112));
    INVX1 U11241 (.I(N8384), .ZN(n24113));
    NANDX1 U11242 (.A1(N5071), .A2(n13930), .ZN(n24114));
    INVX1 U11243 (.I(N9603), .ZN(N24115));
    INVX1 U11244 (.I(N12345), .ZN(n24116));
    INVX1 U11245 (.I(n19433), .ZN(N24117));
    INVX1 U11246 (.I(N5686), .ZN(n24118));
    NANDX1 U11247 (.A1(n18096), .A2(n15320), .ZN(n24119));
    INVX1 U11248 (.I(n13546), .ZN(n24120));
    NOR2X1 U11249 (.A1(n18193), .A2(N2122), .ZN(n24121));
    INVX1 U11250 (.I(N418), .ZN(n24122));
    INVX1 U11251 (.I(N1359), .ZN(n24123));
    INVX1 U11252 (.I(N8286), .ZN(n24124));
    NANDX1 U11253 (.A1(N2515), .A2(N1669), .ZN(n24125));
    INVX1 U11254 (.I(N3535), .ZN(n24126));
    NOR2X1 U11255 (.A1(n19252), .A2(N3147), .ZN(n24127));
    INVX1 U11256 (.I(N5624), .ZN(n24128));
    NOR2X1 U11257 (.A1(n20427), .A2(n17968), .ZN(n24129));
    NOR2X1 U11258 (.A1(n13171), .A2(n18051), .ZN(N24130));
    NANDX1 U11259 (.A1(N7606), .A2(n14916), .ZN(N24131));
    NANDX1 U11260 (.A1(N10594), .A2(N1773), .ZN(n24132));
    NOR2X1 U11261 (.A1(N7556), .A2(N3894), .ZN(N24133));
    INVX1 U11262 (.I(N2515), .ZN(N24134));
    NANDX1 U11263 (.A1(n14866), .A2(N8487), .ZN(n24135));
    INVX1 U11264 (.I(N9990), .ZN(n24136));
    INVX1 U11265 (.I(N6911), .ZN(N24137));
    INVX1 U11266 (.I(N9078), .ZN(N24138));
    INVX1 U11267 (.I(N12665), .ZN(N24139));
    INVX1 U11268 (.I(n14256), .ZN(N24140));
    INVX1 U11269 (.I(n19515), .ZN(n24141));
    INVX1 U11270 (.I(n15026), .ZN(n24142));
    NOR2X1 U11271 (.A1(n21165), .A2(N6388), .ZN(N24143));
    NANDX1 U11272 (.A1(N2082), .A2(n15845), .ZN(N24144));
    INVX1 U11273 (.I(N12675), .ZN(n24145));
    NOR2X1 U11274 (.A1(n15581), .A2(n14772), .ZN(n24146));
    INVX1 U11275 (.I(N7858), .ZN(n24147));
    NANDX1 U11276 (.A1(n18466), .A2(n17266), .ZN(n24148));
    NANDX1 U11277 (.A1(N2478), .A2(N6025), .ZN(n24149));
    INVX1 U11278 (.I(N3930), .ZN(n24150));
    INVX1 U11279 (.I(n19162), .ZN(N24151));
    NANDX1 U11280 (.A1(N12103), .A2(N4697), .ZN(n24152));
    NOR2X1 U11281 (.A1(N3703), .A2(N2982), .ZN(N24153));
    INVX1 U11282 (.I(n18728), .ZN(n24154));
    INVX1 U11283 (.I(N5471), .ZN(n24155));
    INVX1 U11284 (.I(N9404), .ZN(n24156));
    INVX1 U11285 (.I(n14272), .ZN(n24157));
    NOR2X1 U11286 (.A1(n14768), .A2(N10659), .ZN(n24158));
    INVX1 U11287 (.I(N8309), .ZN(n24159));
    INVX1 U11288 (.I(n14067), .ZN(n24160));
    NANDX1 U11289 (.A1(N2716), .A2(N10102), .ZN(N24161));
    INVX1 U11290 (.I(n20965), .ZN(N24162));
    INVX1 U11291 (.I(n13531), .ZN(n24163));
    NOR2X1 U11292 (.A1(N10105), .A2(N6004), .ZN(N24164));
    INVX1 U11293 (.I(n16749), .ZN(n24165));
    NOR2X1 U11294 (.A1(N867), .A2(n20451), .ZN(n24166));
    INVX1 U11295 (.I(N6403), .ZN(n24167));
    NOR2X1 U11296 (.A1(n15935), .A2(N6415), .ZN(N24168));
    INVX1 U11297 (.I(N4109), .ZN(n24169));
    NANDX1 U11298 (.A1(N3959), .A2(n15967), .ZN(n24170));
    NANDX1 U11299 (.A1(n14617), .A2(N945), .ZN(n24171));
    NANDX1 U11300 (.A1(n20097), .A2(N9553), .ZN(N24172));
    INVX1 U11301 (.I(n17354), .ZN(N24173));
    NOR2X1 U11302 (.A1(N12705), .A2(N11630), .ZN(n24174));
    NOR2X1 U11303 (.A1(n20777), .A2(n15293), .ZN(n24175));
    INVX1 U11304 (.I(N5551), .ZN(n24176));
    INVX1 U11305 (.I(N3798), .ZN(n24177));
    NOR2X1 U11306 (.A1(N3109), .A2(N3019), .ZN(N24178));
    NOR2X1 U11307 (.A1(N9512), .A2(n15509), .ZN(n24179));
    INVX1 U11308 (.I(n15926), .ZN(n24180));
    NOR2X1 U11309 (.A1(N6912), .A2(N3204), .ZN(n24181));
    INVX1 U11310 (.I(n17420), .ZN(n24182));
    NANDX1 U11311 (.A1(N2541), .A2(n12907), .ZN(n24183));
    INVX1 U11312 (.I(n17179), .ZN(n24184));
    NANDX1 U11313 (.A1(n19400), .A2(N7844), .ZN(n24185));
    NANDX1 U11314 (.A1(N5416), .A2(n19473), .ZN(n24186));
    NANDX1 U11315 (.A1(N4963), .A2(N8077), .ZN(n24187));
    NANDX1 U11316 (.A1(N5055), .A2(n15777), .ZN(N24188));
    INVX1 U11317 (.I(N10389), .ZN(n24189));
    INVX1 U11318 (.I(N7464), .ZN(n24190));
    INVX1 U11319 (.I(N1708), .ZN(n24191));
    NOR2X1 U11320 (.A1(N61), .A2(N12176), .ZN(N24192));
    NOR2X1 U11321 (.A1(N6973), .A2(N9921), .ZN(n24193));
    NOR2X1 U11322 (.A1(n18934), .A2(N9710), .ZN(n24194));
    INVX1 U11323 (.I(N10610), .ZN(n24195));
    NANDX1 U11324 (.A1(N9120), .A2(N6381), .ZN(N24196));
    INVX1 U11325 (.I(N11505), .ZN(n24197));
    NOR2X1 U11326 (.A1(n17979), .A2(N9747), .ZN(n24198));
    INVX1 U11327 (.I(n17483), .ZN(n24199));
    NOR2X1 U11328 (.A1(N9363), .A2(N1307), .ZN(n24200));
    INVX1 U11329 (.I(n13808), .ZN(n24201));
    NOR2X1 U11330 (.A1(N4566), .A2(N41), .ZN(n24202));
    NOR2X1 U11331 (.A1(N815), .A2(N1782), .ZN(n24203));
    INVX1 U11332 (.I(n12990), .ZN(n24204));
    INVX1 U11333 (.I(N10527), .ZN(n24205));
    NANDX1 U11334 (.A1(n19349), .A2(N8230), .ZN(n24206));
    NANDX1 U11335 (.A1(N11291), .A2(n13382), .ZN(n24207));
    NOR2X1 U11336 (.A1(n14952), .A2(n14304), .ZN(n24208));
    INVX1 U11337 (.I(N5227), .ZN(n24209));
    INVX1 U11338 (.I(N2949), .ZN(n24210));
    NANDX1 U11339 (.A1(N12676), .A2(n20431), .ZN(n24211));
    NOR2X1 U11340 (.A1(N808), .A2(N508), .ZN(n24212));
    NOR2X1 U11341 (.A1(N9157), .A2(N12202), .ZN(n24213));
    NANDX1 U11342 (.A1(N9197), .A2(n21154), .ZN(N24214));
    NANDX1 U11343 (.A1(N5520), .A2(N3478), .ZN(n24215));
    NOR2X1 U11344 (.A1(N8779), .A2(n14004), .ZN(n24216));
    NOR2X1 U11345 (.A1(N1440), .A2(n16775), .ZN(n24217));
    INVX1 U11346 (.I(N12730), .ZN(n24218));
    NANDX1 U11347 (.A1(N488), .A2(N6451), .ZN(n24219));
    NOR2X1 U11348 (.A1(N6688), .A2(N6219), .ZN(n24220));
    INVX1 U11349 (.I(N9636), .ZN(N24221));
    NOR2X1 U11350 (.A1(n13178), .A2(N8836), .ZN(N24222));
    NANDX1 U11351 (.A1(N8527), .A2(N9343), .ZN(n24223));
    NANDX1 U11352 (.A1(n17684), .A2(n16087), .ZN(n24224));
    NANDX1 U11353 (.A1(N192), .A2(N10552), .ZN(n24225));
    NOR2X1 U11354 (.A1(N5712), .A2(n14029), .ZN(n24226));
    NOR2X1 U11355 (.A1(N9032), .A2(N6802), .ZN(n24227));
    NANDX1 U11356 (.A1(N10471), .A2(n18118), .ZN(n24228));
    NOR2X1 U11357 (.A1(n17742), .A2(N356), .ZN(n24229));
    NANDX1 U11358 (.A1(n18735), .A2(N12668), .ZN(N24230));
    INVX1 U11359 (.I(N3723), .ZN(n24231));
    INVX1 U11360 (.I(n18849), .ZN(n24232));
    NANDX1 U11361 (.A1(n20889), .A2(N6454), .ZN(n24233));
    INVX1 U11362 (.I(N2727), .ZN(N24234));
    NOR2X1 U11363 (.A1(N1548), .A2(n20410), .ZN(n24235));
    INVX1 U11364 (.I(n16384), .ZN(n24236));
    NANDX1 U11365 (.A1(n15746), .A2(n17471), .ZN(n24237));
    INVX1 U11366 (.I(N3086), .ZN(N24238));
    NANDX1 U11367 (.A1(N3198), .A2(N4429), .ZN(n24239));
    NANDX1 U11368 (.A1(N8211), .A2(N1316), .ZN(n24240));
    NANDX1 U11369 (.A1(n20494), .A2(N1671), .ZN(N24241));
    NOR2X1 U11370 (.A1(n17998), .A2(N8881), .ZN(n24242));
    NOR2X1 U11371 (.A1(N491), .A2(N820), .ZN(n24243));
    NOR2X1 U11372 (.A1(n14488), .A2(N478), .ZN(N24244));
    NANDX1 U11373 (.A1(N7866), .A2(N3204), .ZN(n24245));
    INVX1 U11374 (.I(N9413), .ZN(N24246));
    NOR2X1 U11375 (.A1(n19679), .A2(n20338), .ZN(n24247));
    NANDX1 U11376 (.A1(N8736), .A2(N11120), .ZN(n24248));
    NANDX1 U11377 (.A1(N11821), .A2(n18001), .ZN(N24249));
    INVX1 U11378 (.I(n16249), .ZN(n24250));
    NOR2X1 U11379 (.A1(N1268), .A2(N12106), .ZN(n24251));
    NANDX1 U11380 (.A1(N532), .A2(N8319), .ZN(n24252));
    INVX1 U11381 (.I(n18529), .ZN(n24253));
    NOR2X1 U11382 (.A1(N546), .A2(n13561), .ZN(N24254));
    INVX1 U11383 (.I(N3696), .ZN(n24255));
    NOR2X1 U11384 (.A1(N7579), .A2(n13300), .ZN(n24256));
    INVX1 U11385 (.I(N5324), .ZN(n24257));
    NOR2X1 U11386 (.A1(n18638), .A2(N2249), .ZN(n24258));
    INVX1 U11387 (.I(N12287), .ZN(N24259));
    NANDX1 U11388 (.A1(N8279), .A2(N2176), .ZN(n24260));
    INVX1 U11389 (.I(n14641), .ZN(n24261));
    NOR2X1 U11390 (.A1(N2693), .A2(N4201), .ZN(n24262));
    NOR2X1 U11391 (.A1(N3960), .A2(n16307), .ZN(n24263));
    INVX1 U11392 (.I(n20263), .ZN(n24264));
    NANDX1 U11393 (.A1(N1805), .A2(n17562), .ZN(n24265));
    NANDX1 U11394 (.A1(n18122), .A2(N4434), .ZN(N24266));
    NANDX1 U11395 (.A1(N588), .A2(N11252), .ZN(n24267));
    NOR2X1 U11396 (.A1(N8429), .A2(n20477), .ZN(n24268));
    INVX1 U11397 (.I(n14983), .ZN(n24269));
    INVX1 U11398 (.I(n16156), .ZN(n24270));
    NOR2X1 U11399 (.A1(N3482), .A2(n19556), .ZN(n24271));
    NOR2X1 U11400 (.A1(N199), .A2(N2503), .ZN(n24272));
    NANDX1 U11401 (.A1(n14917), .A2(n20967), .ZN(N24273));
    NOR2X1 U11402 (.A1(n18160), .A2(n19468), .ZN(N24274));
    NANDX1 U11403 (.A1(N9180), .A2(n18501), .ZN(n24275));
    INVX1 U11404 (.I(N5526), .ZN(n24276));
    NOR2X1 U11405 (.A1(n17646), .A2(n18190), .ZN(N24277));
    INVX1 U11406 (.I(N2879), .ZN(n24278));
    NOR2X1 U11407 (.A1(n19601), .A2(N11462), .ZN(N24279));
    INVX1 U11408 (.I(n13389), .ZN(n24280));
    INVX1 U11409 (.I(N10041), .ZN(n24281));
    INVX1 U11410 (.I(n20293), .ZN(n24282));
    INVX1 U11411 (.I(n18380), .ZN(N24283));
    NOR2X1 U11412 (.A1(n15225), .A2(n18579), .ZN(n24284));
    NOR2X1 U11413 (.A1(N4751), .A2(N12265), .ZN(n24285));
    NANDX1 U11414 (.A1(n19708), .A2(N3736), .ZN(N24286));
    INVX1 U11415 (.I(N3053), .ZN(n24287));
    NANDX1 U11416 (.A1(n21220), .A2(N5564), .ZN(n24288));
    NANDX1 U11417 (.A1(N9363), .A2(N1979), .ZN(n24289));
    INVX1 U11418 (.I(n17712), .ZN(N24290));
    NANDX1 U11419 (.A1(n17801), .A2(n16082), .ZN(n24291));
    NOR2X1 U11420 (.A1(N12860), .A2(N2782), .ZN(n24292));
    NANDX1 U11421 (.A1(N1670), .A2(N1908), .ZN(n24293));
    NANDX1 U11422 (.A1(n20778), .A2(n20288), .ZN(n24294));
    NANDX1 U11423 (.A1(N9314), .A2(n17636), .ZN(N24295));
    NANDX1 U11424 (.A1(n14065), .A2(N3212), .ZN(n24296));
    NOR2X1 U11425 (.A1(N7084), .A2(N1489), .ZN(N24297));
    NANDX1 U11426 (.A1(N10137), .A2(N3487), .ZN(N24298));
    NOR2X1 U11427 (.A1(n15700), .A2(N11010), .ZN(N24299));
    INVX1 U11428 (.I(N12221), .ZN(n24300));
    NOR2X1 U11429 (.A1(N2541), .A2(N11619), .ZN(n24301));
    NANDX1 U11430 (.A1(n13164), .A2(N1249), .ZN(N24302));
    INVX1 U11431 (.I(n15945), .ZN(n24303));
    NOR2X1 U11432 (.A1(n15676), .A2(N12395), .ZN(n24304));
    NANDX1 U11433 (.A1(N9765), .A2(N11452), .ZN(N24305));
    INVX1 U11434 (.I(n19079), .ZN(n24306));
    INVX1 U11435 (.I(n20342), .ZN(n24307));
    NOR2X1 U11436 (.A1(N152), .A2(n19788), .ZN(n24308));
    INVX1 U11437 (.I(n17412), .ZN(N24309));
    NOR2X1 U11438 (.A1(n18216), .A2(n20898), .ZN(n24310));
    NANDX1 U11439 (.A1(N7228), .A2(N10677), .ZN(n24311));
    NANDX1 U11440 (.A1(n19448), .A2(n20711), .ZN(N24312));
    NOR2X1 U11441 (.A1(N4378), .A2(N628), .ZN(n24313));
    NANDX1 U11442 (.A1(N5626), .A2(n14633), .ZN(N24314));
    NANDX1 U11443 (.A1(n16413), .A2(N3620), .ZN(N24315));
    INVX1 U11444 (.I(n20030), .ZN(n24316));
    INVX1 U11445 (.I(N11053), .ZN(n24317));
    NANDX1 U11446 (.A1(N317), .A2(n13451), .ZN(n24318));
    INVX1 U11447 (.I(N6771), .ZN(n24319));
    INVX1 U11448 (.I(N616), .ZN(n24320));
    NANDX1 U11449 (.A1(N4325), .A2(N1338), .ZN(n24321));
    NANDX1 U11450 (.A1(N3992), .A2(n19987), .ZN(n24322));
    INVX1 U11451 (.I(N9210), .ZN(n24323));
    INVX1 U11452 (.I(N6364), .ZN(n24324));
    NANDX1 U11453 (.A1(n13710), .A2(N10741), .ZN(N24325));
    NANDX1 U11454 (.A1(n17118), .A2(N10909), .ZN(n24326));
    NOR2X1 U11455 (.A1(N4325), .A2(N6091), .ZN(N24327));
    INVX1 U11456 (.I(N9384), .ZN(n24328));
    INVX1 U11457 (.I(n19122), .ZN(n24329));
    NOR2X1 U11458 (.A1(N2379), .A2(n19438), .ZN(n24330));
    NANDX1 U11459 (.A1(N4438), .A2(n20750), .ZN(n24331));
    NANDX1 U11460 (.A1(n20825), .A2(n14369), .ZN(n24332));
    INVX1 U11461 (.I(n16705), .ZN(n24333));
    NANDX1 U11462 (.A1(n18198), .A2(n15461), .ZN(n24334));
    NOR2X1 U11463 (.A1(N6178), .A2(n17694), .ZN(n24335));
    NOR2X1 U11464 (.A1(N9410), .A2(N10173), .ZN(n24336));
    INVX1 U11465 (.I(N7811), .ZN(n24337));
    NANDX1 U11466 (.A1(N3528), .A2(n15386), .ZN(n24338));
    NOR2X1 U11467 (.A1(N4160), .A2(N5351), .ZN(n24339));
    NOR2X1 U11468 (.A1(N3592), .A2(n19014), .ZN(n24340));
    NOR2X1 U11469 (.A1(N5970), .A2(N11763), .ZN(n24341));
    NOR2X1 U11470 (.A1(N10407), .A2(N11282), .ZN(N24342));
    INVX1 U11471 (.I(N4544), .ZN(n24343));
    NANDX1 U11472 (.A1(N12657), .A2(N18), .ZN(n24344));
    INVX1 U11473 (.I(N4166), .ZN(n24345));
    NOR2X1 U11474 (.A1(N682), .A2(N10343), .ZN(n24346));
    NANDX1 U11475 (.A1(N9248), .A2(n14294), .ZN(N24347));
    INVX1 U11476 (.I(N1867), .ZN(n24348));
    NANDX1 U11477 (.A1(N11800), .A2(n21166), .ZN(n24349));
    INVX1 U11478 (.I(N11268), .ZN(n24350));
    NANDX1 U11479 (.A1(N10694), .A2(n14662), .ZN(n24351));
    NANDX1 U11480 (.A1(N8478), .A2(n17262), .ZN(N24352));
    NOR2X1 U11481 (.A1(n14782), .A2(n16143), .ZN(n24353));
    NOR2X1 U11482 (.A1(N4834), .A2(n14592), .ZN(n24354));
    INVX1 U11483 (.I(N3796), .ZN(n24355));
    NANDX1 U11484 (.A1(N12249), .A2(N2273), .ZN(n24356));
    NANDX1 U11485 (.A1(n16810), .A2(n18726), .ZN(n24357));
    NANDX1 U11486 (.A1(n17834), .A2(N6744), .ZN(n24358));
    NANDX1 U11487 (.A1(N7801), .A2(N3152), .ZN(n24359));
    INVX1 U11488 (.I(n14142), .ZN(N24360));
    NANDX1 U11489 (.A1(n13746), .A2(N4180), .ZN(n24361));
    INVX1 U11490 (.I(N3210), .ZN(N24362));
    NOR2X1 U11491 (.A1(n19725), .A2(N6229), .ZN(n24363));
    NANDX1 U11492 (.A1(N6692), .A2(n21010), .ZN(n24364));
    NOR2X1 U11493 (.A1(n19838), .A2(n20385), .ZN(n24365));
    NOR2X1 U11494 (.A1(N10839), .A2(N2950), .ZN(n24366));
    NANDX1 U11495 (.A1(n17629), .A2(n20995), .ZN(n24367));
    NOR2X1 U11496 (.A1(n13208), .A2(n18490), .ZN(n24368));
    NANDX1 U11497 (.A1(N9812), .A2(n19775), .ZN(n24369));
    INVX1 U11498 (.I(N12154), .ZN(n24370));
    NOR2X1 U11499 (.A1(N12139), .A2(N5066), .ZN(n24371));
    NANDX1 U11500 (.A1(N4655), .A2(N9245), .ZN(N24372));
    NANDX1 U11501 (.A1(N2406), .A2(N1397), .ZN(n24373));
    INVX1 U11502 (.I(N8634), .ZN(N24374));
    INVX1 U11503 (.I(N5633), .ZN(n24375));
    NOR2X1 U11504 (.A1(N9678), .A2(N4241), .ZN(n24376));
    NOR2X1 U11505 (.A1(n17679), .A2(N9621), .ZN(n24377));
    INVX1 U11506 (.I(N5010), .ZN(n24378));
    NOR2X1 U11507 (.A1(n20595), .A2(N7379), .ZN(n24379));
    NOR2X1 U11508 (.A1(n17855), .A2(n19358), .ZN(N24380));
    NANDX1 U11509 (.A1(n16399), .A2(N1864), .ZN(N24381));
    NANDX1 U11510 (.A1(N12637), .A2(N8545), .ZN(n24382));
    INVX1 U11511 (.I(N6504), .ZN(n24383));
    INVX1 U11512 (.I(N2125), .ZN(n24384));
    INVX1 U11513 (.I(n15604), .ZN(n24385));
    NANDX1 U11514 (.A1(n16808), .A2(n18779), .ZN(n24386));
    NANDX1 U11515 (.A1(N1211), .A2(n16275), .ZN(n24387));
    NOR2X1 U11516 (.A1(n21223), .A2(n12926), .ZN(n24388));
    NANDX1 U11517 (.A1(N4155), .A2(N12527), .ZN(n24389));
    INVX1 U11518 (.I(N10174), .ZN(n24390));
    NOR2X1 U11519 (.A1(n16471), .A2(N2713), .ZN(n24391));
    NANDX1 U11520 (.A1(n14598), .A2(N5062), .ZN(n24392));
    NOR2X1 U11521 (.A1(N11004), .A2(n19565), .ZN(N24393));
    INVX1 U11522 (.I(n19548), .ZN(n24394));
    INVX1 U11523 (.I(N11908), .ZN(n24395));
    NANDX1 U11524 (.A1(n14569), .A2(n18858), .ZN(n24396));
    INVX1 U11525 (.I(n18090), .ZN(n24397));
    NOR2X1 U11526 (.A1(N8293), .A2(N274), .ZN(n24398));
    NOR2X1 U11527 (.A1(N3337), .A2(N7908), .ZN(N24399));
    INVX1 U11528 (.I(N10805), .ZN(n24400));
    INVX1 U11529 (.I(N8876), .ZN(n24401));
    NOR2X1 U11530 (.A1(n21082), .A2(n13592), .ZN(n24402));
    NANDX1 U11531 (.A1(N10864), .A2(n16304), .ZN(N24403));
    INVX1 U11532 (.I(n20004), .ZN(N24404));
    INVX1 U11533 (.I(N9815), .ZN(n24405));
    INVX1 U11534 (.I(n14242), .ZN(n24406));
    INVX1 U11535 (.I(n18408), .ZN(N24407));
    INVX1 U11536 (.I(N437), .ZN(n24408));
    NOR2X1 U11537 (.A1(n20025), .A2(n19295), .ZN(n24409));
    INVX1 U11538 (.I(N11426), .ZN(n24410));
    INVX1 U11539 (.I(N1041), .ZN(n24411));
    INVX1 U11540 (.I(N6313), .ZN(n24412));
    INVX1 U11541 (.I(n14149), .ZN(n24413));
    INVX1 U11542 (.I(N9723), .ZN(n24414));
    NOR2X1 U11543 (.A1(n14451), .A2(N6365), .ZN(n24415));
    INVX1 U11544 (.I(N1354), .ZN(n24416));
    NOR2X1 U11545 (.A1(N4708), .A2(n17657), .ZN(n24417));
    INVX1 U11546 (.I(N3481), .ZN(n24418));
    INVX1 U11547 (.I(n20529), .ZN(n24419));
    NANDX1 U11548 (.A1(n21117), .A2(N9058), .ZN(N24420));
    NOR2X1 U11549 (.A1(N5342), .A2(N9495), .ZN(n24421));
    NOR2X1 U11550 (.A1(N4136), .A2(N2101), .ZN(n24422));
    NOR2X1 U11551 (.A1(N10103), .A2(N3684), .ZN(n24423));
    NOR2X1 U11552 (.A1(n16344), .A2(N9996), .ZN(n24424));
    INVX1 U11553 (.I(N3804), .ZN(n24425));
    INVX1 U11554 (.I(N10037), .ZN(N24426));
    NOR2X1 U11555 (.A1(N3333), .A2(N10943), .ZN(n24427));
    NOR2X1 U11556 (.A1(N4687), .A2(N4610), .ZN(n24428));
    INVX1 U11557 (.I(n16885), .ZN(n24429));
    INVX1 U11558 (.I(n21056), .ZN(n24430));
    NANDX1 U11559 (.A1(N9164), .A2(N2166), .ZN(n24431));
    NANDX1 U11560 (.A1(N12764), .A2(N1683), .ZN(n24432));
    NOR2X1 U11561 (.A1(N1028), .A2(N4434), .ZN(n24433));
    INVX1 U11562 (.I(n18900), .ZN(n24434));
    INVX1 U11563 (.I(n16538), .ZN(n24435));
    NANDX1 U11564 (.A1(N1328), .A2(N11651), .ZN(N24436));
    NANDX1 U11565 (.A1(N1642), .A2(n15454), .ZN(n24437));
    NANDX1 U11566 (.A1(N6220), .A2(n18707), .ZN(n24438));
    NANDX1 U11567 (.A1(n17162), .A2(N10345), .ZN(n24439));
    INVX1 U11568 (.I(N542), .ZN(N24440));
    NOR2X1 U11569 (.A1(n19675), .A2(n15865), .ZN(n24441));
    NOR2X1 U11570 (.A1(n16746), .A2(n19571), .ZN(n24442));
    NANDX1 U11571 (.A1(n19162), .A2(N11104), .ZN(N24443));
    NOR2X1 U11572 (.A1(N5689), .A2(N6673), .ZN(n24444));
    NANDX1 U11573 (.A1(N12123), .A2(N4342), .ZN(N24445));
    NOR2X1 U11574 (.A1(N1972), .A2(N236), .ZN(N24446));
    INVX1 U11575 (.I(n13622), .ZN(n24447));
    NANDX1 U11576 (.A1(n17097), .A2(N2387), .ZN(n24448));
    INVX1 U11577 (.I(N2086), .ZN(n24449));
    INVX1 U11578 (.I(n20229), .ZN(n24450));
    NANDX1 U11579 (.A1(N4750), .A2(n17561), .ZN(n24451));
    NANDX1 U11580 (.A1(n16898), .A2(n16005), .ZN(n24452));
    INVX1 U11581 (.I(n17955), .ZN(n24453));
    INVX1 U11582 (.I(N1847), .ZN(N24454));
    INVX1 U11583 (.I(N3993), .ZN(n24455));
    NOR2X1 U11584 (.A1(N10312), .A2(N4223), .ZN(n24456));
    NOR2X1 U11585 (.A1(n19651), .A2(N10888), .ZN(N24457));
    NANDX1 U11586 (.A1(n18006), .A2(N12859), .ZN(n24458));
    NANDX1 U11587 (.A1(N12231), .A2(N5251), .ZN(n24459));
    INVX1 U11588 (.I(N8097), .ZN(n24460));
    NANDX1 U11589 (.A1(N9385), .A2(N10182), .ZN(n24461));
    INVX1 U11590 (.I(N8383), .ZN(n24462));
    NANDX1 U11591 (.A1(N1333), .A2(N4713), .ZN(n24463));
    INVX1 U11592 (.I(n18230), .ZN(n24464));
    NANDX1 U11593 (.A1(N4804), .A2(n14954), .ZN(n24465));
    NOR2X1 U11594 (.A1(N1192), .A2(n14902), .ZN(N24466));
    NOR2X1 U11595 (.A1(N8683), .A2(N3983), .ZN(n24467));
    NANDX1 U11596 (.A1(N1616), .A2(n18175), .ZN(N24468));
    NOR2X1 U11597 (.A1(n14662), .A2(n14950), .ZN(n24469));
    INVX1 U11598 (.I(N1255), .ZN(n24470));
    INVX1 U11599 (.I(N5155), .ZN(n24471));
    NANDX1 U11600 (.A1(N8589), .A2(N7334), .ZN(N24472));
    NOR2X1 U11601 (.A1(n13313), .A2(N3917), .ZN(n24473));
    NANDX1 U11602 (.A1(n16053), .A2(N5249), .ZN(n24474));
    INVX1 U11603 (.I(N11892), .ZN(n24475));
    NANDX1 U11604 (.A1(n15336), .A2(N11238), .ZN(n24476));
    INVX1 U11605 (.I(n15426), .ZN(n24477));
    NANDX1 U11606 (.A1(n15728), .A2(N8592), .ZN(n24478));
    NANDX1 U11607 (.A1(n19710), .A2(N11439), .ZN(n24479));
    INVX1 U11608 (.I(N11196), .ZN(n24480));
    INVX1 U11609 (.I(N10701), .ZN(n24481));
    NOR2X1 U11610 (.A1(N3848), .A2(N11955), .ZN(n24482));
    NOR2X1 U11611 (.A1(N3544), .A2(N469), .ZN(N24483));
    NOR2X1 U11612 (.A1(N10877), .A2(N3824), .ZN(n24484));
    NANDX1 U11613 (.A1(N9335), .A2(N4646), .ZN(n24485));
    NANDX1 U11614 (.A1(N9125), .A2(N10181), .ZN(N24486));
    INVX1 U11615 (.I(N5914), .ZN(n24487));
    INVX1 U11616 (.I(N7655), .ZN(n24488));
    INVX1 U11617 (.I(n14253), .ZN(N24489));
    INVX1 U11618 (.I(N1238), .ZN(n24490));
    NOR2X1 U11619 (.A1(n14506), .A2(n15490), .ZN(n24491));
    NANDX1 U11620 (.A1(N10545), .A2(N5455), .ZN(n24492));
    NANDX1 U11621 (.A1(n15787), .A2(N4912), .ZN(N24493));
    INVX1 U11622 (.I(N6511), .ZN(n24494));
    NOR2X1 U11623 (.A1(N8012), .A2(N6979), .ZN(n24495));
    NOR2X1 U11624 (.A1(n13430), .A2(N5345), .ZN(n24496));
    INVX1 U11625 (.I(n17307), .ZN(n24497));
    NANDX1 U11626 (.A1(N3400), .A2(N5201), .ZN(n24498));
    NOR2X1 U11627 (.A1(n21047), .A2(N5657), .ZN(n24499));
    NOR2X1 U11628 (.A1(N7471), .A2(N12397), .ZN(n24500));
    INVX1 U11629 (.I(N865), .ZN(n24501));
    NANDX1 U11630 (.A1(N2717), .A2(n15371), .ZN(n24502));
    INVX1 U11631 (.I(N10311), .ZN(n24503));
    NANDX1 U11632 (.A1(N2432), .A2(n16389), .ZN(n24504));
    NOR2X1 U11633 (.A1(N1885), .A2(n15399), .ZN(n24505));
    NOR2X1 U11634 (.A1(N1288), .A2(N2180), .ZN(N24506));
    INVX1 U11635 (.I(N3770), .ZN(n24507));
    NANDX1 U11636 (.A1(N1700), .A2(N1413), .ZN(n24508));
    INVX1 U11637 (.I(N11689), .ZN(n24509));
    NANDX1 U11638 (.A1(N11428), .A2(N5171), .ZN(n24510));
    NOR2X1 U11639 (.A1(N11626), .A2(n18709), .ZN(n24511));
    NANDX1 U11640 (.A1(n18564), .A2(N4040), .ZN(N24512));
    NOR2X1 U11641 (.A1(N5509), .A2(N6756), .ZN(n24513));
    INVX1 U11642 (.I(N2486), .ZN(n24514));
    INVX1 U11643 (.I(N11185), .ZN(N24515));
    NOR2X1 U11644 (.A1(N1308), .A2(N4967), .ZN(N24516));
    NANDX1 U11645 (.A1(n16706), .A2(n21031), .ZN(n24517));
    INVX1 U11646 (.I(n18885), .ZN(n24518));
    NANDX1 U11647 (.A1(N6399), .A2(N7806), .ZN(N24519));
    NANDX1 U11648 (.A1(N2354), .A2(n14032), .ZN(n24520));
    NANDX1 U11649 (.A1(N1707), .A2(n20001), .ZN(n24521));
    NOR2X1 U11650 (.A1(N877), .A2(N10396), .ZN(n24522));
    NANDX1 U11651 (.A1(N7516), .A2(N7729), .ZN(n24523));
    NANDX1 U11652 (.A1(N9562), .A2(N7780), .ZN(n24524));
    NOR2X1 U11653 (.A1(N290), .A2(N10265), .ZN(n24525));
    NOR2X1 U11654 (.A1(N11474), .A2(N9723), .ZN(n24526));
    NANDX1 U11655 (.A1(N10982), .A2(n16523), .ZN(N24527));
    NANDX1 U11656 (.A1(N10783), .A2(n19153), .ZN(n24528));
    NANDX1 U11657 (.A1(N1480), .A2(n20093), .ZN(n24529));
    NOR2X1 U11658 (.A1(n20565), .A2(N1216), .ZN(N24530));
    INVX1 U11659 (.I(N3420), .ZN(N24531));
    NOR2X1 U11660 (.A1(N11432), .A2(N7217), .ZN(n24532));
    NANDX1 U11661 (.A1(n16369), .A2(N8492), .ZN(n24533));
    INVX1 U11662 (.I(n18640), .ZN(N24534));
    NOR2X1 U11663 (.A1(N9960), .A2(N5189), .ZN(N24535));
    NANDX1 U11664 (.A1(N10249), .A2(N9995), .ZN(n24536));
    NANDX1 U11665 (.A1(n16265), .A2(n19717), .ZN(n24537));
    NOR2X1 U11666 (.A1(N6016), .A2(N9551), .ZN(n24538));
    NANDX1 U11667 (.A1(N11340), .A2(N2015), .ZN(N24539));
    NOR2X1 U11668 (.A1(N12820), .A2(N878), .ZN(n24540));
    NOR2X1 U11669 (.A1(N6696), .A2(n17865), .ZN(n24541));
    INVX1 U11670 (.I(N4657), .ZN(n24542));
    NANDX1 U11671 (.A1(n16959), .A2(N11873), .ZN(n24543));
    NOR2X1 U11672 (.A1(N6639), .A2(n14906), .ZN(N24544));
    NANDX1 U11673 (.A1(N4048), .A2(n17796), .ZN(n24545));
    NOR2X1 U11674 (.A1(N3778), .A2(N610), .ZN(n24546));
    NANDX1 U11675 (.A1(N8314), .A2(N11956), .ZN(n24547));
    NANDX1 U11676 (.A1(N6800), .A2(n16140), .ZN(n24548));
    NOR2X1 U11677 (.A1(N10893), .A2(N8637), .ZN(n24549));
    INVX1 U11678 (.I(N7449), .ZN(n24550));
    NOR2X1 U11679 (.A1(n16420), .A2(N2868), .ZN(n24551));
    NANDX1 U11680 (.A1(N1885), .A2(n20733), .ZN(N24552));
    NANDX1 U11681 (.A1(N6541), .A2(N9373), .ZN(n24553));
    NANDX1 U11682 (.A1(n12955), .A2(N1812), .ZN(n24554));
    NANDX1 U11683 (.A1(N1173), .A2(N10420), .ZN(N24555));
    NANDX1 U11684 (.A1(n13510), .A2(N7757), .ZN(n24556));
    NANDX1 U11685 (.A1(N8661), .A2(n15342), .ZN(N24557));
    NOR2X1 U11686 (.A1(n20616), .A2(N12504), .ZN(n24558));
    NANDX1 U11687 (.A1(n15525), .A2(N10223), .ZN(n24559));
    INVX1 U11688 (.I(n18704), .ZN(n24560));
    NANDX1 U11689 (.A1(N12165), .A2(n16120), .ZN(n24561));
    NOR2X1 U11690 (.A1(n15033), .A2(N944), .ZN(n24562));
    INVX1 U11691 (.I(N9077), .ZN(n24563));
    NANDX1 U11692 (.A1(N11980), .A2(n18449), .ZN(n24564));
    INVX1 U11693 (.I(n19476), .ZN(n24565));
    NOR2X1 U11694 (.A1(N7095), .A2(n15190), .ZN(n24566));
    INVX1 U11695 (.I(n14175), .ZN(n24567));
    NOR2X1 U11696 (.A1(N11747), .A2(n19574), .ZN(n24568));
    NANDX1 U11697 (.A1(N401), .A2(n17514), .ZN(n24569));
    INVX1 U11698 (.I(N7446), .ZN(n24570));
    INVX1 U11699 (.I(n20124), .ZN(n24571));
    NOR2X1 U11700 (.A1(N10596), .A2(n17597), .ZN(n24572));
    NANDX1 U11701 (.A1(N1531), .A2(N7028), .ZN(n24573));
    NANDX1 U11702 (.A1(N11105), .A2(N7972), .ZN(N24574));
    INVX1 U11703 (.I(n20181), .ZN(n24575));
    INVX1 U11704 (.I(n15460), .ZN(n24576));
    NANDX1 U11705 (.A1(n19101), .A2(n13705), .ZN(n24577));
    NANDX1 U11706 (.A1(N4966), .A2(N7665), .ZN(N24578));
    NOR2X1 U11707 (.A1(n13682), .A2(N9676), .ZN(n24579));
    NANDX1 U11708 (.A1(N12025), .A2(n20347), .ZN(n24580));
    NANDX1 U11709 (.A1(N2850), .A2(N3716), .ZN(n24581));
    NOR2X1 U11710 (.A1(n14188), .A2(N2610), .ZN(N24582));
    NOR2X1 U11711 (.A1(N3553), .A2(n14748), .ZN(n24583));
    NANDX1 U11712 (.A1(n20855), .A2(n16318), .ZN(N24584));
    INVX1 U11713 (.I(N10729), .ZN(n24585));
    NANDX1 U11714 (.A1(n20939), .A2(N9679), .ZN(n24586));
    NOR2X1 U11715 (.A1(N9710), .A2(N390), .ZN(n24587));
    NOR2X1 U11716 (.A1(n17956), .A2(N5902), .ZN(n24588));
    NOR2X1 U11717 (.A1(n20162), .A2(n15404), .ZN(n24589));
    NOR2X1 U11718 (.A1(N8607), .A2(N9965), .ZN(N24590));
    NOR2X1 U11719 (.A1(N2266), .A2(N4926), .ZN(n24591));
    NANDX1 U11720 (.A1(N5981), .A2(N7332), .ZN(N24592));
    NANDX1 U11721 (.A1(N3132), .A2(n16489), .ZN(N24593));
    NOR2X1 U11722 (.A1(n17880), .A2(n14676), .ZN(n24594));
    INVX1 U11723 (.I(n12967), .ZN(n24595));
    INVX1 U11724 (.I(n13287), .ZN(n24596));
    INVX1 U11725 (.I(N5154), .ZN(n24597));
    NOR2X1 U11726 (.A1(N7433), .A2(N9405), .ZN(N24598));
    INVX1 U11727 (.I(n17941), .ZN(N24599));
    NANDX1 U11728 (.A1(n18340), .A2(N6727), .ZN(n24600));
    INVX1 U11729 (.I(N12513), .ZN(n24601));
    INVX1 U11730 (.I(N8210), .ZN(n24602));
    INVX1 U11731 (.I(N2454), .ZN(N24603));
    INVX1 U11732 (.I(N715), .ZN(n24604));
    NANDX1 U11733 (.A1(n16456), .A2(N2589), .ZN(n24605));
    INVX1 U11734 (.I(n19587), .ZN(n24606));
    INVX1 U11735 (.I(N878), .ZN(N24607));
    INVX1 U11736 (.I(N12522), .ZN(n24608));
    NOR2X1 U11737 (.A1(n18286), .A2(n17967), .ZN(N24609));
    INVX1 U11738 (.I(N7622), .ZN(n24610));
    INVX1 U11739 (.I(N7542), .ZN(n24611));
    NOR2X1 U11740 (.A1(N5836), .A2(n19980), .ZN(n24612));
    INVX1 U11741 (.I(N6508), .ZN(N24613));
    NANDX1 U11742 (.A1(N7575), .A2(N11569), .ZN(n24614));
    NOR2X1 U11743 (.A1(N11309), .A2(n19778), .ZN(N24615));
    NOR2X1 U11744 (.A1(n13762), .A2(N9023), .ZN(n24616));
    NOR2X1 U11745 (.A1(N6867), .A2(n20020), .ZN(n24617));
    NOR2X1 U11746 (.A1(N4811), .A2(n18376), .ZN(n24618));
    NOR2X1 U11747 (.A1(N5689), .A2(N7924), .ZN(N24619));
    NANDX1 U11748 (.A1(N3666), .A2(n20751), .ZN(n24620));
    INVX1 U11749 (.I(n14930), .ZN(N24621));
    NOR2X1 U11750 (.A1(N4939), .A2(n17013), .ZN(N24622));
    NOR2X1 U11751 (.A1(N10774), .A2(n15762), .ZN(n24623));
    NOR2X1 U11752 (.A1(n17281), .A2(N11620), .ZN(N24624));
    INVX1 U11753 (.I(N2161), .ZN(n24625));
    NANDX1 U11754 (.A1(n20095), .A2(N709), .ZN(n24626));
    NANDX1 U11755 (.A1(N7168), .A2(N4273), .ZN(n24627));
    INVX1 U11756 (.I(n14035), .ZN(N24628));
    INVX1 U11757 (.I(N3738), .ZN(n24629));
    NANDX1 U11758 (.A1(n15979), .A2(n13903), .ZN(n24630));
    NOR2X1 U11759 (.A1(n18444), .A2(N9901), .ZN(n24631));
    NANDX1 U11760 (.A1(n17965), .A2(N2635), .ZN(n24632));
    NANDX1 U11761 (.A1(N3877), .A2(N7573), .ZN(N24633));
    NOR2X1 U11762 (.A1(N9698), .A2(n12889), .ZN(n24634));
    INVX1 U11763 (.I(n16368), .ZN(n24635));
    NOR2X1 U11764 (.A1(N2000), .A2(N9381), .ZN(n24636));
    NANDX1 U11765 (.A1(N11074), .A2(N8245), .ZN(n24637));
    NOR2X1 U11766 (.A1(n18849), .A2(n15413), .ZN(N24638));
    INVX1 U11767 (.I(n20583), .ZN(n24639));
    INVX1 U11768 (.I(N2767), .ZN(n24640));
    NANDX1 U11769 (.A1(N10687), .A2(n18745), .ZN(n24641));
    NOR2X1 U11770 (.A1(n18846), .A2(n15959), .ZN(N24642));
    NANDX1 U11771 (.A1(N9440), .A2(N12693), .ZN(n24643));
    NOR2X1 U11772 (.A1(N9505), .A2(N11111), .ZN(N24644));
    NANDX1 U11773 (.A1(N5353), .A2(n15350), .ZN(n24645));
    NANDX1 U11774 (.A1(n16963), .A2(N10487), .ZN(N24646));
    NOR2X1 U11775 (.A1(n13504), .A2(n19868), .ZN(N24647));
    INVX1 U11776 (.I(n19119), .ZN(n24648));
    NANDX1 U11777 (.A1(N564), .A2(N11279), .ZN(n24649));
    NANDX1 U11778 (.A1(n16041), .A2(N5173), .ZN(N24650));
    NOR2X1 U11779 (.A1(n18807), .A2(N2805), .ZN(N24651));
    INVX1 U11780 (.I(N10863), .ZN(n24652));
    INVX1 U11781 (.I(N11522), .ZN(n24653));
    NANDX1 U11782 (.A1(n19398), .A2(n15503), .ZN(n24654));
    INVX1 U11783 (.I(N11320), .ZN(n24655));
    INVX1 U11784 (.I(n13019), .ZN(n24656));
    INVX1 U11785 (.I(N3672), .ZN(N24657));
    NANDX1 U11786 (.A1(N6823), .A2(n15176), .ZN(n24658));
    NOR2X1 U11787 (.A1(N6312), .A2(N1991), .ZN(n24659));
    NANDX1 U11788 (.A1(N5984), .A2(n15651), .ZN(n24660));
    NANDX1 U11789 (.A1(N1089), .A2(N5699), .ZN(n24661));
    NOR2X1 U11790 (.A1(n17129), .A2(N10872), .ZN(n24662));
    INVX1 U11791 (.I(N9247), .ZN(N24663));
    NOR2X1 U11792 (.A1(n14043), .A2(n20109), .ZN(n24664));
    INVX1 U11793 (.I(N4334), .ZN(n24665));
    INVX1 U11794 (.I(N9806), .ZN(n24666));
    INVX1 U11795 (.I(n16692), .ZN(n24667));
    INVX1 U11796 (.I(N7238), .ZN(n24668));
    INVX1 U11797 (.I(n15565), .ZN(n24669));
    INVX1 U11798 (.I(N10161), .ZN(n24670));
    INVX1 U11799 (.I(n20626), .ZN(n24671));
    NANDX1 U11800 (.A1(N2010), .A2(n17158), .ZN(n24672));
    NANDX1 U11801 (.A1(N7993), .A2(N11578), .ZN(n24673));
    NOR2X1 U11802 (.A1(N3623), .A2(n17277), .ZN(n24674));
    NOR2X1 U11803 (.A1(n20751), .A2(N1460), .ZN(N24675));
    NOR2X1 U11804 (.A1(N8767), .A2(N4219), .ZN(n24676));
    NOR2X1 U11805 (.A1(N7645), .A2(n15857), .ZN(n24677));
    INVX1 U11806 (.I(n16970), .ZN(n24678));
    NANDX1 U11807 (.A1(N10870), .A2(N12432), .ZN(n24679));
    NOR2X1 U11808 (.A1(n18108), .A2(n15454), .ZN(n24680));
    NANDX1 U11809 (.A1(N2328), .A2(N4384), .ZN(n24681));
    NANDX1 U11810 (.A1(n17496), .A2(N10938), .ZN(n24682));
    NOR2X1 U11811 (.A1(n13423), .A2(n17380), .ZN(n24683));
    NANDX1 U11812 (.A1(N3771), .A2(N9361), .ZN(n24684));
    NOR2X1 U11813 (.A1(n15589), .A2(n19489), .ZN(n24685));
    INVX1 U11814 (.I(N11590), .ZN(n24686));
    INVX1 U11815 (.I(N10208), .ZN(n24687));
    NANDX1 U11816 (.A1(N6140), .A2(N12395), .ZN(n24688));
    NANDX1 U11817 (.A1(N2632), .A2(N2676), .ZN(n24689));
    INVX1 U11818 (.I(n13502), .ZN(n24690));
    NANDX1 U11819 (.A1(N2217), .A2(N4921), .ZN(n24691));
    NOR2X1 U11820 (.A1(N5733), .A2(N7248), .ZN(n24692));
    NOR2X1 U11821 (.A1(n20720), .A2(N3513), .ZN(n24693));
    NOR2X1 U11822 (.A1(N11027), .A2(N11478), .ZN(n24694));
    INVX1 U11823 (.I(N9327), .ZN(n24695));
    NOR2X1 U11824 (.A1(n19245), .A2(N5790), .ZN(N24696));
    NANDX1 U11825 (.A1(n17503), .A2(N1774), .ZN(n24697));
    NANDX1 U11826 (.A1(n20566), .A2(N6523), .ZN(n24698));
    INVX1 U11827 (.I(N17), .ZN(n24699));
    INVX1 U11828 (.I(n20145), .ZN(n24700));
    NOR2X1 U11829 (.A1(n16135), .A2(n18637), .ZN(n24701));
    INVX1 U11830 (.I(N10011), .ZN(n24702));
    NANDX1 U11831 (.A1(N10154), .A2(n13883), .ZN(n24703));
    NANDX1 U11832 (.A1(n17401), .A2(N907), .ZN(n24704));
    NANDX1 U11833 (.A1(n15456), .A2(n14641), .ZN(n24705));
    NANDX1 U11834 (.A1(N5703), .A2(N3295), .ZN(N24706));
    INVX1 U11835 (.I(N10034), .ZN(n24707));
    NANDX1 U11836 (.A1(N9154), .A2(n14181), .ZN(n24708));
    INVX1 U11837 (.I(N10927), .ZN(n24709));
    NOR2X1 U11838 (.A1(N7230), .A2(n17450), .ZN(n24710));
    INVX1 U11839 (.I(N1789), .ZN(N24711));
    NOR2X1 U11840 (.A1(N11854), .A2(n20209), .ZN(n24712));
    NOR2X1 U11841 (.A1(N3802), .A2(N4212), .ZN(n24713));
    NOR2X1 U11842 (.A1(n19196), .A2(n14365), .ZN(n24714));
    NANDX1 U11843 (.A1(n13635), .A2(N5077), .ZN(N24715));
    NANDX1 U11844 (.A1(N7562), .A2(n15074), .ZN(n24716));
    NANDX1 U11845 (.A1(N7058), .A2(n15318), .ZN(N24717));
    NOR2X1 U11846 (.A1(n15880), .A2(N4121), .ZN(n24718));
    INVX1 U11847 (.I(n19576), .ZN(n24719));
    NOR2X1 U11848 (.A1(n18914), .A2(N9272), .ZN(n24720));
    NOR2X1 U11849 (.A1(N4913), .A2(N5491), .ZN(n24721));
    NOR2X1 U11850 (.A1(N6701), .A2(N9711), .ZN(n24722));
    NOR2X1 U11851 (.A1(N221), .A2(n14292), .ZN(n24723));
    NOR2X1 U11852 (.A1(N4432), .A2(N2196), .ZN(N24724));
    INVX1 U11853 (.I(n13338), .ZN(n24725));
    NANDX1 U11854 (.A1(n18661), .A2(n12957), .ZN(n24726));
    NANDX1 U11855 (.A1(N4992), .A2(N6800), .ZN(n24727));
    NOR2X1 U11856 (.A1(N6592), .A2(n16660), .ZN(n24728));
    NANDX1 U11857 (.A1(n17013), .A2(n20780), .ZN(n24729));
    NOR2X1 U11858 (.A1(n15358), .A2(N6935), .ZN(n24730));
    NANDX1 U11859 (.A1(N3400), .A2(N12089), .ZN(n24731));
    NANDX1 U11860 (.A1(N3432), .A2(N8953), .ZN(N24732));
    INVX1 U11861 (.I(n13142), .ZN(n24733));
    INVX1 U11862 (.I(n16048), .ZN(n24734));
    INVX1 U11863 (.I(N3500), .ZN(n24735));
    NANDX1 U11864 (.A1(N2941), .A2(N3068), .ZN(N24736));
    NANDX1 U11865 (.A1(n17237), .A2(N498), .ZN(n24737));
    INVX1 U11866 (.I(N7537), .ZN(n24738));
    INVX1 U11867 (.I(N197), .ZN(N24739));
    NANDX1 U11868 (.A1(N6623), .A2(n16856), .ZN(n24740));
    INVX1 U11869 (.I(N2405), .ZN(n24741));
    INVX1 U11870 (.I(N1441), .ZN(N24742));
    NANDX1 U11871 (.A1(N12423), .A2(N11113), .ZN(n24743));
    NOR2X1 U11872 (.A1(N3282), .A2(n20239), .ZN(n24744));
    INVX1 U11873 (.I(N6776), .ZN(n24745));
    NANDX1 U11874 (.A1(N11047), .A2(n18987), .ZN(n24746));
    NOR2X1 U11875 (.A1(N11792), .A2(n17028), .ZN(N24747));
    NANDX1 U11876 (.A1(n14732), .A2(n20096), .ZN(n24748));
    INVX1 U11877 (.I(N5280), .ZN(N24749));
    NANDX1 U11878 (.A1(n14284), .A2(N12816), .ZN(n24750));
    NANDX1 U11879 (.A1(N9022), .A2(N11611), .ZN(n24751));
    NOR2X1 U11880 (.A1(n20419), .A2(n16834), .ZN(N24752));
    INVX1 U11881 (.I(N10135), .ZN(n24753));
    INVX1 U11882 (.I(n15267), .ZN(n24754));
    INVX1 U11883 (.I(N2698), .ZN(n24755));
    NANDX1 U11884 (.A1(n20381), .A2(N1707), .ZN(n24756));
    NANDX1 U11885 (.A1(N5926), .A2(N11084), .ZN(N24757));
    NANDX1 U11886 (.A1(N3682), .A2(N9821), .ZN(n24758));
    NOR2X1 U11887 (.A1(n20709), .A2(n18121), .ZN(n24759));
    NOR2X1 U11888 (.A1(n14116), .A2(N12320), .ZN(n24760));
    NANDX1 U11889 (.A1(n13479), .A2(N5373), .ZN(N24761));
    INVX1 U11890 (.I(N7414), .ZN(n24762));
    NOR2X1 U11891 (.A1(n16084), .A2(N2514), .ZN(n24763));
    NANDX1 U11892 (.A1(N11688), .A2(N5476), .ZN(n24764));
    NANDX1 U11893 (.A1(N3273), .A2(n15284), .ZN(n24765));
    NANDX1 U11894 (.A1(N5971), .A2(N3793), .ZN(n24766));
    NOR2X1 U11895 (.A1(N2219), .A2(N5978), .ZN(n24767));
    INVX1 U11896 (.I(N7844), .ZN(n24768));
    NANDX1 U11897 (.A1(N6509), .A2(N12207), .ZN(n24769));
    NANDX1 U11898 (.A1(N530), .A2(N9097), .ZN(n24770));
    NANDX1 U11899 (.A1(n14645), .A2(N186), .ZN(n24771));
    INVX1 U11900 (.I(N1435), .ZN(n24772));
    INVX1 U11901 (.I(N6113), .ZN(n24773));
    NOR2X1 U11902 (.A1(N9035), .A2(N966), .ZN(n24774));
    NANDX1 U11903 (.A1(N11700), .A2(N7195), .ZN(N24775));
    NANDX1 U11904 (.A1(n19042), .A2(N10468), .ZN(N24776));
    INVX1 U11905 (.I(N1022), .ZN(N24777));
    INVX1 U11906 (.I(n19538), .ZN(n24778));
    INVX1 U11907 (.I(N7740), .ZN(n24779));
    INVX1 U11908 (.I(N6210), .ZN(n24780));
    INVX1 U11909 (.I(N7722), .ZN(n24781));
    NOR2X1 U11910 (.A1(N6559), .A2(N9494), .ZN(N24782));
    NOR2X1 U11911 (.A1(N10198), .A2(N8559), .ZN(N24783));
    NANDX1 U11912 (.A1(N10383), .A2(N4740), .ZN(N24784));
    NOR2X1 U11913 (.A1(N5025), .A2(N10852), .ZN(N24785));
    NANDX1 U11914 (.A1(N8601), .A2(N6360), .ZN(n24786));
    INVX1 U11915 (.I(n20301), .ZN(n24787));
    NOR2X1 U11916 (.A1(N6936), .A2(N12654), .ZN(n24788));
    NOR2X1 U11917 (.A1(N1451), .A2(n13675), .ZN(n24789));
    INVX1 U11918 (.I(n20988), .ZN(n24790));
    INVX1 U11919 (.I(N10593), .ZN(n24791));
    INVX1 U11920 (.I(n17809), .ZN(n24792));
    INVX1 U11921 (.I(N6306), .ZN(n24793));
    INVX1 U11922 (.I(N588), .ZN(n24794));
    NOR2X1 U11923 (.A1(N11628), .A2(N10785), .ZN(n24795));
    NANDX1 U11924 (.A1(N7373), .A2(n15710), .ZN(n24796));
    INVX1 U11925 (.I(N4553), .ZN(n24797));
    NANDX1 U11926 (.A1(N2344), .A2(n20895), .ZN(n24798));
    INVX1 U11927 (.I(N8703), .ZN(n24799));
    NOR2X1 U11928 (.A1(N1716), .A2(n16799), .ZN(n24800));
    INVX1 U11929 (.I(n14369), .ZN(n24801));
    INVX1 U11930 (.I(N9065), .ZN(n24802));
    INVX1 U11931 (.I(N6069), .ZN(n24803));
    INVX1 U11932 (.I(n18412), .ZN(n24804));
    NANDX1 U11933 (.A1(N7406), .A2(n14990), .ZN(n24805));
    NOR2X1 U11934 (.A1(N8253), .A2(n18828), .ZN(n24806));
    INVX1 U11935 (.I(n18593), .ZN(N24807));
    INVX1 U11936 (.I(N11146), .ZN(n24808));
    INVX1 U11937 (.I(N11140), .ZN(n24809));
    NANDX1 U11938 (.A1(N7753), .A2(n15692), .ZN(n24810));
    NOR2X1 U11939 (.A1(N10097), .A2(n15357), .ZN(n24811));
    NANDX1 U11940 (.A1(n13341), .A2(N10578), .ZN(n24812));
    NANDX1 U11941 (.A1(N3451), .A2(n18193), .ZN(N24813));
    NANDX1 U11942 (.A1(N6666), .A2(N569), .ZN(N24814));
    NOR2X1 U11943 (.A1(N7276), .A2(n19705), .ZN(N24815));
    NANDX1 U11944 (.A1(n18478), .A2(N5880), .ZN(n24816));
    INVX1 U11945 (.I(n18252), .ZN(n24817));
    INVX1 U11946 (.I(n13149), .ZN(n24818));
    NANDX1 U11947 (.A1(N6036), .A2(n16916), .ZN(n24819));
    NOR2X1 U11948 (.A1(n16838), .A2(N6825), .ZN(n24820));
    NANDX1 U11949 (.A1(n19133), .A2(n17058), .ZN(n24821));
    NANDX1 U11950 (.A1(N2541), .A2(N5726), .ZN(n24822));
    INVX1 U11951 (.I(N10423), .ZN(N24823));
    NANDX1 U11952 (.A1(n14108), .A2(n13874), .ZN(N24824));
    INVX1 U11953 (.I(N5819), .ZN(n24825));
    INVX1 U11954 (.I(N2918), .ZN(N24826));
    NANDX1 U11955 (.A1(N1126), .A2(N1392), .ZN(n24827));
    NOR2X1 U11956 (.A1(n14145), .A2(N1813), .ZN(n24828));
    INVX1 U11957 (.I(N11166), .ZN(N24829));
    NOR2X1 U11958 (.A1(N1458), .A2(N8548), .ZN(N24830));
    NANDX1 U11959 (.A1(n18373), .A2(N11618), .ZN(n24831));
    NOR2X1 U11960 (.A1(n19739), .A2(n14854), .ZN(N24832));
    INVX1 U11961 (.I(n15566), .ZN(n24833));
    NANDX1 U11962 (.A1(N7113), .A2(n15834), .ZN(n24834));
    INVX1 U11963 (.I(n17535), .ZN(n24835));
    NANDX1 U11964 (.A1(n20713), .A2(N4720), .ZN(n24836));
    NANDX1 U11965 (.A1(n21073), .A2(n19800), .ZN(n24837));
    NANDX1 U11966 (.A1(N9041), .A2(n15467), .ZN(n24838));
    NANDX1 U11967 (.A1(N3028), .A2(N2924), .ZN(n24839));
    NOR2X1 U11968 (.A1(n18025), .A2(N8631), .ZN(N24840));
    INVX1 U11969 (.I(n14024), .ZN(n24841));
    NANDX1 U11970 (.A1(n14237), .A2(N5708), .ZN(n24842));
    NANDX1 U11971 (.A1(n20907), .A2(N4216), .ZN(n24843));
    NANDX1 U11972 (.A1(n20021), .A2(n14323), .ZN(N24844));
    INVX1 U11973 (.I(N445), .ZN(n24845));
    INVX1 U11974 (.I(N3720), .ZN(n24846));
    NOR2X1 U11975 (.A1(N8916), .A2(n18974), .ZN(N24847));
    NOR2X1 U11976 (.A1(n16713), .A2(n18816), .ZN(N24848));
    INVX1 U11977 (.I(N6198), .ZN(n24849));
    NOR2X1 U11978 (.A1(N4589), .A2(n18304), .ZN(n24850));
    NANDX1 U11979 (.A1(N2054), .A2(N5534), .ZN(n24851));
    NANDX1 U11980 (.A1(N10685), .A2(N3250), .ZN(n24852));
    NOR2X1 U11981 (.A1(N1175), .A2(N12029), .ZN(n24853));
    INVX1 U11982 (.I(n19054), .ZN(n24854));
    NANDX1 U11983 (.A1(n19477), .A2(N3868), .ZN(N24855));
    INVX1 U11984 (.I(N7111), .ZN(N24856));
    INVX1 U11985 (.I(N5482), .ZN(n24857));
    NANDX1 U11986 (.A1(n20474), .A2(n18003), .ZN(N24858));
    NOR2X1 U11987 (.A1(n18217), .A2(n14014), .ZN(N24859));
    INVX1 U11988 (.I(N10345), .ZN(n24860));
    NANDX1 U11989 (.A1(n15716), .A2(N11512), .ZN(n24861));
    INVX1 U11990 (.I(N7331), .ZN(n24862));
    NOR2X1 U11991 (.A1(N4320), .A2(N12864), .ZN(n24863));
    INVX1 U11992 (.I(N9546), .ZN(N24864));
    INVX1 U11993 (.I(n15334), .ZN(n24865));
    NOR2X1 U11994 (.A1(n17226), .A2(N9365), .ZN(n24866));
    NANDX1 U11995 (.A1(N2242), .A2(N2153), .ZN(n24867));
    NANDX1 U11996 (.A1(N1821), .A2(N3806), .ZN(n24868));
    NANDX1 U11997 (.A1(N7303), .A2(n14384), .ZN(N24869));
    NANDX1 U11998 (.A1(n19847), .A2(N7189), .ZN(N24870));
    NOR2X1 U11999 (.A1(N7172), .A2(n16707), .ZN(N24871));
    NOR2X1 U12000 (.A1(N10307), .A2(N11192), .ZN(N24872));
    INVX1 U12001 (.I(N7115), .ZN(n24873));
    NOR2X1 U12002 (.A1(N4121), .A2(N5976), .ZN(n24874));
    NOR2X1 U12003 (.A1(n15358), .A2(n15521), .ZN(n24875));
    NOR2X1 U12004 (.A1(N9462), .A2(n20782), .ZN(n24876));
    NANDX1 U12005 (.A1(n13368), .A2(N2636), .ZN(N24877));
    INVX1 U12006 (.I(n15521), .ZN(n24878));
    NOR2X1 U12007 (.A1(N9952), .A2(n13868), .ZN(n24879));
    NANDX1 U12008 (.A1(N11796), .A2(N7021), .ZN(n24880));
    INVX1 U12009 (.I(N10412), .ZN(n24881));
    NOR2X1 U12010 (.A1(N1567), .A2(n17584), .ZN(n24882));
    NANDX1 U12011 (.A1(N5157), .A2(N1202), .ZN(n24883));
    NOR2X1 U12012 (.A1(n20258), .A2(N2858), .ZN(N24884));
    NOR2X1 U12013 (.A1(N3148), .A2(N3375), .ZN(N24885));
    NANDX1 U12014 (.A1(n13048), .A2(n18895), .ZN(n24886));
    NANDX1 U12015 (.A1(n17051), .A2(n12988), .ZN(N24887));
    NOR2X1 U12016 (.A1(N9188), .A2(n15623), .ZN(n24888));
    INVX1 U12017 (.I(n19250), .ZN(n24889));
    NOR2X1 U12018 (.A1(N3354), .A2(N11887), .ZN(N24890));
    NANDX1 U12019 (.A1(N9691), .A2(n13449), .ZN(n24891));
    NANDX1 U12020 (.A1(n14645), .A2(N970), .ZN(n24892));
    NANDX1 U12021 (.A1(N5540), .A2(N5197), .ZN(n24893));
    NANDX1 U12022 (.A1(N1283), .A2(n20615), .ZN(N24894));
    INVX1 U12023 (.I(n19913), .ZN(N24895));
    NOR2X1 U12024 (.A1(N5967), .A2(N2057), .ZN(N24896));
    INVX1 U12025 (.I(n19014), .ZN(n24897));
    NANDX1 U12026 (.A1(N3427), .A2(n14834), .ZN(n24898));
    INVX1 U12027 (.I(n15387), .ZN(n24899));
    INVX1 U12028 (.I(N1644), .ZN(n24900));
    NOR2X1 U12029 (.A1(n16583), .A2(N10478), .ZN(n24901));
    NANDX1 U12030 (.A1(N1781), .A2(N10143), .ZN(n24902));
    INVX1 U12031 (.I(n15230), .ZN(N24903));
    NANDX1 U12032 (.A1(n20104), .A2(n16199), .ZN(n24904));
    INVX1 U12033 (.I(N4413), .ZN(n24905));
    INVX1 U12034 (.I(N4782), .ZN(n24906));
    NANDX1 U12035 (.A1(n15321), .A2(N7601), .ZN(n24907));
    NOR2X1 U12036 (.A1(N728), .A2(n13567), .ZN(n24908));
    NANDX1 U12037 (.A1(n19313), .A2(N11350), .ZN(n24909));
    INVX1 U12038 (.I(N1510), .ZN(n24910));
    NANDX1 U12039 (.A1(N7947), .A2(N11438), .ZN(n24911));
    NANDX1 U12040 (.A1(N4132), .A2(n14769), .ZN(n24912));
    NOR2X1 U12041 (.A1(N9152), .A2(n15996), .ZN(n24913));
    NANDX1 U12042 (.A1(n19294), .A2(N5683), .ZN(n24914));
    NOR2X1 U12043 (.A1(N5276), .A2(N4556), .ZN(n24915));
    INVX1 U12044 (.I(N808), .ZN(n24916));
    NANDX1 U12045 (.A1(n14635), .A2(N5590), .ZN(N24917));
    NOR2X1 U12046 (.A1(N3267), .A2(n13190), .ZN(n24918));
    INVX1 U12047 (.I(N3994), .ZN(n24919));
    INVX1 U12048 (.I(n19412), .ZN(n24920));
    NANDX1 U12049 (.A1(N5959), .A2(n14650), .ZN(n24921));
    NOR2X1 U12050 (.A1(N5453), .A2(n17138), .ZN(N24922));
    INVX1 U12051 (.I(n18051), .ZN(n24923));
    INVX1 U12052 (.I(n18876), .ZN(n24924));
    NOR2X1 U12053 (.A1(N3733), .A2(n13641), .ZN(n24925));
    NANDX1 U12054 (.A1(N1796), .A2(n13865), .ZN(n24926));
    NANDX1 U12055 (.A1(N7071), .A2(n12962), .ZN(N24927));
    NANDX1 U12056 (.A1(N2421), .A2(n16471), .ZN(n24928));
    NOR2X1 U12057 (.A1(N2552), .A2(n14758), .ZN(N24929));
    INVX1 U12058 (.I(N10283), .ZN(n24930));
    INVX1 U12059 (.I(N11535), .ZN(n24931));
    INVX1 U12060 (.I(N10145), .ZN(n24932));
    NANDX1 U12061 (.A1(n16308), .A2(n19336), .ZN(N24933));
    NANDX1 U12062 (.A1(n16302), .A2(n15244), .ZN(n24934));
    NANDX1 U12063 (.A1(N7664), .A2(N4367), .ZN(n24935));
    INVX1 U12064 (.I(N12435), .ZN(n24936));
    INVX1 U12065 (.I(N10755), .ZN(N24937));
    NANDX1 U12066 (.A1(N4436), .A2(N3389), .ZN(N24938));
    NOR2X1 U12067 (.A1(N6049), .A2(n16350), .ZN(N24939));
    INVX1 U12068 (.I(N8469), .ZN(n24940));
    INVX1 U12069 (.I(N12395), .ZN(N24941));
    NOR2X1 U12070 (.A1(n20890), .A2(n19936), .ZN(n24942));
    NOR2X1 U12071 (.A1(N6165), .A2(N10240), .ZN(N24943));
    NOR2X1 U12072 (.A1(N10852), .A2(n12934), .ZN(n24944));
    NOR2X1 U12073 (.A1(N8957), .A2(n13755), .ZN(N24945));
    INVX1 U12074 (.I(n18742), .ZN(N24946));
    INVX1 U12075 (.I(n13088), .ZN(n24947));
    NANDX1 U12076 (.A1(N10339), .A2(n20065), .ZN(n24948));
    NOR2X1 U12077 (.A1(n15635), .A2(n14855), .ZN(n24949));
    NANDX1 U12078 (.A1(n19024), .A2(N11504), .ZN(N24950));
    NOR2X1 U12079 (.A1(N8685), .A2(n14166), .ZN(n24951));
    NOR2X1 U12080 (.A1(N9359), .A2(n21103), .ZN(n24952));
    NANDX1 U12081 (.A1(N3560), .A2(n19808), .ZN(n24953));
    INVX1 U12082 (.I(N9724), .ZN(N24954));
    INVX1 U12083 (.I(n17690), .ZN(n24955));
    INVX1 U12084 (.I(n16292), .ZN(N24956));
    INVX1 U12085 (.I(N2844), .ZN(n24957));
    INVX1 U12086 (.I(N12237), .ZN(n24958));
    NOR2X1 U12087 (.A1(n16581), .A2(n19866), .ZN(n24959));
    NOR2X1 U12088 (.A1(N231), .A2(n18700), .ZN(n24960));
    NANDX1 U12089 (.A1(n15866), .A2(N6867), .ZN(n24961));
    NOR2X1 U12090 (.A1(N8201), .A2(n18370), .ZN(n24962));
    NOR2X1 U12091 (.A1(N11427), .A2(N11305), .ZN(n24963));
    NANDX1 U12092 (.A1(n20785), .A2(N5719), .ZN(N24964));
    NOR2X1 U12093 (.A1(N3114), .A2(N4296), .ZN(n24965));
    INVX1 U12094 (.I(N7380), .ZN(n24966));
    NOR2X1 U12095 (.A1(N1409), .A2(N1266), .ZN(n24967));
    INVX1 U12096 (.I(N2763), .ZN(N24968));
    INVX1 U12097 (.I(N6072), .ZN(N24969));
    NANDX1 U12098 (.A1(n14778), .A2(n17195), .ZN(n24970));
    INVX1 U12099 (.I(N6094), .ZN(n24971));
    NANDX1 U12100 (.A1(N5646), .A2(n17699), .ZN(n24972));
    NOR2X1 U12101 (.A1(N12512), .A2(n17028), .ZN(N24973));
    NOR2X1 U12102 (.A1(N4193), .A2(N10127), .ZN(n24974));
    NANDX1 U12103 (.A1(N10040), .A2(n15780), .ZN(N24975));
    INVX1 U12104 (.I(n15758), .ZN(n24976));
    NANDX1 U12105 (.A1(N12523), .A2(n20054), .ZN(n24977));
    NOR2X1 U12106 (.A1(n19902), .A2(N1019), .ZN(N24978));
    INVX1 U12107 (.I(n21167), .ZN(N24979));
    NOR2X1 U12108 (.A1(N749), .A2(n19818), .ZN(n24980));
    NOR2X1 U12109 (.A1(n15747), .A2(N7907), .ZN(n24981));
    NOR2X1 U12110 (.A1(N2693), .A2(N8542), .ZN(n24982));
    NANDX1 U12111 (.A1(N2881), .A2(N5010), .ZN(N24983));
    NANDX1 U12112 (.A1(N9934), .A2(n16579), .ZN(n24984));
    NANDX1 U12113 (.A1(n14127), .A2(N5476), .ZN(n24985));
    INVX1 U12114 (.I(n18708), .ZN(n24986));
    NANDX1 U12115 (.A1(N10483), .A2(n13235), .ZN(n24987));
    NOR2X1 U12116 (.A1(N1775), .A2(N6600), .ZN(n24988));
    NOR2X1 U12117 (.A1(N446), .A2(N7619), .ZN(n24989));
    NANDX1 U12118 (.A1(n16155), .A2(N5894), .ZN(N24990));
    NANDX1 U12119 (.A1(N9284), .A2(n15698), .ZN(n24991));
    INVX1 U12120 (.I(n17190), .ZN(N24992));
    NOR2X1 U12121 (.A1(N5402), .A2(n20273), .ZN(n24993));
    NANDX1 U12122 (.A1(N8282), .A2(N4052), .ZN(n24994));
    NOR2X1 U12123 (.A1(N12757), .A2(n20631), .ZN(n24995));
    NANDX1 U12124 (.A1(N5653), .A2(n20648), .ZN(n24996));
    NANDX1 U12125 (.A1(n18902), .A2(N9756), .ZN(n24997));
    INVX1 U12126 (.I(N10907), .ZN(n24998));
    NANDX1 U12127 (.A1(N8653), .A2(N12048), .ZN(n24999));
    NOR2X1 U12128 (.A1(N3641), .A2(n19666), .ZN(n25000));
    NANDX1 U12129 (.A1(n19795), .A2(N4329), .ZN(n25001));
    NOR2X1 U12130 (.A1(N2390), .A2(n14569), .ZN(n25002));
    INVX1 U12131 (.I(n19579), .ZN(N25003));
    INVX1 U12132 (.I(n19441), .ZN(n25004));
    NOR2X1 U12133 (.A1(N5486), .A2(N1034), .ZN(n25005));
    NOR2X1 U12134 (.A1(n20503), .A2(n13791), .ZN(N25006));
    INVX1 U12135 (.I(N53), .ZN(n25007));
    NOR2X1 U12136 (.A1(N5115), .A2(n17678), .ZN(n25008));
    INVX1 U12137 (.I(n14870), .ZN(n25009));
    INVX1 U12138 (.I(n17105), .ZN(n25010));
    INVX1 U12139 (.I(N11979), .ZN(n25011));
    INVX1 U12140 (.I(N11370), .ZN(N25012));
    NANDX1 U12141 (.A1(N900), .A2(N3593), .ZN(n25013));
    NOR2X1 U12142 (.A1(n21000), .A2(n14924), .ZN(n25014));
    INVX1 U12143 (.I(n14338), .ZN(n25015));
    INVX1 U12144 (.I(N4004), .ZN(N25016));
    NOR2X1 U12145 (.A1(N486), .A2(n17166), .ZN(N25017));
    NANDX1 U12146 (.A1(N1519), .A2(n13149), .ZN(n25018));
    NANDX1 U12147 (.A1(N9851), .A2(n18847), .ZN(n25019));
    NANDX1 U12148 (.A1(N2606), .A2(n18503), .ZN(n25020));
    INVX1 U12149 (.I(N8804), .ZN(N25021));
    NOR2X1 U12150 (.A1(N6435), .A2(N4678), .ZN(n25022));
    INVX1 U12151 (.I(n12955), .ZN(n25023));
    NOR2X1 U12152 (.A1(n13100), .A2(N7343), .ZN(n25024));
    INVX1 U12153 (.I(n16692), .ZN(n25025));
    NANDX1 U12154 (.A1(N7810), .A2(N4927), .ZN(n25026));
    NANDX1 U12155 (.A1(n16689), .A2(N7201), .ZN(n25027));
    NOR2X1 U12156 (.A1(N2769), .A2(N7686), .ZN(n25028));
    INVX1 U12157 (.I(n15563), .ZN(n25029));
    INVX1 U12158 (.I(n13578), .ZN(n25030));
    INVX1 U12159 (.I(n13597), .ZN(n25031));
    NANDX1 U12160 (.A1(N2145), .A2(N10744), .ZN(n25032));
    INVX1 U12161 (.I(n21026), .ZN(N25033));
    INVX1 U12162 (.I(N9693), .ZN(n25034));
    INVX1 U12163 (.I(n18766), .ZN(n25035));
    INVX1 U12164 (.I(n13726), .ZN(n25036));
    NOR2X1 U12165 (.A1(n19064), .A2(n21068), .ZN(n25037));
    NOR2X1 U12166 (.A1(n14525), .A2(N10446), .ZN(n25038));
    INVX1 U12167 (.I(n19451), .ZN(n25039));
    INVX1 U12168 (.I(N5068), .ZN(n25040));
    NOR2X1 U12169 (.A1(n20889), .A2(N7836), .ZN(n25041));
    INVX1 U12170 (.I(N88), .ZN(N25042));
    INVX1 U12171 (.I(N11395), .ZN(n25043));
    INVX1 U12172 (.I(n13424), .ZN(n25044));
    NANDX1 U12173 (.A1(n13943), .A2(n15568), .ZN(N25045));
    NANDX1 U12174 (.A1(N11493), .A2(n15363), .ZN(n25046));
    NANDX1 U12175 (.A1(n21185), .A2(N10676), .ZN(n25047));
    NANDX1 U12176 (.A1(N5919), .A2(N3171), .ZN(n25048));
    INVX1 U12177 (.I(N3752), .ZN(n25049));
    NANDX1 U12178 (.A1(N10772), .A2(N12818), .ZN(n25050));
    NANDX1 U12179 (.A1(n20381), .A2(N5580), .ZN(n25051));
    NANDX1 U12180 (.A1(N4218), .A2(N5542), .ZN(n25052));
    NOR2X1 U12181 (.A1(N12053), .A2(N7732), .ZN(n25053));
    NANDX1 U12182 (.A1(N3304), .A2(n19126), .ZN(N25054));
    NOR2X1 U12183 (.A1(n16727), .A2(N11971), .ZN(n25055));
    NOR2X1 U12184 (.A1(N5607), .A2(N10101), .ZN(n25056));
    NOR2X1 U12185 (.A1(n15511), .A2(N6547), .ZN(N25057));
    INVX1 U12186 (.I(N4957), .ZN(n25058));
    INVX1 U12187 (.I(n15127), .ZN(n25059));
    INVX1 U12188 (.I(n19815), .ZN(n25060));
    NANDX1 U12189 (.A1(N5677), .A2(N9357), .ZN(n25061));
    NANDX1 U12190 (.A1(n13671), .A2(N8507), .ZN(N25062));
    NOR2X1 U12191 (.A1(N11372), .A2(N7266), .ZN(n25063));
    INVX1 U12192 (.I(N8730), .ZN(N25064));
    NANDX1 U12193 (.A1(n18401), .A2(N718), .ZN(n25065));
    INVX1 U12194 (.I(N10838), .ZN(N25066));
    NOR2X1 U12195 (.A1(N7202), .A2(N1578), .ZN(N25067));
    NANDX1 U12196 (.A1(N12808), .A2(N11678), .ZN(n25068));
    NANDX1 U12197 (.A1(N7088), .A2(N12767), .ZN(N25069));
    NANDX1 U12198 (.A1(N12044), .A2(N2379), .ZN(n25070));
    INVX1 U12199 (.I(n14713), .ZN(n25071));
    NANDX1 U12200 (.A1(n19595), .A2(n20389), .ZN(n25072));
    NOR2X1 U12201 (.A1(N3371), .A2(N7371), .ZN(n25073));
    INVX1 U12202 (.I(N8498), .ZN(n25074));
    INVX1 U12203 (.I(n15175), .ZN(n25075));
    INVX1 U12204 (.I(N784), .ZN(n25076));
    INVX1 U12205 (.I(n16336), .ZN(n25077));
    NOR2X1 U12206 (.A1(n19508), .A2(N5944), .ZN(n25078));
    NOR2X1 U12207 (.A1(N5479), .A2(N2063), .ZN(N25079));
    INVX1 U12208 (.I(n18286), .ZN(N25080));
    NOR2X1 U12209 (.A1(N3554), .A2(n19916), .ZN(n25081));
    NANDX1 U12210 (.A1(N10375), .A2(N5271), .ZN(n25082));
    NANDX1 U12211 (.A1(N11092), .A2(n19983), .ZN(n25083));
    NOR2X1 U12212 (.A1(N3998), .A2(n13683), .ZN(n25084));
    NANDX1 U12213 (.A1(N7368), .A2(n21054), .ZN(n25085));
    NOR2X1 U12214 (.A1(N10407), .A2(n13107), .ZN(n25086));
    NANDX1 U12215 (.A1(N2884), .A2(N8432), .ZN(n25087));
    NOR2X1 U12216 (.A1(n13762), .A2(N4474), .ZN(N25088));
    NANDX1 U12217 (.A1(n19705), .A2(N11741), .ZN(n25089));
    NOR2X1 U12218 (.A1(n16309), .A2(n17681), .ZN(n25090));
    INVX1 U12219 (.I(N3361), .ZN(N25091));
    NOR2X1 U12220 (.A1(N11114), .A2(n18951), .ZN(N25092));
    NANDX1 U12221 (.A1(n16384), .A2(n15690), .ZN(n25093));
    INVX1 U12222 (.I(N9679), .ZN(n25094));
    NANDX1 U12223 (.A1(n20008), .A2(N2131), .ZN(n25095));
    NANDX1 U12224 (.A1(N687), .A2(n17726), .ZN(n25096));
    INVX1 U12225 (.I(N5635), .ZN(n25097));
    INVX1 U12226 (.I(N8407), .ZN(n25098));
    NOR2X1 U12227 (.A1(n18034), .A2(N4251), .ZN(n25099));
    NANDX1 U12228 (.A1(n17050), .A2(n14145), .ZN(n25100));
    NOR2X1 U12229 (.A1(N2102), .A2(N8288), .ZN(n25101));
    NOR2X1 U12230 (.A1(n19783), .A2(n20716), .ZN(n25102));
    NANDX1 U12231 (.A1(n14328), .A2(N5141), .ZN(n25103));
    NOR2X1 U12232 (.A1(n13790), .A2(N294), .ZN(n25104));
    NOR2X1 U12233 (.A1(N8570), .A2(N4514), .ZN(n25105));
    NANDX1 U12234 (.A1(N1890), .A2(N6645), .ZN(n25106));
    INVX1 U12235 (.I(N2576), .ZN(n25107));
    NOR2X1 U12236 (.A1(N11958), .A2(N8211), .ZN(n25108));
    INVX1 U12237 (.I(n14906), .ZN(n25109));
    NOR2X1 U12238 (.A1(n19860), .A2(n19157), .ZN(n25110));
    INVX1 U12239 (.I(N10221), .ZN(n25111));
    INVX1 U12240 (.I(N927), .ZN(n25112));
    NANDX1 U12241 (.A1(n14900), .A2(N5842), .ZN(N25113));
    INVX1 U12242 (.I(N8927), .ZN(N25114));
    NANDX1 U12243 (.A1(n14286), .A2(N8609), .ZN(N25115));
    NANDX1 U12244 (.A1(N6845), .A2(N8903), .ZN(n25116));
    INVX1 U12245 (.I(n15414), .ZN(n25117));
    NANDX1 U12246 (.A1(N11982), .A2(n17303), .ZN(N25118));
    NOR2X1 U12247 (.A1(N3575), .A2(n14421), .ZN(n25119));
    INVX1 U12248 (.I(N10075), .ZN(N25120));
    NANDX1 U12249 (.A1(n14109), .A2(N3750), .ZN(N25121));
    INVX1 U12250 (.I(N12738), .ZN(N25122));
    NANDX1 U12251 (.A1(n14074), .A2(N1728), .ZN(N25123));
    NOR2X1 U12252 (.A1(n15000), .A2(N8592), .ZN(n25124));
    NOR2X1 U12253 (.A1(n20841), .A2(n14007), .ZN(n25125));
    INVX1 U12254 (.I(N8271), .ZN(n25126));
    NOR2X1 U12255 (.A1(N3119), .A2(N12011), .ZN(n25127));
    INVX1 U12256 (.I(N6563), .ZN(n25128));
    NOR2X1 U12257 (.A1(N2632), .A2(n14521), .ZN(n25129));
    INVX1 U12258 (.I(n14476), .ZN(n25130));
    INVX1 U12259 (.I(N9930), .ZN(n25131));
    NANDX1 U12260 (.A1(n14717), .A2(n20004), .ZN(N25132));
    INVX1 U12261 (.I(N7596), .ZN(n25133));
    NANDX1 U12262 (.A1(N5362), .A2(n14875), .ZN(n25134));
    INVX1 U12263 (.I(n19435), .ZN(N25135));
    NOR2X1 U12264 (.A1(N11885), .A2(n13204), .ZN(N25136));
    NANDX1 U12265 (.A1(N2927), .A2(N7357), .ZN(n25137));
    INVX1 U12266 (.I(n13209), .ZN(n25138));
    NANDX1 U12267 (.A1(n14116), .A2(n16327), .ZN(n25139));
    INVX1 U12268 (.I(N1333), .ZN(n25140));
    NANDX1 U12269 (.A1(n16552), .A2(N3964), .ZN(n25141));
    NANDX1 U12270 (.A1(N7135), .A2(n12982), .ZN(n25142));
    NANDX1 U12271 (.A1(n17065), .A2(n15189), .ZN(N25143));
    INVX1 U12272 (.I(N10380), .ZN(N25144));
    NOR2X1 U12273 (.A1(N8779), .A2(N7445), .ZN(n25145));
    NOR2X1 U12274 (.A1(n18195), .A2(N728), .ZN(n25146));
    NOR2X1 U12275 (.A1(N8109), .A2(N12612), .ZN(n25147));
    NOR2X1 U12276 (.A1(N6614), .A2(N10080), .ZN(n25148));
    INVX1 U12277 (.I(n13668), .ZN(n25149));
    NOR2X1 U12278 (.A1(N10028), .A2(N6553), .ZN(n25150));
    NOR2X1 U12279 (.A1(N5518), .A2(N7885), .ZN(n25151));
    INVX1 U12280 (.I(n16612), .ZN(n25152));
    NOR2X1 U12281 (.A1(n14391), .A2(N2516), .ZN(n25153));
    NANDX1 U12282 (.A1(N6315), .A2(n14122), .ZN(n25154));
    NOR2X1 U12283 (.A1(N2040), .A2(N3272), .ZN(n25155));
    NANDX1 U12284 (.A1(N5360), .A2(N5258), .ZN(n25156));
    NOR2X1 U12285 (.A1(N2325), .A2(N5985), .ZN(N25157));
    NOR2X1 U12286 (.A1(N10433), .A2(n13139), .ZN(N25158));
    NANDX1 U12287 (.A1(N11589), .A2(N1988), .ZN(n25159));
    INVX1 U12288 (.I(N4026), .ZN(n25160));
    NOR2X1 U12289 (.A1(N11286), .A2(N5120), .ZN(n25161));
    NOR2X1 U12290 (.A1(N11346), .A2(n13004), .ZN(n25162));
    NOR2X1 U12291 (.A1(N1269), .A2(n13936), .ZN(n25163));
    NANDX1 U12292 (.A1(N3784), .A2(N12077), .ZN(n25164));
    NOR2X1 U12293 (.A1(N12448), .A2(n19949), .ZN(N25165));
    NANDX1 U12294 (.A1(N10261), .A2(n19928), .ZN(n25166));
    NOR2X1 U12295 (.A1(n15518), .A2(n17377), .ZN(n25167));
    INVX1 U12296 (.I(n16045), .ZN(n25168));
    NANDX1 U12297 (.A1(N2667), .A2(N7953), .ZN(n25169));
    NANDX1 U12298 (.A1(N8797), .A2(N4482), .ZN(N25170));
    NANDX1 U12299 (.A1(N12822), .A2(n18841), .ZN(N25171));
    NANDX1 U12300 (.A1(n17941), .A2(N3666), .ZN(N25172));
    NOR2X1 U12301 (.A1(N4256), .A2(n13390), .ZN(n25173));
    NANDX1 U12302 (.A1(N12734), .A2(N502), .ZN(n25174));
    INVX1 U12303 (.I(n19352), .ZN(n25175));
    NOR2X1 U12304 (.A1(n20538), .A2(n18070), .ZN(n25176));
    NANDX1 U12305 (.A1(N4110), .A2(n16768), .ZN(n25177));
    NANDX1 U12306 (.A1(n19627), .A2(N7456), .ZN(n25178));
    NOR2X1 U12307 (.A1(N8983), .A2(N7040), .ZN(N25179));
    NANDX1 U12308 (.A1(N11477), .A2(n18336), .ZN(n25180));
    INVX1 U12309 (.I(n15959), .ZN(N25181));
    NANDX1 U12310 (.A1(N5533), .A2(N8111), .ZN(n25182));
    NOR2X1 U12311 (.A1(n18015), .A2(N11777), .ZN(n25183));
    INVX1 U12312 (.I(n16812), .ZN(n25184));
    NOR2X1 U12313 (.A1(N9300), .A2(N8315), .ZN(n25185));
    NOR2X1 U12314 (.A1(N11932), .A2(N6437), .ZN(N25186));
    NOR2X1 U12315 (.A1(N5781), .A2(N3276), .ZN(n25187));
    INVX1 U12316 (.I(N9890), .ZN(n25188));
    NOR2X1 U12317 (.A1(N7717), .A2(N2829), .ZN(n25189));
    NOR2X1 U12318 (.A1(n15654), .A2(N11811), .ZN(N25190));
    NANDX1 U12319 (.A1(N5027), .A2(N2058), .ZN(n25191));
    NANDX1 U12320 (.A1(n18968), .A2(N12558), .ZN(N25192));
    INVX1 U12321 (.I(N3270), .ZN(N25193));
    NOR2X1 U12322 (.A1(N194), .A2(N54), .ZN(n25194));
    NANDX1 U12323 (.A1(n20959), .A2(n16866), .ZN(n25195));
    NOR2X1 U12324 (.A1(N3571), .A2(n19722), .ZN(n25196));
    NOR2X1 U12325 (.A1(n15502), .A2(N4928), .ZN(n25197));
    NANDX1 U12326 (.A1(N53), .A2(N2746), .ZN(n25198));
    NOR2X1 U12327 (.A1(N9942), .A2(n17330), .ZN(N25199));
    NANDX1 U12328 (.A1(N12770), .A2(N12682), .ZN(N25200));
    INVX1 U12329 (.I(n19123), .ZN(n25201));
    NANDX1 U12330 (.A1(n15325), .A2(n21180), .ZN(n25202));
    INVX1 U12331 (.I(n13063), .ZN(n25203));
    INVX1 U12332 (.I(n18266), .ZN(n25204));
    NOR2X1 U12333 (.A1(N1028), .A2(n18460), .ZN(n25205));
    INVX1 U12334 (.I(N1326), .ZN(n25206));
    NANDX1 U12335 (.A1(N1105), .A2(N101), .ZN(N25207));
    NANDX1 U12336 (.A1(n20826), .A2(n19085), .ZN(n25208));
    NOR2X1 U12337 (.A1(n20296), .A2(N9144), .ZN(n25209));
    NANDX1 U12338 (.A1(N1811), .A2(N1530), .ZN(N25210));
    NANDX1 U12339 (.A1(n13682), .A2(N1632), .ZN(n25211));
    INVX1 U12340 (.I(N5134), .ZN(n25212));
    NOR2X1 U12341 (.A1(n20311), .A2(n20206), .ZN(n25213));
    INVX1 U12342 (.I(n20260), .ZN(n25214));
    NOR2X1 U12343 (.A1(n13629), .A2(N620), .ZN(n25215));
    NOR2X1 U12344 (.A1(N3272), .A2(N1647), .ZN(n25216));
    INVX1 U12345 (.I(N3283), .ZN(n25217));
    NOR2X1 U12346 (.A1(N9623), .A2(N4387), .ZN(n25218));
    NANDX1 U12347 (.A1(N4692), .A2(n19755), .ZN(n25219));
    INVX1 U12348 (.I(n15263), .ZN(n25220));
    NOR2X1 U12349 (.A1(n20383), .A2(n20428), .ZN(n25221));
    NOR2X1 U12350 (.A1(N682), .A2(n14305), .ZN(n25222));
    INVX1 U12351 (.I(n18086), .ZN(n25223));
    INVX1 U12352 (.I(N7298), .ZN(n25224));
    NOR2X1 U12353 (.A1(n14573), .A2(N816), .ZN(n25225));
    INVX1 U12354 (.I(N8144), .ZN(n25226));
    NANDX1 U12355 (.A1(N1749), .A2(N8763), .ZN(n25227));
    INVX1 U12356 (.I(n20793), .ZN(n25228));
    INVX1 U12357 (.I(n15772), .ZN(N25229));
    NANDX1 U12358 (.A1(N2465), .A2(n19936), .ZN(n25230));
    INVX1 U12359 (.I(N78), .ZN(n25231));
    INVX1 U12360 (.I(n16070), .ZN(n25232));
    NOR2X1 U12361 (.A1(n13202), .A2(N8201), .ZN(N25233));
    INVX1 U12362 (.I(N6941), .ZN(n25234));
    NOR2X1 U12363 (.A1(N5694), .A2(N15), .ZN(N25235));
    INVX1 U12364 (.I(N2549), .ZN(n25236));
    NOR2X1 U12365 (.A1(N6146), .A2(N5875), .ZN(N25237));
    NOR2X1 U12366 (.A1(N6961), .A2(n15226), .ZN(N25238));
    NOR2X1 U12367 (.A1(N4946), .A2(N11516), .ZN(N25239));
    INVX1 U12368 (.I(N2594), .ZN(N25240));
    NOR2X1 U12369 (.A1(N4017), .A2(n18365), .ZN(n25241));
    NOR2X1 U12370 (.A1(N6481), .A2(N11612), .ZN(n25242));
    NOR2X1 U12371 (.A1(N6558), .A2(N9551), .ZN(n25243));
    INVX1 U12372 (.I(N12417), .ZN(n25244));
    NANDX1 U12373 (.A1(N2361), .A2(n17429), .ZN(n25245));
    NANDX1 U12374 (.A1(n20274), .A2(n17664), .ZN(n25246));
    NANDX1 U12375 (.A1(n19121), .A2(n14754), .ZN(N25247));
    NANDX1 U12376 (.A1(n19808), .A2(n20628), .ZN(n25248));
    NOR2X1 U12377 (.A1(N5538), .A2(N9165), .ZN(n25249));
    NOR2X1 U12378 (.A1(N10483), .A2(n20681), .ZN(n25250));
    INVX1 U12379 (.I(n13077), .ZN(n25251));
    NOR2X1 U12380 (.A1(N9843), .A2(N4753), .ZN(n25252));
    NANDX1 U12381 (.A1(N10865), .A2(n16365), .ZN(n25253));
    NANDX1 U12382 (.A1(n17422), .A2(n20457), .ZN(n25254));
    NANDX1 U12383 (.A1(N3151), .A2(n16520), .ZN(n25255));
    NANDX1 U12384 (.A1(n20579), .A2(n14065), .ZN(N25256));
    INVX1 U12385 (.I(N11554), .ZN(N25257));
    NANDX1 U12386 (.A1(N5707), .A2(N5077), .ZN(n25258));
    NANDX1 U12387 (.A1(n20056), .A2(n20246), .ZN(n25259));
    INVX1 U12388 (.I(N4364), .ZN(N25260));
    NANDX1 U12389 (.A1(N5449), .A2(N9388), .ZN(n25261));
    NANDX1 U12390 (.A1(N11275), .A2(n17006), .ZN(n25262));
    INVX1 U12391 (.I(n15659), .ZN(n25263));
    INVX1 U12392 (.I(N4402), .ZN(n25264));
    NANDX1 U12393 (.A1(N11435), .A2(N6340), .ZN(N25265));
    NOR2X1 U12394 (.A1(N5203), .A2(n18211), .ZN(N25266));
    NOR2X1 U12395 (.A1(N492), .A2(N11211), .ZN(N25267));
    INVX1 U12396 (.I(n14556), .ZN(N25268));
    INVX1 U12397 (.I(N4620), .ZN(n25269));
    NANDX1 U12398 (.A1(n13817), .A2(N4238), .ZN(n25270));
    INVX1 U12399 (.I(N12642), .ZN(n25271));
    INVX1 U12400 (.I(N1642), .ZN(N25272));
    NANDX1 U12401 (.A1(N11433), .A2(N1632), .ZN(n25273));
    NANDX1 U12402 (.A1(n13605), .A2(N7449), .ZN(n25274));
    INVX1 U12403 (.I(n15389), .ZN(n25275));
    NOR2X1 U12404 (.A1(N11780), .A2(n14332), .ZN(n25276));
    NANDX1 U12405 (.A1(n17756), .A2(n15213), .ZN(n25277));
    NANDX1 U12406 (.A1(N1728), .A2(N6735), .ZN(N25278));
    INVX1 U12407 (.I(n17991), .ZN(n25279));
    NOR2X1 U12408 (.A1(N5752), .A2(N5859), .ZN(n25280));
    NOR2X1 U12409 (.A1(N4913), .A2(N5351), .ZN(N25281));
    NOR2X1 U12410 (.A1(N9150), .A2(N8304), .ZN(N25282));
    NOR2X1 U12411 (.A1(N12402), .A2(N9945), .ZN(n25283));
    NOR2X1 U12412 (.A1(N2605), .A2(N6118), .ZN(n25284));
    INVX1 U12413 (.I(N10751), .ZN(N25285));
    NANDX1 U12414 (.A1(N11325), .A2(n20681), .ZN(n25286));
    NANDX1 U12415 (.A1(n17647), .A2(n13782), .ZN(n25287));
    INVX1 U12416 (.I(n14172), .ZN(N25288));
    NANDX1 U12417 (.A1(n14891), .A2(n15900), .ZN(n25289));
    INVX1 U12418 (.I(N6346), .ZN(n25290));
    NOR2X1 U12419 (.A1(N298), .A2(N12097), .ZN(n25291));
    NOR2X1 U12420 (.A1(N5123), .A2(n17009), .ZN(n25292));
    NANDX1 U12421 (.A1(N2534), .A2(N4928), .ZN(n25293));
    INVX1 U12422 (.I(N7129), .ZN(n25294));
    NOR2X1 U12423 (.A1(N9969), .A2(N7498), .ZN(N25295));
    NOR2X1 U12424 (.A1(n16087), .A2(N2113), .ZN(N25296));
    NANDX1 U12425 (.A1(N8422), .A2(n13437), .ZN(n25297));
    NOR2X1 U12426 (.A1(n18406), .A2(N9853), .ZN(n25298));
    NOR2X1 U12427 (.A1(n14329), .A2(n18567), .ZN(n25299));
    INVX1 U12428 (.I(N2531), .ZN(n25300));
    NOR2X1 U12429 (.A1(n17658), .A2(N8876), .ZN(n25301));
    NANDX1 U12430 (.A1(N12498), .A2(n15514), .ZN(n25302));
    NOR2X1 U12431 (.A1(n17620), .A2(N5834), .ZN(n25303));
    INVX1 U12432 (.I(n14696), .ZN(n25304));
    INVX1 U12433 (.I(N4013), .ZN(n25305));
    NOR2X1 U12434 (.A1(n17174), .A2(n13981), .ZN(n25306));
    NOR2X1 U12435 (.A1(N4960), .A2(N3379), .ZN(n25307));
    INVX1 U12436 (.I(N3497), .ZN(n25308));
    NANDX1 U12437 (.A1(n18181), .A2(N1485), .ZN(N25309));
    NOR2X1 U12438 (.A1(N1346), .A2(N2338), .ZN(N25310));
    NOR2X1 U12439 (.A1(n19912), .A2(N10955), .ZN(n25311));
    NOR2X1 U12440 (.A1(N6459), .A2(N1924), .ZN(n25312));
    NOR2X1 U12441 (.A1(N207), .A2(n14421), .ZN(N25313));
    INVX1 U12442 (.I(N7015), .ZN(n25314));
    NANDX1 U12443 (.A1(N2682), .A2(N5545), .ZN(n25315));
    NOR2X1 U12444 (.A1(N7984), .A2(N9557), .ZN(N25316));
    NANDX1 U12445 (.A1(N3927), .A2(n18079), .ZN(n25317));
    NANDX1 U12446 (.A1(N8887), .A2(N228), .ZN(N25318));
    NOR2X1 U12447 (.A1(N12383), .A2(N6570), .ZN(N25319));
    NOR2X1 U12448 (.A1(N8409), .A2(N10087), .ZN(n25320));
    NOR2X1 U12449 (.A1(N10746), .A2(N6703), .ZN(n25321));
    INVX1 U12450 (.I(n16242), .ZN(n25322));
    INVX1 U12451 (.I(n20535), .ZN(n25323));
    NANDX1 U12452 (.A1(N8414), .A2(n20742), .ZN(N25324));
    NOR2X1 U12453 (.A1(N5261), .A2(N1068), .ZN(n25325));
    NANDX1 U12454 (.A1(N2484), .A2(N6612), .ZN(n25326));
    NANDX1 U12455 (.A1(N10468), .A2(N10710), .ZN(n25327));
    INVX1 U12456 (.I(n14394), .ZN(n25328));
    INVX1 U12457 (.I(n16977), .ZN(n25329));
    INVX1 U12458 (.I(N2328), .ZN(N25330));
    NANDX1 U12459 (.A1(N8975), .A2(N8897), .ZN(n25331));
    NOR2X1 U12460 (.A1(n17383), .A2(n13525), .ZN(n25332));
    NOR2X1 U12461 (.A1(N6899), .A2(n14770), .ZN(n25333));
    INVX1 U12462 (.I(n17682), .ZN(n25334));
    NANDX1 U12463 (.A1(N8960), .A2(n14617), .ZN(n25335));
    INVX1 U12464 (.I(N3013), .ZN(n25336));
    NOR2X1 U12465 (.A1(N2146), .A2(N4081), .ZN(N25337));
    NANDX1 U12466 (.A1(N4630), .A2(N10692), .ZN(n25338));
    NANDX1 U12467 (.A1(N9639), .A2(n15944), .ZN(N25339));
    NOR2X1 U12468 (.A1(N2802), .A2(N2272), .ZN(N25340));
    NOR2X1 U12469 (.A1(n20624), .A2(n20371), .ZN(n25341));
    INVX1 U12470 (.I(N8368), .ZN(n25342));
    NOR2X1 U12471 (.A1(n18853), .A2(N4520), .ZN(n25343));
    INVX1 U12472 (.I(N8974), .ZN(n25344));
    NOR2X1 U12473 (.A1(N9642), .A2(n13171), .ZN(N25345));
    INVX1 U12474 (.I(N3572), .ZN(n25346));
    NOR2X1 U12475 (.A1(N11570), .A2(N457), .ZN(N25347));
    INVX1 U12476 (.I(N10854), .ZN(n25348));
    NANDX1 U12477 (.A1(N2535), .A2(n15930), .ZN(n25349));
    NANDX1 U12478 (.A1(n13226), .A2(n15300), .ZN(N25350));
    NOR2X1 U12479 (.A1(N2481), .A2(N2916), .ZN(n25351));
    NOR2X1 U12480 (.A1(N4752), .A2(N2051), .ZN(n25352));
    INVX1 U12481 (.I(N3892), .ZN(n25353));
    NOR2X1 U12482 (.A1(n16515), .A2(N6470), .ZN(n25354));
    INVX1 U12483 (.I(n15577), .ZN(n25355));
    NOR2X1 U12484 (.A1(n15772), .A2(N306), .ZN(N25356));
    INVX1 U12485 (.I(N7712), .ZN(n25357));
    NOR2X1 U12486 (.A1(N9098), .A2(N3154), .ZN(N25358));
    NOR2X1 U12487 (.A1(N9554), .A2(N1608), .ZN(N25359));
    NANDX1 U12488 (.A1(N6698), .A2(N4142), .ZN(n25360));
    NOR2X1 U12489 (.A1(N3013), .A2(N11909), .ZN(n25361));
    NOR2X1 U12490 (.A1(N8966), .A2(n14390), .ZN(n25362));
    NOR2X1 U12491 (.A1(n17721), .A2(n13683), .ZN(n25363));
    INVX1 U12492 (.I(N4638), .ZN(n25364));
    INVX1 U12493 (.I(N6218), .ZN(n25365));
    NANDX1 U12494 (.A1(n18586), .A2(N7559), .ZN(n25366));
    INVX1 U12495 (.I(n14470), .ZN(n25367));
    NOR2X1 U12496 (.A1(N10346), .A2(n19996), .ZN(N25368));
    NOR2X1 U12497 (.A1(N7605), .A2(N7863), .ZN(n25369));
    NOR2X1 U12498 (.A1(N10975), .A2(n17416), .ZN(n25370));
    NOR2X1 U12499 (.A1(n19740), .A2(n18656), .ZN(n25371));
    NANDX1 U12500 (.A1(N1975), .A2(N438), .ZN(n25372));
    NOR2X1 U12501 (.A1(n20738), .A2(N9404), .ZN(N25373));
    NANDX1 U12502 (.A1(N10271), .A2(N5894), .ZN(n25374));
    INVX1 U12503 (.I(N1855), .ZN(N25375));
    INVX1 U12504 (.I(N11975), .ZN(N25376));
    INVX1 U12505 (.I(n20767), .ZN(n25377));
    NANDX1 U12506 (.A1(n15630), .A2(N9577), .ZN(n25378));
    NANDX1 U12507 (.A1(N12272), .A2(n19923), .ZN(n25379));
    NOR2X1 U12508 (.A1(N11167), .A2(N839), .ZN(N25380));
    NOR2X1 U12509 (.A1(n13215), .A2(N6355), .ZN(N25381));
    INVX1 U12510 (.I(N11412), .ZN(n25382));
    NANDX1 U12511 (.A1(N7663), .A2(n13750), .ZN(n25383));
    INVX1 U12512 (.I(N2643), .ZN(n25384));
    INVX1 U12513 (.I(N888), .ZN(n25385));
    INVX1 U12514 (.I(n14172), .ZN(n25386));
    NANDX1 U12515 (.A1(N12481), .A2(N8572), .ZN(n25387));
    NANDX1 U12516 (.A1(n17553), .A2(n20546), .ZN(n25388));
    INVX1 U12517 (.I(n17090), .ZN(n25389));
    NOR2X1 U12518 (.A1(N4567), .A2(N5436), .ZN(N25390));
    NANDX1 U12519 (.A1(N11380), .A2(n19900), .ZN(n25391));
    NANDX1 U12520 (.A1(N1316), .A2(n15280), .ZN(n25392));
    INVX1 U12521 (.I(N9072), .ZN(n25393));
    INVX1 U12522 (.I(N9548), .ZN(n25394));
    INVX1 U12523 (.I(N5268), .ZN(n25395));
    NOR2X1 U12524 (.A1(n13002), .A2(N6647), .ZN(N25396));
    NANDX1 U12525 (.A1(n19768), .A2(N7534), .ZN(N25397));
    NOR2X1 U12526 (.A1(N7251), .A2(n13234), .ZN(n25398));
    INVX1 U12527 (.I(n15822), .ZN(N25399));
    NANDX1 U12528 (.A1(N3096), .A2(n15137), .ZN(N25400));
    NOR2X1 U12529 (.A1(n14727), .A2(N12865), .ZN(N25401));
    INVX1 U12530 (.I(n14704), .ZN(n25402));
    NOR2X1 U12531 (.A1(N9898), .A2(n13374), .ZN(n25403));
    NANDX1 U12532 (.A1(N5756), .A2(N1965), .ZN(n25404));
    NOR2X1 U12533 (.A1(n14827), .A2(N2369), .ZN(n25405));
    NOR2X1 U12534 (.A1(N8622), .A2(N2178), .ZN(n25406));
    NANDX1 U12535 (.A1(N393), .A2(N8824), .ZN(N25407));
    NANDX1 U12536 (.A1(n14702), .A2(n16358), .ZN(n25408));
    INVX1 U12537 (.I(N722), .ZN(n25409));
    NANDX1 U12538 (.A1(N2341), .A2(n16543), .ZN(n25410));
    INVX1 U12539 (.I(n21208), .ZN(n25411));
    NANDX1 U12540 (.A1(n17641), .A2(n14704), .ZN(N25412));
    INVX1 U12541 (.I(N10701), .ZN(n25413));
    INVX1 U12542 (.I(n20102), .ZN(n25414));
    NANDX1 U12543 (.A1(n16092), .A2(N7605), .ZN(n25415));
    NOR2X1 U12544 (.A1(n18057), .A2(n15648), .ZN(n25416));
    INVX1 U12545 (.I(n14967), .ZN(n25417));
    INVX1 U12546 (.I(n17655), .ZN(n25418));
    INVX1 U12547 (.I(n14662), .ZN(n25419));
    INVX1 U12548 (.I(N4737), .ZN(N25420));
    INVX1 U12549 (.I(N11519), .ZN(n25421));
    NOR2X1 U12550 (.A1(N588), .A2(N6782), .ZN(n25422));
    NANDX1 U12551 (.A1(n18700), .A2(N2095), .ZN(n25423));
    NOR2X1 U12552 (.A1(n18677), .A2(N1627), .ZN(n25424));
    INVX1 U12553 (.I(N12150), .ZN(N25425));
    NOR2X1 U12554 (.A1(N6877), .A2(n14869), .ZN(N25426));
    NOR2X1 U12555 (.A1(N786), .A2(N4272), .ZN(n25427));
    NANDX1 U12556 (.A1(N451), .A2(n16870), .ZN(n25428));
    NOR2X1 U12557 (.A1(N9484), .A2(N10606), .ZN(N25429));
    INVX1 U12558 (.I(N5908), .ZN(N25430));
    INVX1 U12559 (.I(n19754), .ZN(N25431));
    INVX1 U12560 (.I(N340), .ZN(n25432));
    INVX1 U12561 (.I(N3326), .ZN(n25433));
    NANDX1 U12562 (.A1(n19903), .A2(N10108), .ZN(N25434));
    INVX1 U12563 (.I(n17373), .ZN(n25435));
    NOR2X1 U12564 (.A1(n13049), .A2(n14819), .ZN(n25436));
    NANDX1 U12565 (.A1(N9225), .A2(N281), .ZN(N25437));
    NOR2X1 U12566 (.A1(n16101), .A2(N9691), .ZN(n25438));
    NANDX1 U12567 (.A1(n16886), .A2(n13962), .ZN(N25439));
    INVX1 U12568 (.I(N11878), .ZN(n25440));
    NANDX1 U12569 (.A1(N5810), .A2(N131), .ZN(n25441));
    NANDX1 U12570 (.A1(N10902), .A2(N580), .ZN(n25442));
    NOR2X1 U12571 (.A1(N3967), .A2(n13618), .ZN(N25443));
    NANDX1 U12572 (.A1(N2052), .A2(n16943), .ZN(n25444));
    INVX1 U12573 (.I(N724), .ZN(n25445));
    INVX1 U12574 (.I(n13259), .ZN(n25446));
    NOR2X1 U12575 (.A1(N12563), .A2(N5077), .ZN(n25447));
    NOR2X1 U12576 (.A1(n15475), .A2(n14301), .ZN(N25448));
    NANDX1 U12577 (.A1(N11180), .A2(N3713), .ZN(n25449));
    NOR2X1 U12578 (.A1(N8863), .A2(n20599), .ZN(n25450));
    NOR2X1 U12579 (.A1(n16130), .A2(N11246), .ZN(N25451));
    NANDX1 U12580 (.A1(n16481), .A2(N5919), .ZN(N25452));
    INVX1 U12581 (.I(N6152), .ZN(n25453));
    NANDX1 U12582 (.A1(N567), .A2(N10118), .ZN(n25454));
    INVX1 U12583 (.I(N5799), .ZN(n25455));
    NANDX1 U12584 (.A1(N10370), .A2(N5775), .ZN(N25456));
    NANDX1 U12585 (.A1(N10731), .A2(n13576), .ZN(n25457));
    NOR2X1 U12586 (.A1(n17836), .A2(n18652), .ZN(N25458));
    NANDX1 U12587 (.A1(N12080), .A2(N6265), .ZN(n25459));
    NOR2X1 U12588 (.A1(n17801), .A2(N9977), .ZN(n25460));
    NOR2X1 U12589 (.A1(n21205), .A2(N3887), .ZN(N25461));
    NANDX1 U12590 (.A1(N10646), .A2(n15133), .ZN(n25462));
    INVX1 U12591 (.I(N5896), .ZN(n25463));
    NOR2X1 U12592 (.A1(n17549), .A2(N12047), .ZN(N25464));
    NANDX1 U12593 (.A1(n18115), .A2(n16706), .ZN(n25465));
    NOR2X1 U12594 (.A1(n18455), .A2(n17958), .ZN(n25466));
    INVX1 U12595 (.I(N2999), .ZN(n25467));
    INVX1 U12596 (.I(N9928), .ZN(N25468));
    NANDX1 U12597 (.A1(n13317), .A2(N6533), .ZN(n25469));
    INVX1 U12598 (.I(N7468), .ZN(N25470));
    NOR2X1 U12599 (.A1(N3886), .A2(N8125), .ZN(n25471));
    INVX1 U12600 (.I(n13862), .ZN(N25472));
    INVX1 U12601 (.I(N4241), .ZN(N25473));
    NANDX1 U12602 (.A1(N12552), .A2(n14886), .ZN(n25474));
    NANDX1 U12603 (.A1(N2883), .A2(n15324), .ZN(n25475));
    NANDX1 U12604 (.A1(n14973), .A2(N682), .ZN(n25476));
    INVX1 U12605 (.I(N11857), .ZN(n25477));
    NOR2X1 U12606 (.A1(N6014), .A2(N3623), .ZN(n25478));
    NOR2X1 U12607 (.A1(N5211), .A2(N1164), .ZN(n25479));
    NOR2X1 U12608 (.A1(N9681), .A2(N12279), .ZN(N25480));
    NANDX1 U12609 (.A1(n16213), .A2(n15358), .ZN(n25481));
    NOR2X1 U12610 (.A1(N2679), .A2(n19243), .ZN(n25482));
    INVX1 U12611 (.I(N6944), .ZN(N25483));
    NOR2X1 U12612 (.A1(n18182), .A2(N11184), .ZN(n25484));
    INVX1 U12613 (.I(N9504), .ZN(n25485));
    NANDX1 U12614 (.A1(n19441), .A2(N6928), .ZN(n25486));
    NANDX1 U12615 (.A1(n14537), .A2(N671), .ZN(n25487));
    NANDX1 U12616 (.A1(N5034), .A2(N7069), .ZN(n25488));
    INVX1 U12617 (.I(N5590), .ZN(N25489));
    NANDX1 U12618 (.A1(N9284), .A2(N5342), .ZN(n25490));
    NANDX1 U12619 (.A1(N11185), .A2(n15022), .ZN(N25491));
    INVX1 U12620 (.I(N10631), .ZN(n25492));
    NANDX1 U12621 (.A1(N7345), .A2(N12085), .ZN(n25493));
    NOR2X1 U12622 (.A1(n21129), .A2(n16206), .ZN(n25494));
    INVX1 U12623 (.I(N857), .ZN(n25495));
    NANDX1 U12624 (.A1(n19894), .A2(n14105), .ZN(n25496));
    NOR2X1 U12625 (.A1(n13817), .A2(N6857), .ZN(n25497));
    NANDX1 U12626 (.A1(N1833), .A2(n15935), .ZN(n25498));
    NANDX1 U12627 (.A1(N11760), .A2(n20969), .ZN(n25499));
    NOR2X1 U12628 (.A1(N12387), .A2(N5328), .ZN(N25500));
    NANDX1 U12629 (.A1(n16212), .A2(N10669), .ZN(N25501));
    NOR2X1 U12630 (.A1(N6166), .A2(n20233), .ZN(n25502));
    INVX1 U12631 (.I(n18687), .ZN(n25503));
    INVX1 U12632 (.I(n20855), .ZN(n25504));
    NANDX1 U12633 (.A1(N4466), .A2(n13322), .ZN(N25505));
    NANDX1 U12634 (.A1(N3363), .A2(n20880), .ZN(N25506));
    NANDX1 U12635 (.A1(n20469), .A2(n17990), .ZN(n25507));
    NOR2X1 U12636 (.A1(n23674), .A2(N4145), .ZN(n25508));
    NOR2X1 U12637 (.A1(N4524), .A2(N11820), .ZN(n25509));
    NANDX1 U12638 (.A1(N788), .A2(n14503), .ZN(n25510));
    NANDX1 U12639 (.A1(n14513), .A2(N1192), .ZN(n25511));
    NANDX1 U12640 (.A1(N7996), .A2(n13386), .ZN(N25512));
    NANDX1 U12641 (.A1(n13894), .A2(N509), .ZN(n25513));
    NOR2X1 U12642 (.A1(N7078), .A2(n21058), .ZN(N25514));
    INVX1 U12643 (.I(n16816), .ZN(n25515));
    NOR2X1 U12644 (.A1(N3570), .A2(N2237), .ZN(n25516));
    INVX1 U12645 (.I(n24449), .ZN(n25517));
    NANDX1 U12646 (.A1(N12620), .A2(N5704), .ZN(n25518));
    INVX1 U12647 (.I(N10791), .ZN(n25519));
    NANDX1 U12648 (.A1(n19783), .A2(N4083), .ZN(N25520));
    NOR2X1 U12649 (.A1(n19069), .A2(N4870), .ZN(N25521));
    INVX1 U12650 (.I(N11971), .ZN(n25522));
    INVX1 U12651 (.I(N627), .ZN(N25523));
    NANDX1 U12652 (.A1(n16146), .A2(n14012), .ZN(n25524));
    NOR2X1 U12653 (.A1(n18807), .A2(N3289), .ZN(n25525));
    NOR2X1 U12654 (.A1(N382), .A2(n13114), .ZN(n25526));
    NOR2X1 U12655 (.A1(N5965), .A2(N1903), .ZN(N25527));
    NANDX1 U12656 (.A1(n22471), .A2(n19556), .ZN(n25528));
    NANDX1 U12657 (.A1(N7304), .A2(n20944), .ZN(n25529));
    INVX1 U12658 (.I(N3556), .ZN(N25530));
    NANDX1 U12659 (.A1(n22967), .A2(n23338), .ZN(n25531));
    INVX1 U12660 (.I(N7899), .ZN(n25532));
    INVX1 U12661 (.I(N3952), .ZN(n25533));
    INVX1 U12662 (.I(N3372), .ZN(n25534));
    NOR2X1 U12663 (.A1(n22230), .A2(n19169), .ZN(N25535));
    INVX1 U12664 (.I(n25010), .ZN(n25536));
    NOR2X1 U12665 (.A1(N10319), .A2(N2796), .ZN(n25537));
    NOR2X1 U12666 (.A1(n24970), .A2(n15909), .ZN(N25538));
    NOR2X1 U12667 (.A1(n19702), .A2(N6580), .ZN(n25539));
    NANDX1 U12668 (.A1(n16670), .A2(N633), .ZN(N25540));
    NOR2X1 U12669 (.A1(N12742), .A2(n21576), .ZN(N25541));
    INVX1 U12670 (.I(n16297), .ZN(N25542));
    NOR2X1 U12671 (.A1(n18747), .A2(N2900), .ZN(N25543));
    NOR2X1 U12672 (.A1(n15414), .A2(N8571), .ZN(n25544));
    NANDX1 U12673 (.A1(N11515), .A2(N11942), .ZN(N25545));
    NANDX1 U12674 (.A1(n22513), .A2(n19878), .ZN(n25546));
    NANDX1 U12675 (.A1(n22020), .A2(N4759), .ZN(n25547));
    NOR2X1 U12676 (.A1(n13583), .A2(N12486), .ZN(n25548));
    NANDX1 U12677 (.A1(n18259), .A2(n22075), .ZN(N25549));
    NOR2X1 U12678 (.A1(n24838), .A2(N11592), .ZN(n25550));
    INVX1 U12679 (.I(n14239), .ZN(n25551));
    INVX1 U12680 (.I(N11688), .ZN(N25552));
    NANDX1 U12681 (.A1(N4304), .A2(n16752), .ZN(n25553));
    NANDX1 U12682 (.A1(n23051), .A2(n19651), .ZN(N25554));
    NOR2X1 U12683 (.A1(N1730), .A2(N2719), .ZN(n25555));
    INVX1 U12684 (.I(N2012), .ZN(N25556));
    NOR2X1 U12685 (.A1(N966), .A2(n24524), .ZN(n25557));
    INVX1 U12686 (.I(N1722), .ZN(N25558));
    INVX1 U12687 (.I(n16831), .ZN(N25559));
    NOR2X1 U12688 (.A1(N12159), .A2(N3815), .ZN(N25560));
    INVX1 U12689 (.I(n19186), .ZN(n25561));
    NANDX1 U12690 (.A1(N8653), .A2(n18521), .ZN(n25562));
    NOR2X1 U12691 (.A1(N7599), .A2(N7257), .ZN(n25563));
    NOR2X1 U12692 (.A1(N8054), .A2(N6337), .ZN(n25564));
    NOR2X1 U12693 (.A1(n24805), .A2(N10759), .ZN(n25565));
    NANDX1 U12694 (.A1(N7721), .A2(N5336), .ZN(n25566));
    NOR2X1 U12695 (.A1(n24709), .A2(n22559), .ZN(n25567));
    NOR2X1 U12696 (.A1(N2634), .A2(n23524), .ZN(n25568));
    NANDX1 U12697 (.A1(n14706), .A2(n25245), .ZN(n25569));
    NOR2X1 U12698 (.A1(N6034), .A2(n15577), .ZN(n25570));
    NANDX1 U12699 (.A1(n24118), .A2(n16451), .ZN(n25571));
    INVX1 U12700 (.I(N2040), .ZN(n25572));
    NOR2X1 U12701 (.A1(N6163), .A2(N5823), .ZN(n25573));
    INVX1 U12702 (.I(n13419), .ZN(n25574));
    INVX1 U12703 (.I(N4020), .ZN(N25575));
    NOR2X1 U12704 (.A1(n20469), .A2(n17592), .ZN(N25576));
    INVX1 U12705 (.I(n23394), .ZN(N25577));
    NOR2X1 U12706 (.A1(n24617), .A2(N2547), .ZN(N25578));
    NANDX1 U12707 (.A1(n21673), .A2(n23483), .ZN(n25579));
    INVX1 U12708 (.I(N8462), .ZN(n25580));
    NANDX1 U12709 (.A1(n19392), .A2(N8205), .ZN(n25581));
    NANDX1 U12710 (.A1(n14193), .A2(n23781), .ZN(n25582));
    INVX1 U12711 (.I(N12809), .ZN(n25583));
    NOR2X1 U12712 (.A1(n15034), .A2(N3616), .ZN(n25584));
    NANDX1 U12713 (.A1(n21196), .A2(N9439), .ZN(N25585));
    NOR2X1 U12714 (.A1(n23383), .A2(N2065), .ZN(n25586));
    NOR2X1 U12715 (.A1(N6403), .A2(N11301), .ZN(N25587));
    INVX1 U12716 (.I(n14452), .ZN(n25588));
    NANDX1 U12717 (.A1(N12288), .A2(N2335), .ZN(N25589));
    NANDX1 U12718 (.A1(N71), .A2(n24007), .ZN(n25590));
    NANDX1 U12719 (.A1(N4757), .A2(N6967), .ZN(n25591));
    INVX1 U12720 (.I(n24148), .ZN(n25592));
    NOR2X1 U12721 (.A1(n16162), .A2(N12839), .ZN(n25593));
    NANDX1 U12722 (.A1(N6820), .A2(n14415), .ZN(n25594));
    NOR2X1 U12723 (.A1(N10621), .A2(N6798), .ZN(N25595));
    NANDX1 U12724 (.A1(n20585), .A2(n16236), .ZN(N25596));
    NOR2X1 U12725 (.A1(n18465), .A2(N7069), .ZN(n25597));
    NANDX1 U12726 (.A1(n13635), .A2(N7137), .ZN(n25598));
    NOR2X1 U12727 (.A1(N2585), .A2(N5097), .ZN(N25599));
    NOR2X1 U12728 (.A1(N4919), .A2(n19873), .ZN(n25600));
    NANDX1 U12729 (.A1(n17693), .A2(N7127), .ZN(n25601));
    NANDX1 U12730 (.A1(n13427), .A2(N12319), .ZN(n25602));
    NANDX1 U12731 (.A1(N6133), .A2(n17248), .ZN(n25603));
    INVX1 U12732 (.I(N11388), .ZN(n25604));
    NANDX1 U12733 (.A1(n22437), .A2(n20139), .ZN(n25605));
    NOR2X1 U12734 (.A1(N3732), .A2(n23792), .ZN(N25606));
    INVX1 U12735 (.I(N8736), .ZN(n25607));
    NANDX1 U12736 (.A1(N11499), .A2(N4572), .ZN(n25608));
    INVX1 U12737 (.I(n13902), .ZN(N25609));
    NOR2X1 U12738 (.A1(N6574), .A2(n16486), .ZN(N25610));
    NANDX1 U12739 (.A1(n20749), .A2(N10172), .ZN(N25611));
    INVX1 U12740 (.I(n23763), .ZN(N25612));
    NANDX1 U12741 (.A1(N7070), .A2(N6032), .ZN(n25613));
    NANDX1 U12742 (.A1(N8156), .A2(N1216), .ZN(n25614));
    NOR2X1 U12743 (.A1(n25403), .A2(N9238), .ZN(n25615));
    INVX1 U12744 (.I(N12735), .ZN(N25616));
    NOR2X1 U12745 (.A1(n19750), .A2(N10687), .ZN(N25617));
    NANDX1 U12746 (.A1(N6808), .A2(N3722), .ZN(N25618));
    NANDX1 U12747 (.A1(N10851), .A2(N3988), .ZN(n25619));
    NOR2X1 U12748 (.A1(N4304), .A2(n17889), .ZN(N25620));
    INVX1 U12749 (.I(N10877), .ZN(n25621));
    NOR2X1 U12750 (.A1(N6793), .A2(N6124), .ZN(N25622));
    NANDX1 U12751 (.A1(N6735), .A2(N4384), .ZN(N25623));
    NANDX1 U12752 (.A1(N2572), .A2(n24685), .ZN(n25624));
    NOR2X1 U12753 (.A1(N10727), .A2(N398), .ZN(n25625));
    NANDX1 U12754 (.A1(n24897), .A2(N9635), .ZN(n25626));
    INVX1 U12755 (.I(N12129), .ZN(n25627));
    NANDX1 U12756 (.A1(n25352), .A2(n22816), .ZN(N25628));
    INVX1 U12757 (.I(N6657), .ZN(N25629));
    NOR2X1 U12758 (.A1(n24920), .A2(N6276), .ZN(n25630));
    INVX1 U12759 (.I(N163), .ZN(n25631));
    INVX1 U12760 (.I(N11679), .ZN(n25632));
    NOR2X1 U12761 (.A1(n21456), .A2(N9318), .ZN(n25633));
    NANDX1 U12762 (.A1(n16347), .A2(N5897), .ZN(N25634));
    NOR2X1 U12763 (.A1(N9498), .A2(n19107), .ZN(n25635));
    NOR2X1 U12764 (.A1(N8681), .A2(N139), .ZN(n25636));
    INVX1 U12765 (.I(n23348), .ZN(N25637));
    INVX1 U12766 (.I(n19408), .ZN(n25638));
    NANDX1 U12767 (.A1(N499), .A2(N6034), .ZN(n25639));
    INVX1 U12768 (.I(n14619), .ZN(n25640));
    NANDX1 U12769 (.A1(N4066), .A2(N10043), .ZN(n25641));
    NANDX1 U12770 (.A1(n17754), .A2(N5086), .ZN(n25642));
    NOR2X1 U12771 (.A1(N6684), .A2(n15665), .ZN(N25643));
    NOR2X1 U12772 (.A1(n22336), .A2(N386), .ZN(n25644));
    NANDX1 U12773 (.A1(n19278), .A2(N5500), .ZN(N25645));
    NOR2X1 U12774 (.A1(N11722), .A2(n14997), .ZN(N25646));
    NOR2X1 U12775 (.A1(N6738), .A2(N12445), .ZN(N25647));
    INVX1 U12776 (.I(N1249), .ZN(N25648));
    NOR2X1 U12777 (.A1(N8545), .A2(n20656), .ZN(n25649));
    NANDX1 U12778 (.A1(N9043), .A2(n15457), .ZN(n25650));
    NANDX1 U12779 (.A1(N12429), .A2(n18804), .ZN(n25651));
    INVX1 U12780 (.I(N11240), .ZN(N25652));
    INVX1 U12781 (.I(n17947), .ZN(n25653));
    NANDX1 U12782 (.A1(N1928), .A2(n24630), .ZN(n25654));
    NANDX1 U12783 (.A1(n14814), .A2(n21463), .ZN(N25655));
    NANDX1 U12784 (.A1(n14554), .A2(N4006), .ZN(n25656));
    NOR2X1 U12785 (.A1(N5919), .A2(n15727), .ZN(n25657));
    NOR2X1 U12786 (.A1(N5159), .A2(n22465), .ZN(n25658));
    NANDX1 U12787 (.A1(n18806), .A2(N12481), .ZN(N25659));
    INVX1 U12788 (.I(N1848), .ZN(n25660));
    NANDX1 U12789 (.A1(n22944), .A2(n25161), .ZN(n25661));
    INVX1 U12790 (.I(N4802), .ZN(n25662));
    INVX1 U12791 (.I(n19429), .ZN(n25663));
    NANDX1 U12792 (.A1(N12094), .A2(n20149), .ZN(n25664));
    INVX1 U12793 (.I(N2917), .ZN(n25665));
    NANDX1 U12794 (.A1(N10836), .A2(N12441), .ZN(N25666));
    NOR2X1 U12795 (.A1(n21066), .A2(n22351), .ZN(N25667));
    NANDX1 U12796 (.A1(n25071), .A2(N12257), .ZN(n25668));
    NOR2X1 U12797 (.A1(N4063), .A2(n17160), .ZN(n25669));
    NANDX1 U12798 (.A1(n15295), .A2(n23276), .ZN(N25670));
    NANDX1 U12799 (.A1(N2273), .A2(n14179), .ZN(n25671));
    INVX1 U12800 (.I(n24176), .ZN(n25672));
    NOR2X1 U12801 (.A1(N12400), .A2(n24802), .ZN(N25673));
    NANDX1 U12802 (.A1(n13255), .A2(n18728), .ZN(N25674));
    INVX1 U12803 (.I(n14116), .ZN(N25675));
    INVX1 U12804 (.I(N10660), .ZN(n25676));
    NANDX1 U12805 (.A1(n12986), .A2(n21495), .ZN(n25677));
    INVX1 U12806 (.I(n16179), .ZN(N25678));
    INVX1 U12807 (.I(n15089), .ZN(n25679));
    INVX1 U12808 (.I(n19664), .ZN(n25680));
    INVX1 U12809 (.I(n17817), .ZN(n25681));
    NANDX1 U12810 (.A1(n22041), .A2(n21138), .ZN(N25682));
    NANDX1 U12811 (.A1(n19814), .A2(N6530), .ZN(n25683));
    NANDX1 U12812 (.A1(n22760), .A2(n19271), .ZN(N25684));
    NANDX1 U12813 (.A1(N8878), .A2(n20439), .ZN(n25685));
    NANDX1 U12814 (.A1(N2835), .A2(n22461), .ZN(N25686));
    NANDX1 U12815 (.A1(N1786), .A2(N11074), .ZN(N25687));
    NOR2X1 U12816 (.A1(N12445), .A2(n16874), .ZN(N25688));
    NANDX1 U12817 (.A1(n22707), .A2(n23882), .ZN(n25689));
    NANDX1 U12818 (.A1(N3030), .A2(N2236), .ZN(N25690));
    NANDX1 U12819 (.A1(N11461), .A2(n18348), .ZN(n25691));
    NANDX1 U12820 (.A1(N9685), .A2(n14886), .ZN(n25692));
    NANDX1 U12821 (.A1(n23203), .A2(n23467), .ZN(n25693));
    INVX1 U12822 (.I(N2259), .ZN(n25694));
    INVX1 U12823 (.I(N4305), .ZN(N25695));
    NOR2X1 U12824 (.A1(n18370), .A2(n24743), .ZN(n25696));
    NANDX1 U12825 (.A1(n21205), .A2(n21701), .ZN(n25697));
    INVX1 U12826 (.I(n22990), .ZN(n25698));
    NANDX1 U12827 (.A1(N7753), .A2(n24203), .ZN(n25699));
    NANDX1 U12828 (.A1(n21674), .A2(n21407), .ZN(n25700));
    INVX1 U12829 (.I(N769), .ZN(n25701));
    NANDX1 U12830 (.A1(N2295), .A2(n13788), .ZN(n25702));
    NOR2X1 U12831 (.A1(n20643), .A2(n19121), .ZN(n25703));
    NOR2X1 U12832 (.A1(n24296), .A2(n20090), .ZN(n25704));
    NANDX1 U12833 (.A1(N11029), .A2(N5123), .ZN(N25705));
    INVX1 U12834 (.I(n20521), .ZN(n25706));
    INVX1 U12835 (.I(N6102), .ZN(n25707));
    NOR2X1 U12836 (.A1(N8667), .A2(n17162), .ZN(n25708));
    INVX1 U12837 (.I(n19135), .ZN(N25709));
    NOR2X1 U12838 (.A1(N9616), .A2(N3943), .ZN(n25710));
    NANDX1 U12839 (.A1(n22586), .A2(n16855), .ZN(N25711));
    INVX1 U12840 (.I(n18490), .ZN(n25712));
    NOR2X1 U12841 (.A1(N9243), .A2(n20462), .ZN(N25713));
    NANDX1 U12842 (.A1(n23030), .A2(n19625), .ZN(N25714));
    NANDX1 U12843 (.A1(n16648), .A2(n17239), .ZN(N25715));
    NOR2X1 U12844 (.A1(N3), .A2(N12554), .ZN(n25716));
    NANDX1 U12845 (.A1(N5126), .A2(n24397), .ZN(n25717));
    NOR2X1 U12846 (.A1(n14552), .A2(n19266), .ZN(n25718));
    NANDX1 U12847 (.A1(N11987), .A2(n25195), .ZN(n25719));
    INVX1 U12848 (.I(n19889), .ZN(n25720));
    INVX1 U12849 (.I(N12429), .ZN(n25721));
    NOR2X1 U12850 (.A1(N10471), .A2(N9512), .ZN(N25722));
    NANDX1 U12851 (.A1(n18945), .A2(n16769), .ZN(n25723));
    INVX1 U12852 (.I(N2685), .ZN(N25724));
    NANDX1 U12853 (.A1(N6378), .A2(N212), .ZN(n25725));
    NOR2X1 U12854 (.A1(n23765), .A2(N5628), .ZN(N25726));
    NOR2X1 U12855 (.A1(N3211), .A2(N5630), .ZN(N25727));
    NOR2X1 U12856 (.A1(N7955), .A2(n25025), .ZN(n25728));
    NOR2X1 U12857 (.A1(N7717), .A2(N2843), .ZN(N25729));
    NOR2X1 U12858 (.A1(N9634), .A2(N3597), .ZN(n25730));
    INVX1 U12859 (.I(n23679), .ZN(n25731));
    NANDX1 U12860 (.A1(N9772), .A2(N10605), .ZN(n25732));
    NANDX1 U12861 (.A1(n20242), .A2(N8884), .ZN(N25733));
    INVX1 U12862 (.I(N2453), .ZN(n25734));
    NOR2X1 U12863 (.A1(N1702), .A2(N5137), .ZN(N25735));
    NANDX1 U12864 (.A1(N8079), .A2(n19619), .ZN(N25736));
    INVX1 U12865 (.I(n20611), .ZN(N25737));
    INVX1 U12866 (.I(n21391), .ZN(n25738));
    NOR2X1 U12867 (.A1(N8411), .A2(N9067), .ZN(N25739));
    NOR2X1 U12868 (.A1(N7934), .A2(N9906), .ZN(N25740));
    INVX1 U12869 (.I(n25046), .ZN(n25741));
    NOR2X1 U12870 (.A1(N12391), .A2(N3140), .ZN(N25742));
    NANDX1 U12871 (.A1(n24837), .A2(n15392), .ZN(n25743));
    INVX1 U12872 (.I(n24210), .ZN(N25744));
    NANDX1 U12873 (.A1(n20623), .A2(N7591), .ZN(n25745));
    NOR2X1 U12874 (.A1(n23075), .A2(N7741), .ZN(N25746));
    INVX1 U12875 (.I(n16980), .ZN(n25747));
    INVX1 U12876 (.I(N5357), .ZN(n25748));
    NANDX1 U12877 (.A1(n17921), .A2(n14735), .ZN(N25749));
    NANDX1 U12878 (.A1(n13810), .A2(n13054), .ZN(n25750));
    NANDX1 U12879 (.A1(N11644), .A2(n22364), .ZN(n25751));
    INVX1 U12880 (.I(n21549), .ZN(N25752));
    INVX1 U12881 (.I(N7299), .ZN(n25753));
    NOR2X1 U12882 (.A1(N777), .A2(N10438), .ZN(n25754));
    INVX1 U12883 (.I(N111), .ZN(N25755));
    NOR2X1 U12884 (.A1(n17049), .A2(n24320), .ZN(n25756));
    NANDX1 U12885 (.A1(N937), .A2(n20679), .ZN(N25757));
    NANDX1 U12886 (.A1(n24012), .A2(n17187), .ZN(n25758));
    NANDX1 U12887 (.A1(N4257), .A2(n14342), .ZN(n25759));
    NANDX1 U12888 (.A1(N4120), .A2(N6760), .ZN(n25760));
    NANDX1 U12889 (.A1(N6764), .A2(N9337), .ZN(N25761));
    NANDX1 U12890 (.A1(N6586), .A2(n20980), .ZN(N25762));
    INVX1 U12891 (.I(n14342), .ZN(N25763));
    NANDX1 U12892 (.A1(n15081), .A2(n21640), .ZN(n25764));
    INVX1 U12893 (.I(n15857), .ZN(n25765));
    NOR2X1 U12894 (.A1(n14823), .A2(N4736), .ZN(n25766));
    NOR2X1 U12895 (.A1(n20639), .A2(N3553), .ZN(N25767));
    NANDX1 U12896 (.A1(n21575), .A2(n12999), .ZN(n25768));
    NOR2X1 U12897 (.A1(N8852), .A2(N4684), .ZN(N25769));
    NOR2X1 U12898 (.A1(N1876), .A2(n19025), .ZN(N25770));
    INVX1 U12899 (.I(n20265), .ZN(n25771));
    NOR2X1 U12900 (.A1(N11395), .A2(n15796), .ZN(N25772));
    INVX1 U12901 (.I(n15726), .ZN(n25773));
    NOR2X1 U12902 (.A1(n19366), .A2(N5687), .ZN(n25774));
    INVX1 U12903 (.I(n25160), .ZN(n25775));
    INVX1 U12904 (.I(n21628), .ZN(n25776));
    NOR2X1 U12905 (.A1(n25392), .A2(N2701), .ZN(n25777));
    INVX1 U12906 (.I(N4625), .ZN(n25778));
    NOR2X1 U12907 (.A1(n22041), .A2(n22447), .ZN(N25779));
    NANDX1 U12908 (.A1(N6882), .A2(N9944), .ZN(N25780));
    NANDX1 U12909 (.A1(n15733), .A2(n14627), .ZN(N25781));
    INVX1 U12910 (.I(N6377), .ZN(n25782));
    INVX1 U12911 (.I(N4324), .ZN(n25783));
    NANDX1 U12912 (.A1(n22700), .A2(n15718), .ZN(n25784));
    INVX1 U12913 (.I(N9854), .ZN(n25785));
    INVX1 U12914 (.I(n13814), .ZN(n25786));
    INVX1 U12915 (.I(N396), .ZN(n25787));
    INVX1 U12916 (.I(n17645), .ZN(n25788));
    INVX1 U12917 (.I(N9927), .ZN(n25789));
    INVX1 U12918 (.I(N9819), .ZN(n25790));
    NANDX1 U12919 (.A1(N2590), .A2(N3211), .ZN(N25791));
    NANDX1 U12920 (.A1(n24631), .A2(n14426), .ZN(n25792));
    NOR2X1 U12921 (.A1(n20280), .A2(n24369), .ZN(N25793));
    NANDX1 U12922 (.A1(n24780), .A2(N2261), .ZN(n25794));
    NOR2X1 U12923 (.A1(N5654), .A2(n24679), .ZN(n25795));
    NANDX1 U12924 (.A1(N6793), .A2(N10644), .ZN(n25796));
    INVX1 U12925 (.I(n23727), .ZN(N25797));
    NOR2X1 U12926 (.A1(n16776), .A2(N806), .ZN(N25798));
    NOR2X1 U12927 (.A1(N5939), .A2(n14607), .ZN(n25799));
    NOR2X1 U12928 (.A1(N4636), .A2(n24533), .ZN(n25800));
    INVX1 U12929 (.I(N3223), .ZN(n25801));
    NOR2X1 U12930 (.A1(n23172), .A2(N6433), .ZN(n25802));
    NANDX1 U12931 (.A1(N11068), .A2(n20858), .ZN(n25803));
    INVX1 U12932 (.I(N5845), .ZN(n25804));
    INVX1 U12933 (.I(N2302), .ZN(n25805));
    NANDX1 U12934 (.A1(N10752), .A2(N4328), .ZN(n25806));
    INVX1 U12935 (.I(N9928), .ZN(N25807));
    NANDX1 U12936 (.A1(n17568), .A2(n20572), .ZN(n25808));
    NANDX1 U12937 (.A1(N4560), .A2(n15567), .ZN(N25809));
    NOR2X1 U12938 (.A1(N5365), .A2(N3047), .ZN(n25810));
    NOR2X1 U12939 (.A1(n19971), .A2(N8171), .ZN(N25811));
    NANDX1 U12940 (.A1(N7769), .A2(n14483), .ZN(N25812));
    NOR2X1 U12941 (.A1(N11233), .A2(N12152), .ZN(n25813));
    INVX1 U12942 (.I(N3230), .ZN(n25814));
    INVX1 U12943 (.I(N5903), .ZN(n25815));
    NOR2X1 U12944 (.A1(n17831), .A2(n14394), .ZN(n25816));
    NOR2X1 U12945 (.A1(n22952), .A2(n13914), .ZN(n25817));
    NOR2X1 U12946 (.A1(N8225), .A2(n23841), .ZN(N25818));
    INVX1 U12947 (.I(n14560), .ZN(n25819));
    INVX1 U12948 (.I(n18332), .ZN(n25820));
    INVX1 U12949 (.I(N12012), .ZN(n25821));
    NOR2X1 U12950 (.A1(n13251), .A2(n15058), .ZN(n25822));
    INVX1 U12951 (.I(N7719), .ZN(n25823));
    NOR2X1 U12952 (.A1(N2761), .A2(N4256), .ZN(n25824));
    NANDX1 U12953 (.A1(N6875), .A2(n15488), .ZN(n25825));
    INVX1 U12954 (.I(n17421), .ZN(n25826));
    NOR2X1 U12955 (.A1(n13882), .A2(N12091), .ZN(n25827));
    NOR2X1 U12956 (.A1(N6210), .A2(n15253), .ZN(N25828));
    NOR2X1 U12957 (.A1(N3659), .A2(N3664), .ZN(n25829));
    NOR2X1 U12958 (.A1(N652), .A2(n16272), .ZN(n25830));
    INVX1 U12959 (.I(n15211), .ZN(n25831));
    NANDX1 U12960 (.A1(N12010), .A2(n23098), .ZN(n25832));
    INVX1 U12961 (.I(N6389), .ZN(n25833));
    NOR2X1 U12962 (.A1(N3053), .A2(n22527), .ZN(n25834));
    NANDX1 U12963 (.A1(n15049), .A2(n14055), .ZN(N25835));
    INVX1 U12964 (.I(n16025), .ZN(n25836));
    NANDX1 U12965 (.A1(n15843), .A2(n17920), .ZN(n25837));
    NANDX1 U12966 (.A1(n23327), .A2(n20569), .ZN(N25838));
    NANDX1 U12967 (.A1(N7290), .A2(N1276), .ZN(n25839));
    NANDX1 U12968 (.A1(N6769), .A2(n19204), .ZN(N25840));
    INVX1 U12969 (.I(N3625), .ZN(n25841));
    INVX1 U12970 (.I(N927), .ZN(n25842));
    NANDX1 U12971 (.A1(n23834), .A2(n13644), .ZN(N25843));
    NOR2X1 U12972 (.A1(n21429), .A2(N1638), .ZN(n25844));
    NANDX1 U12973 (.A1(n21042), .A2(N4690), .ZN(n25845));
    NOR2X1 U12974 (.A1(N2872), .A2(n19738), .ZN(n25846));
    INVX1 U12975 (.I(N3227), .ZN(n25847));
    INVX1 U12976 (.I(N2780), .ZN(N25848));
    INVX1 U12977 (.I(N5715), .ZN(n25849));
    NOR2X1 U12978 (.A1(n19931), .A2(N781), .ZN(n25850));
    NOR2X1 U12979 (.A1(N1719), .A2(N2056), .ZN(N25851));
    NANDX1 U12980 (.A1(N8487), .A2(n21260), .ZN(n25852));
    NOR2X1 U12981 (.A1(N879), .A2(N4380), .ZN(N25853));
    NANDX1 U12982 (.A1(n23684), .A2(N2711), .ZN(N25854));
    NOR2X1 U12983 (.A1(N7493), .A2(n12907), .ZN(N25855));
    INVX1 U12984 (.I(N729), .ZN(n25856));
    NOR2X1 U12985 (.A1(n24989), .A2(n16492), .ZN(n25857));
    INVX1 U12986 (.I(N7992), .ZN(n25858));
    INVX1 U12987 (.I(N3313), .ZN(N25859));
    NOR2X1 U12988 (.A1(N12354), .A2(N11149), .ZN(n25860));
    NANDX1 U12989 (.A1(n19787), .A2(n19848), .ZN(N25861));
    NANDX1 U12990 (.A1(N4191), .A2(N10334), .ZN(n25862));
    NOR2X1 U12991 (.A1(N9358), .A2(N7588), .ZN(n25863));
    NANDX1 U12992 (.A1(n24682), .A2(N8466), .ZN(n25864));
    INVX1 U12993 (.I(n15430), .ZN(n25865));
    NOR2X1 U12994 (.A1(n21455), .A2(n22859), .ZN(n25866));
    NOR2X1 U12995 (.A1(N8860), .A2(n17656), .ZN(N25867));
    NOR2X1 U12996 (.A1(n17306), .A2(N5910), .ZN(n25868));
    INVX1 U12997 (.I(n17391), .ZN(n25869));
    INVX1 U12998 (.I(n18469), .ZN(N25870));
    INVX1 U12999 (.I(n20920), .ZN(n25871));
    NOR2X1 U13000 (.A1(n20620), .A2(n22422), .ZN(n25872));
    NOR2X1 U13001 (.A1(N3733), .A2(N10434), .ZN(n25873));
    NANDX1 U13002 (.A1(n14066), .A2(n14771), .ZN(n25874));
    NANDX1 U13003 (.A1(n21653), .A2(N3634), .ZN(n25875));
    NOR2X1 U13004 (.A1(n18886), .A2(n22378), .ZN(n25876));
    NANDX1 U13005 (.A1(n14301), .A2(N7098), .ZN(n25877));
    INVX1 U13006 (.I(n17208), .ZN(n25878));
    INVX1 U13007 (.I(n23347), .ZN(n25879));
    NANDX1 U13008 (.A1(N10798), .A2(N3754), .ZN(n25880));
    NOR2X1 U13009 (.A1(N2687), .A2(n17654), .ZN(n25881));
    NOR2X1 U13010 (.A1(N12157), .A2(N1840), .ZN(n25882));
    NOR2X1 U13011 (.A1(n21544), .A2(n24261), .ZN(n25883));
    NOR2X1 U13012 (.A1(n14044), .A2(n23462), .ZN(n25884));
    INVX1 U13013 (.I(N2607), .ZN(n25885));
    INVX1 U13014 (.I(n19992), .ZN(n25886));
    INVX1 U13015 (.I(n19401), .ZN(n25887));
    INVX1 U13016 (.I(n20681), .ZN(N25888));
    NOR2X1 U13017 (.A1(n18193), .A2(N9479), .ZN(n25889));
    NANDX1 U13018 (.A1(n23884), .A2(n15454), .ZN(n25890));
    NANDX1 U13019 (.A1(n21728), .A2(n13832), .ZN(n25891));
    NANDX1 U13020 (.A1(n14249), .A2(N6835), .ZN(N25892));
    INVX1 U13021 (.I(n20671), .ZN(n25893));
    INVX1 U13022 (.I(N5772), .ZN(n25894));
    INVX1 U13023 (.I(N1402), .ZN(n25895));
    INVX1 U13024 (.I(N10036), .ZN(N25896));
    INVX1 U13025 (.I(N4625), .ZN(n25897));
    NANDX1 U13026 (.A1(n13405), .A2(n21502), .ZN(n25898));
    NANDX1 U13027 (.A1(N7894), .A2(n23296), .ZN(n25899));
    NOR2X1 U13028 (.A1(N6520), .A2(n18474), .ZN(n25900));
    NOR2X1 U13029 (.A1(n13481), .A2(n16720), .ZN(n25901));
    INVX1 U13030 (.I(N630), .ZN(n25902));
    NOR2X1 U13031 (.A1(N707), .A2(n22358), .ZN(n25903));
    INVX1 U13032 (.I(n17138), .ZN(n25904));
    NANDX1 U13033 (.A1(n16105), .A2(n21985), .ZN(n25905));
    NANDX1 U13034 (.A1(N11947), .A2(n16524), .ZN(n25906));
    NOR2X1 U13035 (.A1(n13349), .A2(n21375), .ZN(N25907));
    NOR2X1 U13036 (.A1(N11720), .A2(N498), .ZN(N25908));
    INVX1 U13037 (.I(n13892), .ZN(n25909));
    NANDX1 U13038 (.A1(N142), .A2(N10554), .ZN(N25910));
    NOR2X1 U13039 (.A1(n17802), .A2(n17073), .ZN(n25911));
    NOR2X1 U13040 (.A1(N3771), .A2(n19321), .ZN(n25912));
    INVX1 U13041 (.I(n13114), .ZN(N25913));
    NANDX1 U13042 (.A1(N2458), .A2(N2588), .ZN(N25914));
    INVX1 U13043 (.I(n22960), .ZN(n25915));
    NANDX1 U13044 (.A1(N5445), .A2(N2330), .ZN(n25916));
    INVX1 U13045 (.I(N485), .ZN(n25917));
    NANDX1 U13046 (.A1(N10266), .A2(N6801), .ZN(N25918));
    NANDX1 U13047 (.A1(N6139), .A2(N11921), .ZN(n25919));
    NOR2X1 U13048 (.A1(N6636), .A2(n13802), .ZN(n25920));
    NANDX1 U13049 (.A1(n17402), .A2(n13943), .ZN(n25921));
    INVX1 U13050 (.I(n14729), .ZN(n25922));
    NANDX1 U13051 (.A1(n21663), .A2(n19298), .ZN(N25923));
    NANDX1 U13052 (.A1(n15481), .A2(N815), .ZN(n25924));
    NOR2X1 U13053 (.A1(n24199), .A2(N3272), .ZN(n25925));
    NOR2X1 U13054 (.A1(N4270), .A2(n14999), .ZN(n25926));
    NANDX1 U13055 (.A1(N9715), .A2(n17328), .ZN(n25927));
    NANDX1 U13056 (.A1(n24469), .A2(n20372), .ZN(N25928));
    NANDX1 U13057 (.A1(N5767), .A2(N11262), .ZN(n25929));
    NOR2X1 U13058 (.A1(N6455), .A2(N2639), .ZN(n25930));
    NANDX1 U13059 (.A1(n20257), .A2(n22178), .ZN(n25931));
    NANDX1 U13060 (.A1(N8697), .A2(N12497), .ZN(n25932));
    NOR2X1 U13061 (.A1(n17977), .A2(n22927), .ZN(n25933));
    NANDX1 U13062 (.A1(n16757), .A2(n12906), .ZN(n25934));
    NOR2X1 U13063 (.A1(N6186), .A2(N370), .ZN(N25935));
    NANDX1 U13064 (.A1(N9434), .A2(N4640), .ZN(N25936));
    NANDX1 U13065 (.A1(N9942), .A2(N3122), .ZN(n25937));
    NOR2X1 U13066 (.A1(N1154), .A2(N2088), .ZN(n25938));
    NANDX1 U13067 (.A1(n16901), .A2(N7854), .ZN(n25939));
    NANDX1 U13068 (.A1(n13285), .A2(N3077), .ZN(n25940));
    INVX1 U13069 (.I(N5071), .ZN(n25941));
    NOR2X1 U13070 (.A1(n17677), .A2(n14259), .ZN(n25942));
    INVX1 U13071 (.I(n18942), .ZN(n25943));
    NANDX1 U13072 (.A1(n13271), .A2(n16366), .ZN(N25944));
    NOR2X1 U13073 (.A1(n18795), .A2(n18039), .ZN(n25945));
    NOR2X1 U13074 (.A1(n24980), .A2(n18409), .ZN(N25946));
    INVX1 U13075 (.I(n23181), .ZN(n25947));
    NOR2X1 U13076 (.A1(n23721), .A2(N7620), .ZN(N25948));
    NANDX1 U13077 (.A1(n21683), .A2(n23043), .ZN(n25949));
    INVX1 U13078 (.I(n14514), .ZN(n25950));
    NANDX1 U13079 (.A1(n13645), .A2(N7375), .ZN(n25951));
    NOR2X1 U13080 (.A1(n16721), .A2(n17145), .ZN(n25952));
    NANDX1 U13081 (.A1(n14551), .A2(n23589), .ZN(n25953));
    INVX1 U13082 (.I(n24116), .ZN(n25954));
    NOR2X1 U13083 (.A1(n14798), .A2(N652), .ZN(n25955));
    INVX1 U13084 (.I(N11486), .ZN(n25956));
    NANDX1 U13085 (.A1(N3466), .A2(n18505), .ZN(n25957));
    NOR2X1 U13086 (.A1(n21874), .A2(n13624), .ZN(N25958));
    NANDX1 U13087 (.A1(n22457), .A2(N610), .ZN(N25959));
    NOR2X1 U13088 (.A1(N11891), .A2(n22292), .ZN(N25960));
    NANDX1 U13089 (.A1(n17682), .A2(N72), .ZN(n25961));
    INVX1 U13090 (.I(N5825), .ZN(n25962));
    NANDX1 U13091 (.A1(n19001), .A2(N11313), .ZN(n25963));
    INVX1 U13092 (.I(N3830), .ZN(n25964));
    NOR2X1 U13093 (.A1(N11445), .A2(N2918), .ZN(n25965));
    NOR2X1 U13094 (.A1(n17240), .A2(n17715), .ZN(n25966));
    INVX1 U13095 (.I(N2667), .ZN(n25967));
    NOR2X1 U13096 (.A1(n22110), .A2(N6133), .ZN(N25968));
    INVX1 U13097 (.I(N4300), .ZN(n25969));
    INVX1 U13098 (.I(n24594), .ZN(N25970));
    NANDX1 U13099 (.A1(n13729), .A2(n25203), .ZN(N25971));
    INVX1 U13100 (.I(n14387), .ZN(N25972));
    NOR2X1 U13101 (.A1(n13763), .A2(N6567), .ZN(n25973));
    INVX1 U13102 (.I(n16270), .ZN(n25974));
    NOR2X1 U13103 (.A1(n21315), .A2(n24038), .ZN(n25975));
    NOR2X1 U13104 (.A1(n23441), .A2(n16636), .ZN(N25976));
    NANDX1 U13105 (.A1(n23653), .A2(n19553), .ZN(n25977));
    INVX1 U13106 (.I(N4158), .ZN(N25978));
    NANDX1 U13107 (.A1(n17508), .A2(N6825), .ZN(n25979));
    NANDX1 U13108 (.A1(n14115), .A2(n12957), .ZN(n25980));
    NOR2X1 U13109 (.A1(N7182), .A2(n18498), .ZN(n25981));
    INVX1 U13110 (.I(N5619), .ZN(n25982));
    NOR2X1 U13111 (.A1(n17030), .A2(n20084), .ZN(n25983));
    INVX1 U13112 (.I(n16558), .ZN(n25984));
    INVX1 U13113 (.I(n16445), .ZN(n25985));
    NANDX1 U13114 (.A1(n13382), .A2(n17603), .ZN(n25986));
    INVX1 U13115 (.I(N685), .ZN(n25987));
    INVX1 U13116 (.I(n24177), .ZN(N25988));
    INVX1 U13117 (.I(N6171), .ZN(n25989));
    INVX1 U13118 (.I(N138), .ZN(n25990));
    INVX1 U13119 (.I(N983), .ZN(n25991));
    NANDX1 U13120 (.A1(N1787), .A2(N7807), .ZN(n25992));
    INVX1 U13121 (.I(n15902), .ZN(n25993));
    INVX1 U13122 (.I(n23138), .ZN(n25994));
    NOR2X1 U13123 (.A1(N2526), .A2(n14965), .ZN(n25995));
    INVX1 U13124 (.I(n23520), .ZN(n25996));
    INVX1 U13125 (.I(N12051), .ZN(n25997));
    INVX1 U13126 (.I(N11817), .ZN(n25998));
    NOR2X1 U13127 (.A1(n24340), .A2(n16741), .ZN(n25999));
    NANDX1 U13128 (.A1(N5208), .A2(n17477), .ZN(N26000));
    NANDX1 U13129 (.A1(N9778), .A2(n16152), .ZN(n26001));
    NANDX1 U13130 (.A1(N4716), .A2(N1744), .ZN(N26002));
    NANDX1 U13131 (.A1(n14498), .A2(N2726), .ZN(n26003));
    INVX1 U13132 (.I(n16284), .ZN(n26004));
    INVX1 U13133 (.I(N12559), .ZN(N26005));
    NOR2X1 U13134 (.A1(n23100), .A2(n24464), .ZN(N26006));
    INVX1 U13135 (.I(n14394), .ZN(n26007));
    INVX1 U13136 (.I(n24771), .ZN(n26008));
    NANDX1 U13137 (.A1(N9185), .A2(N87), .ZN(N26009));
    NANDX1 U13138 (.A1(N9769), .A2(n23518), .ZN(N26010));
    INVX1 U13139 (.I(N1007), .ZN(n26011));
    NANDX1 U13140 (.A1(N1886), .A2(N7252), .ZN(n26012));
    NOR2X1 U13141 (.A1(N431), .A2(n23403), .ZN(n26013));
    NANDX1 U13142 (.A1(N5147), .A2(n13914), .ZN(n26014));
    INVX1 U13143 (.I(N8412), .ZN(n26015));
    NANDX1 U13144 (.A1(N6084), .A2(n13463), .ZN(n26016));
    NOR2X1 U13145 (.A1(N7410), .A2(N8914), .ZN(n26017));
    NANDX1 U13146 (.A1(N6372), .A2(N4983), .ZN(n26018));
    INVX1 U13147 (.I(n20297), .ZN(n26019));
    INVX1 U13148 (.I(n20914), .ZN(N26020));
    NOR2X1 U13149 (.A1(n18607), .A2(N4485), .ZN(n26021));
    NOR2X1 U13150 (.A1(n16622), .A2(n15433), .ZN(n26022));
    NOR2X1 U13151 (.A1(N446), .A2(N6086), .ZN(N26023));
    NANDX1 U13152 (.A1(n24805), .A2(N6516), .ZN(N26024));
    NANDX1 U13153 (.A1(N5011), .A2(N430), .ZN(n26025));
    INVX1 U13154 (.I(n17706), .ZN(n26026));
    NANDX1 U13155 (.A1(n19800), .A2(n23790), .ZN(n26027));
    NANDX1 U13156 (.A1(n13275), .A2(n19967), .ZN(N26028));
    NANDX1 U13157 (.A1(n18617), .A2(N836), .ZN(N26029));
    NANDX1 U13158 (.A1(N12850), .A2(N9901), .ZN(n26030));
    NOR2X1 U13159 (.A1(N8261), .A2(n16918), .ZN(n26031));
    NOR2X1 U13160 (.A1(N1513), .A2(N8201), .ZN(N26032));
    NANDX1 U13161 (.A1(n16945), .A2(n14761), .ZN(n26033));
    NOR2X1 U13162 (.A1(n23030), .A2(N3070), .ZN(N26034));
    INVX1 U13163 (.I(n18313), .ZN(n26035));
    NANDX1 U13164 (.A1(N10004), .A2(N7511), .ZN(n26036));
    NOR2X1 U13165 (.A1(n16478), .A2(N5119), .ZN(n26037));
    NANDX1 U13166 (.A1(n14765), .A2(N4958), .ZN(n26038));
    INVX1 U13167 (.I(n23499), .ZN(N26039));
    NANDX1 U13168 (.A1(n21665), .A2(n24335), .ZN(n26040));
    INVX1 U13169 (.I(N9012), .ZN(n26041));
    NOR2X1 U13170 (.A1(n22964), .A2(N6040), .ZN(N26042));
    NOR2X1 U13171 (.A1(n22820), .A2(N7552), .ZN(n26043));
    NANDX1 U13172 (.A1(n13796), .A2(n24496), .ZN(n26044));
    NANDX1 U13173 (.A1(n19487), .A2(N10791), .ZN(n26045));
    NOR2X1 U13174 (.A1(n24480), .A2(n17872), .ZN(n26046));
    NANDX1 U13175 (.A1(n23252), .A2(n25382), .ZN(n26047));
    NANDX1 U13176 (.A1(n14227), .A2(n19268), .ZN(N26048));
    INVX1 U13177 (.I(n17759), .ZN(n26049));
    INVX1 U13178 (.I(N6795), .ZN(N26050));
    NOR2X1 U13179 (.A1(n15471), .A2(N2957), .ZN(n26051));
    NANDX1 U13180 (.A1(N6181), .A2(N737), .ZN(N26052));
    INVX1 U13181 (.I(N3642), .ZN(N26053));
    NOR2X1 U13182 (.A1(N4040), .A2(n15230), .ZN(n26054));
    INVX1 U13183 (.I(n15426), .ZN(N26055));
    NOR2X1 U13184 (.A1(N2089), .A2(n16070), .ZN(N26056));
    INVX1 U13185 (.I(n12880), .ZN(n26057));
    NANDX1 U13186 (.A1(n25024), .A2(N5249), .ZN(N26058));
    INVX1 U13187 (.I(n22773), .ZN(n26059));
    INVX1 U13188 (.I(N4282), .ZN(n26060));
    INVX1 U13189 (.I(N1931), .ZN(n26061));
    NOR2X1 U13190 (.A1(N6791), .A2(n14924), .ZN(N26062));
    INVX1 U13191 (.I(N11314), .ZN(n26063));
    INVX1 U13192 (.I(N6546), .ZN(n26064));
    NANDX1 U13193 (.A1(n25343), .A2(N7282), .ZN(N26065));
    INVX1 U13194 (.I(n17752), .ZN(n26066));
    NOR2X1 U13195 (.A1(n22600), .A2(N7479), .ZN(n26067));
    NOR2X1 U13196 (.A1(N12523), .A2(n25271), .ZN(n26068));
    NOR2X1 U13197 (.A1(N3090), .A2(N11545), .ZN(n26069));
    INVX1 U13198 (.I(N11641), .ZN(n26070));
    NANDX1 U13199 (.A1(N634), .A2(N1951), .ZN(n26071));
    NOR2X1 U13200 (.A1(N8799), .A2(n20503), .ZN(N26072));
    NANDX1 U13201 (.A1(N10730), .A2(n17298), .ZN(N26073));
    INVX1 U13202 (.I(n14421), .ZN(n26074));
    INVX1 U13203 (.I(n18511), .ZN(n26075));
    NOR2X1 U13204 (.A1(N1930), .A2(N10715), .ZN(N26076));
    INVX1 U13205 (.I(N9212), .ZN(N26077));
    NOR2X1 U13206 (.A1(N3209), .A2(N12037), .ZN(N26078));
    INVX1 U13207 (.I(N10687), .ZN(N26079));
    NOR2X1 U13208 (.A1(n16431), .A2(n24726), .ZN(N26080));
    NANDX1 U13209 (.A1(N8288), .A2(N10768), .ZN(n26081));
    NOR2X1 U13210 (.A1(n19928), .A2(N10602), .ZN(n26082));
    NANDX1 U13211 (.A1(N10647), .A2(N7707), .ZN(n26083));
    NOR2X1 U13212 (.A1(N5647), .A2(N8114), .ZN(n26084));
    NOR2X1 U13213 (.A1(n22944), .A2(n15311), .ZN(n26085));
    NANDX1 U13214 (.A1(n18328), .A2(n22590), .ZN(n26086));
    NOR2X1 U13215 (.A1(N9025), .A2(N7802), .ZN(n26087));
    INVX1 U13216 (.I(n18236), .ZN(n26088));
    NOR2X1 U13217 (.A1(n15943), .A2(n19040), .ZN(n26089));
    INVX1 U13218 (.I(n15398), .ZN(n26090));
    NANDX1 U13219 (.A1(n20679), .A2(n14621), .ZN(N26091));
    INVX1 U13220 (.I(N3465), .ZN(n26092));
    INVX1 U13221 (.I(n12961), .ZN(n26093));
    NANDX1 U13222 (.A1(n24758), .A2(n20674), .ZN(N26094));
    INVX1 U13223 (.I(N6962), .ZN(n26095));
    NANDX1 U13224 (.A1(N2950), .A2(N3843), .ZN(N26096));
    INVX1 U13225 (.I(n14661), .ZN(N26097));
    INVX1 U13226 (.I(n21389), .ZN(n26098));
    INVX1 U13227 (.I(N5008), .ZN(n26099));
    NOR2X1 U13228 (.A1(N5279), .A2(N12809), .ZN(N26100));
    INVX1 U13229 (.I(N12282), .ZN(n26101));
    INVX1 U13230 (.I(n15108), .ZN(n26102));
    NANDX1 U13231 (.A1(N6167), .A2(n19273), .ZN(N26103));
    NOR2X1 U13232 (.A1(N1343), .A2(N8391), .ZN(N26104));
    INVX1 U13233 (.I(n19077), .ZN(n26105));
    NANDX1 U13234 (.A1(n24921), .A2(N5735), .ZN(N26106));
    NOR2X1 U13235 (.A1(n20093), .A2(n17308), .ZN(n26107));
    NANDX1 U13236 (.A1(n20544), .A2(N9026), .ZN(n26108));
    NOR2X1 U13237 (.A1(n22735), .A2(n23686), .ZN(n26109));
    NANDX1 U13238 (.A1(n18621), .A2(n19940), .ZN(n26110));
    NOR2X1 U13239 (.A1(N5051), .A2(n25218), .ZN(n26111));
    NANDX1 U13240 (.A1(N4215), .A2(N11997), .ZN(N26112));
    NANDX1 U13241 (.A1(N8090), .A2(N6584), .ZN(N26113));
    INVX1 U13242 (.I(N1860), .ZN(n26114));
    NANDX1 U13243 (.A1(n22839), .A2(N10250), .ZN(n26115));
    NANDX1 U13244 (.A1(n16413), .A2(n21564), .ZN(N26116));
    INVX1 U13245 (.I(N10915), .ZN(n26117));
    NOR2X1 U13246 (.A1(n18634), .A2(n16991), .ZN(N26118));
    NANDX1 U13247 (.A1(n13675), .A2(N514), .ZN(n26119));
    NANDX1 U13248 (.A1(n25177), .A2(n12967), .ZN(N26120));
    NOR2X1 U13249 (.A1(n18295), .A2(N7404), .ZN(n26121));
    INVX1 U13250 (.I(n23345), .ZN(n26122));
    INVX1 U13251 (.I(n20527), .ZN(N26123));
    INVX1 U13252 (.I(n22154), .ZN(N26124));
    INVX1 U13253 (.I(n13185), .ZN(n26125));
    NOR2X1 U13254 (.A1(N3310), .A2(n15045), .ZN(n26126));
    NANDX1 U13255 (.A1(N646), .A2(n14062), .ZN(n26127));
    INVX1 U13256 (.I(N5826), .ZN(n26128));
    NANDX1 U13257 (.A1(n21757), .A2(N5509), .ZN(n26129));
    NANDX1 U13258 (.A1(N3656), .A2(n22499), .ZN(n26130));
    NOR2X1 U13259 (.A1(n17330), .A2(n23012), .ZN(N26131));
    NANDX1 U13260 (.A1(n17005), .A2(N10476), .ZN(N26132));
    NOR2X1 U13261 (.A1(n24067), .A2(N6648), .ZN(n26133));
    NOR2X1 U13262 (.A1(N10678), .A2(n16804), .ZN(N26134));
    NANDX1 U13263 (.A1(n15773), .A2(n13455), .ZN(n26135));
    NOR2X1 U13264 (.A1(N3455), .A2(N5458), .ZN(n26136));
    NANDX1 U13265 (.A1(n18499), .A2(N7086), .ZN(N26137));
    NOR2X1 U13266 (.A1(n21329), .A2(n19069), .ZN(N26138));
    INVX1 U13267 (.I(n20219), .ZN(N26139));
    NANDX1 U13268 (.A1(N218), .A2(N237), .ZN(n26140));
    NOR2X1 U13269 (.A1(N11484), .A2(n18684), .ZN(N26141));
    INVX1 U13270 (.I(n23263), .ZN(n26142));
    NANDX1 U13271 (.A1(N5346), .A2(n22506), .ZN(n26143));
    INVX1 U13272 (.I(n18180), .ZN(n26144));
    NOR2X1 U13273 (.A1(n14306), .A2(N3355), .ZN(n26145));
    INVX1 U13274 (.I(N11346), .ZN(N26146));
    INVX1 U13275 (.I(N11445), .ZN(n26147));
    NANDX1 U13276 (.A1(N11350), .A2(n16902), .ZN(n26148));
    INVX1 U13277 (.I(n18616), .ZN(n26149));
    NOR2X1 U13278 (.A1(n21363), .A2(n14442), .ZN(n26150));
    NOR2X1 U13279 (.A1(N4840), .A2(n23429), .ZN(n26151));
    NOR2X1 U13280 (.A1(n19327), .A2(n23665), .ZN(N26152));
    NANDX1 U13281 (.A1(N5308), .A2(N5615), .ZN(N26153));
    NOR2X1 U13282 (.A1(N3068), .A2(n14808), .ZN(N26154));
    INVX1 U13283 (.I(N72), .ZN(n26155));
    NOR2X1 U13284 (.A1(n18792), .A2(n17992), .ZN(n26156));
    INVX1 U13285 (.I(N10914), .ZN(n26157));
    NOR2X1 U13286 (.A1(N4781), .A2(n18809), .ZN(n26158));
    NANDX1 U13287 (.A1(N12287), .A2(N4656), .ZN(n26159));
    INVX1 U13288 (.I(n19264), .ZN(n26160));
    NANDX1 U13289 (.A1(N6079), .A2(N3893), .ZN(N26161));
    INVX1 U13290 (.I(N12401), .ZN(N26162));
    NANDX1 U13291 (.A1(N10137), .A2(N8543), .ZN(N26163));
    NANDX1 U13292 (.A1(n22569), .A2(N1198), .ZN(n26164));
    NANDX1 U13293 (.A1(N2681), .A2(N7697), .ZN(n26165));
    NOR2X1 U13294 (.A1(N6256), .A2(N8308), .ZN(N26166));
    NANDX1 U13295 (.A1(n22120), .A2(N1597), .ZN(n26167));
    INVX1 U13296 (.I(N1285), .ZN(n26168));
    NOR2X1 U13297 (.A1(N11280), .A2(N6065), .ZN(n26169));
    NOR2X1 U13298 (.A1(n13204), .A2(n18352), .ZN(N26170));
    NOR2X1 U13299 (.A1(n20797), .A2(N881), .ZN(N26171));
    INVX1 U13300 (.I(N1374), .ZN(n26172));
    NOR2X1 U13301 (.A1(n23488), .A2(n13774), .ZN(n26173));
    NANDX1 U13302 (.A1(n22392), .A2(N11084), .ZN(n26174));
    NOR2X1 U13303 (.A1(N8227), .A2(N1049), .ZN(n26175));
    NANDX1 U13304 (.A1(n25177), .A2(N8745), .ZN(n26176));
    INVX1 U13305 (.I(N5931), .ZN(n26177));
    NOR2X1 U13306 (.A1(N929), .A2(N2548), .ZN(n26178));
    NOR2X1 U13307 (.A1(n21729), .A2(n18103), .ZN(n26179));
    NANDX1 U13308 (.A1(n21776), .A2(n24167), .ZN(n26180));
    NANDX1 U13309 (.A1(N9477), .A2(N5784), .ZN(N26181));
    NANDX1 U13310 (.A1(N4771), .A2(N6665), .ZN(n26182));
    NOR2X1 U13311 (.A1(n20414), .A2(N205), .ZN(N26183));
    NANDX1 U13312 (.A1(N8685), .A2(n13709), .ZN(n26184));
    NANDX1 U13313 (.A1(n19768), .A2(n18537), .ZN(n26185));
    NOR2X1 U13314 (.A1(N9585), .A2(n19997), .ZN(n26186));
    INVX1 U13315 (.I(N7097), .ZN(n26187));
    NANDX1 U13316 (.A1(N37), .A2(n12917), .ZN(N26188));
    NANDX1 U13317 (.A1(n16855), .A2(N9102), .ZN(N26189));
    NANDX1 U13318 (.A1(N9455), .A2(N6564), .ZN(n26190));
    NOR2X1 U13319 (.A1(n22389), .A2(n24113), .ZN(N26191));
    INVX1 U13320 (.I(n16941), .ZN(N26192));
    NANDX1 U13321 (.A1(n20635), .A2(N12373), .ZN(n26193));
    NANDX1 U13322 (.A1(N4315), .A2(N12577), .ZN(n26194));
    INVX1 U13323 (.I(n12999), .ZN(n26195));
    INVX1 U13324 (.I(N4716), .ZN(n26196));
    INVX1 U13325 (.I(n22358), .ZN(N26197));
    NANDX1 U13326 (.A1(N5617), .A2(n16852), .ZN(n26198));
    NANDX1 U13327 (.A1(N12713), .A2(N12505), .ZN(N26199));
    NOR2X1 U13328 (.A1(n14398), .A2(n23356), .ZN(N26200));
    INVX1 U13329 (.I(N12267), .ZN(N26201));
    NANDX1 U13330 (.A1(N11405), .A2(n18830), .ZN(n26202));
    INVX1 U13331 (.I(N8291), .ZN(n26203));
    NANDX1 U13332 (.A1(N1681), .A2(n25231), .ZN(N26204));
    INVX1 U13333 (.I(N11083), .ZN(n26205));
    NANDX1 U13334 (.A1(n14064), .A2(n15397), .ZN(N26206));
    NOR2X1 U13335 (.A1(n21341), .A2(N2894), .ZN(n26207));
    NOR2X1 U13336 (.A1(N554), .A2(n13196), .ZN(N26208));
    NOR2X1 U13337 (.A1(n13971), .A2(N7580), .ZN(n26209));
    INVX1 U13338 (.I(N7225), .ZN(n26210));
    NANDX1 U13339 (.A1(n17976), .A2(N3553), .ZN(n26211));
    INVX1 U13340 (.I(N4597), .ZN(n26212));
    NOR2X1 U13341 (.A1(N10221), .A2(n23797), .ZN(n26213));
    NANDX1 U13342 (.A1(N3549), .A2(N9613), .ZN(N26214));
    INVX1 U13343 (.I(n24026), .ZN(N26215));
    NOR2X1 U13344 (.A1(n13694), .A2(n20129), .ZN(n26216));
    NOR2X1 U13345 (.A1(n14562), .A2(n22961), .ZN(n26217));
    NANDX1 U13346 (.A1(N2505), .A2(N7567), .ZN(n26218));
    NANDX1 U13347 (.A1(n19771), .A2(N8121), .ZN(N26219));
    NOR2X1 U13348 (.A1(N8391), .A2(n22091), .ZN(n26220));
    NOR2X1 U13349 (.A1(N2630), .A2(n18083), .ZN(N26221));
    NANDX1 U13350 (.A1(n20605), .A2(N10403), .ZN(n26222));
    NOR2X1 U13351 (.A1(n25201), .A2(N1635), .ZN(N26223));
    NOR2X1 U13352 (.A1(n23495), .A2(N4271), .ZN(n26224));
    NANDX1 U13353 (.A1(n21875), .A2(n18236), .ZN(n26225));
    NOR2X1 U13354 (.A1(N7665), .A2(N6427), .ZN(n26226));
    INVX1 U13355 (.I(n18807), .ZN(N26227));
    INVX1 U13356 (.I(n16669), .ZN(N26228));
    NANDX1 U13357 (.A1(N12261), .A2(n24236), .ZN(n26229));
    INVX1 U13358 (.I(N6529), .ZN(N26230));
    NOR2X1 U13359 (.A1(n18435), .A2(N3687), .ZN(N26231));
    NOR2X1 U13360 (.A1(n20675), .A2(N6316), .ZN(n26232));
    NOR2X1 U13361 (.A1(n17705), .A2(n15688), .ZN(n26233));
    NOR2X1 U13362 (.A1(N1457), .A2(n15386), .ZN(N26234));
    NANDX1 U13363 (.A1(N6661), .A2(N2146), .ZN(N26235));
    NANDX1 U13364 (.A1(n18452), .A2(N12788), .ZN(N26236));
    NOR2X1 U13365 (.A1(N3264), .A2(N9220), .ZN(N26237));
    NOR2X1 U13366 (.A1(n22474), .A2(n16795), .ZN(N26238));
    NANDX1 U13367 (.A1(n13641), .A2(N11136), .ZN(n26239));
    NOR2X1 U13368 (.A1(N1142), .A2(N12446), .ZN(n26240));
    INVX1 U13369 (.I(n22265), .ZN(n26241));
    NOR2X1 U13370 (.A1(n13062), .A2(N3242), .ZN(n26242));
    NOR2X1 U13371 (.A1(n19377), .A2(n16572), .ZN(n26243));
    NANDX1 U13372 (.A1(N9563), .A2(n14803), .ZN(N26244));
    NOR2X1 U13373 (.A1(n13716), .A2(n14668), .ZN(n26245));
    INVX1 U13374 (.I(N4630), .ZN(N26246));
    NANDX1 U13375 (.A1(N11126), .A2(N6185), .ZN(N26247));
    NANDX1 U13376 (.A1(N3157), .A2(n15405), .ZN(n26248));
    NANDX1 U13377 (.A1(N129), .A2(N6697), .ZN(N26249));
    NOR2X1 U13378 (.A1(N2537), .A2(N6600), .ZN(n26250));
    NANDX1 U13379 (.A1(N3678), .A2(n19045), .ZN(N26251));
    NOR2X1 U13380 (.A1(N440), .A2(n13191), .ZN(n26252));
    NANDX1 U13381 (.A1(n17951), .A2(n16779), .ZN(n26253));
    NOR2X1 U13382 (.A1(N9021), .A2(N1337), .ZN(N26254));
    INVX1 U13383 (.I(n23823), .ZN(n26255));
    NOR2X1 U13384 (.A1(N10096), .A2(N1756), .ZN(n26256));
    INVX1 U13385 (.I(N3493), .ZN(n26257));
    NANDX1 U13386 (.A1(N5421), .A2(N9677), .ZN(n26258));
    NOR2X1 U13387 (.A1(N8577), .A2(n25081), .ZN(N26259));
    NANDX1 U13388 (.A1(n22975), .A2(N6275), .ZN(n26260));
    NANDX1 U13389 (.A1(N9), .A2(N1643), .ZN(N26261));
    INVX1 U13390 (.I(N3686), .ZN(n26262));
    NOR2X1 U13391 (.A1(n19094), .A2(n18395), .ZN(n26263));
    NANDX1 U13392 (.A1(N8999), .A2(N10844), .ZN(N26264));
    INVX1 U13393 (.I(N7048), .ZN(n26265));
    NOR2X1 U13394 (.A1(N4025), .A2(N3428), .ZN(n26266));
    NOR2X1 U13395 (.A1(n16877), .A2(n13523), .ZN(n26267));
    NOR2X1 U13396 (.A1(n22404), .A2(n17015), .ZN(n26268));
    INVX1 U13397 (.I(N2322), .ZN(n26269));
    NANDX1 U13398 (.A1(n18447), .A2(N10898), .ZN(n26270));
    NOR2X1 U13399 (.A1(n15363), .A2(N8371), .ZN(n26271));
    INVX1 U13400 (.I(N2404), .ZN(n26272));
    NOR2X1 U13401 (.A1(N11722), .A2(n19151), .ZN(N26273));
    INVX1 U13402 (.I(n21177), .ZN(N26274));
    NOR2X1 U13403 (.A1(n19227), .A2(n18319), .ZN(n26275));
    NANDX1 U13404 (.A1(N4568), .A2(N9776), .ZN(N26276));
    INVX1 U13405 (.I(n13199), .ZN(N26277));
    NOR2X1 U13406 (.A1(n24021), .A2(n20150), .ZN(n26278));
    NANDX1 U13407 (.A1(N12041), .A2(N6392), .ZN(N26279));
    NOR2X1 U13408 (.A1(n17823), .A2(n16230), .ZN(n26280));
    NOR2X1 U13409 (.A1(N7779), .A2(n23444), .ZN(n26281));
    INVX1 U13410 (.I(n22816), .ZN(n26282));
    NANDX1 U13411 (.A1(n15470), .A2(n21664), .ZN(n26283));
    NOR2X1 U13412 (.A1(N12617), .A2(N7883), .ZN(N26284));
    NOR2X1 U13413 (.A1(n13449), .A2(N3557), .ZN(N26285));
    NANDX1 U13414 (.A1(n21443), .A2(N10644), .ZN(N26286));
    NANDX1 U13415 (.A1(n14779), .A2(n20419), .ZN(n26287));
    NANDX1 U13416 (.A1(N2475), .A2(n22986), .ZN(N26288));
    INVX1 U13417 (.I(N11393), .ZN(N26289));
    INVX1 U13418 (.I(n18828), .ZN(n26290));
    INVX1 U13419 (.I(n22041), .ZN(n26291));
    NANDX1 U13420 (.A1(n22781), .A2(n15205), .ZN(n26292));
    NOR2X1 U13421 (.A1(n20722), .A2(n22305), .ZN(n26293));
    NOR2X1 U13422 (.A1(N8523), .A2(N12272), .ZN(n26294));
    NANDX1 U13423 (.A1(n12998), .A2(n24888), .ZN(n26295));
    NANDX1 U13424 (.A1(N11121), .A2(N1602), .ZN(n26296));
    NANDX1 U13425 (.A1(n25023), .A2(n23045), .ZN(n26297));
    NANDX1 U13426 (.A1(N12699), .A2(N1089), .ZN(N26298));
    NANDX1 U13427 (.A1(n20968), .A2(N3563), .ZN(n26299));
    NANDX1 U13428 (.A1(N2253), .A2(n14955), .ZN(n26300));
    INVX1 U13429 (.I(N9848), .ZN(n26301));
    INVX1 U13430 (.I(N1496), .ZN(n26302));
    NOR2X1 U13431 (.A1(n18785), .A2(N5469), .ZN(n26303));
    NOR2X1 U13432 (.A1(N2773), .A2(N2271), .ZN(N26304));
    NOR2X1 U13433 (.A1(N63), .A2(n14542), .ZN(n26305));
    INVX1 U13434 (.I(n13060), .ZN(n26306));
    INVX1 U13435 (.I(N8100), .ZN(n26307));
    NOR2X1 U13436 (.A1(N4297), .A2(N1281), .ZN(n26308));
    NANDX1 U13437 (.A1(n16109), .A2(N5105), .ZN(n26309));
    INVX1 U13438 (.I(n17197), .ZN(n26310));
    INVX1 U13439 (.I(n20633), .ZN(n26311));
    INVX1 U13440 (.I(N6145), .ZN(n26312));
    NANDX1 U13441 (.A1(n24482), .A2(n25372), .ZN(n26313));
    INVX1 U13442 (.I(N9254), .ZN(n26314));
    INVX1 U13443 (.I(N5761), .ZN(n26315));
    INVX1 U13444 (.I(N6833), .ZN(n26316));
    INVX1 U13445 (.I(n19579), .ZN(N26317));
    NANDX1 U13446 (.A1(n15022), .A2(n19641), .ZN(n26318));
    NOR2X1 U13447 (.A1(n22265), .A2(N7199), .ZN(n26319));
    INVX1 U13448 (.I(N4863), .ZN(n26320));
    NANDX1 U13449 (.A1(n22442), .A2(N6143), .ZN(n26321));
    INVX1 U13450 (.I(n13049), .ZN(N26322));
    INVX1 U13451 (.I(n18009), .ZN(n26323));
    INVX1 U13452 (.I(n21168), .ZN(n26324));
    NOR2X1 U13453 (.A1(N3038), .A2(n16080), .ZN(n26325));
    INVX1 U13454 (.I(n16288), .ZN(N26326));
    NANDX1 U13455 (.A1(N6519), .A2(N39), .ZN(n26327));
    INVX1 U13456 (.I(N12280), .ZN(n26328));
    INVX1 U13457 (.I(n12914), .ZN(N26329));
    NOR2X1 U13458 (.A1(N10921), .A2(N10785), .ZN(n26330));
    INVX1 U13459 (.I(n19330), .ZN(n26331));
    INVX1 U13460 (.I(N2352), .ZN(n26332));
    INVX1 U13461 (.I(n15840), .ZN(n26333));
    NOR2X1 U13462 (.A1(N6901), .A2(N1547), .ZN(n26334));
    INVX1 U13463 (.I(n14013), .ZN(n26335));
    NANDX1 U13464 (.A1(n16410), .A2(N6519), .ZN(n26336));
    INVX1 U13465 (.I(N12075), .ZN(N26337));
    NANDX1 U13466 (.A1(n14181), .A2(n16923), .ZN(n26338));
    NOR2X1 U13467 (.A1(n19236), .A2(N7369), .ZN(N26339));
    NANDX1 U13468 (.A1(N8043), .A2(n13450), .ZN(n26340));
    NANDX1 U13469 (.A1(n13655), .A2(n15132), .ZN(n26341));
    NANDX1 U13470 (.A1(n13344), .A2(n14684), .ZN(n26342));
    NOR2X1 U13471 (.A1(N7171), .A2(n15416), .ZN(n26343));
    NANDX1 U13472 (.A1(N8196), .A2(n20023), .ZN(n26344));
    INVX1 U13473 (.I(N3864), .ZN(n26345));
    NANDX1 U13474 (.A1(n23124), .A2(n17876), .ZN(N26346));
    NANDX1 U13475 (.A1(N2799), .A2(n24394), .ZN(N26347));
    NANDX1 U13476 (.A1(N3642), .A2(N7316), .ZN(n26348));
    INVX1 U13477 (.I(n20564), .ZN(N26349));
    NOR2X1 U13478 (.A1(n18487), .A2(N2430), .ZN(n26350));
    NANDX1 U13479 (.A1(N1027), .A2(N4648), .ZN(N26351));
    INVX1 U13480 (.I(n14681), .ZN(n26352));
    NOR2X1 U13481 (.A1(n21843), .A2(n16792), .ZN(N26353));
    INVX1 U13482 (.I(N4738), .ZN(N26354));
    NOR2X1 U13483 (.A1(n24375), .A2(N4254), .ZN(n26355));
    NANDX1 U13484 (.A1(N7663), .A2(n25253), .ZN(n26356));
    INVX1 U13485 (.I(N3729), .ZN(n26357));
    NOR2X1 U13486 (.A1(n17162), .A2(N3158), .ZN(N26358));
    NOR2X1 U13487 (.A1(N4822), .A2(n24962), .ZN(N26359));
    INVX1 U13488 (.I(N12137), .ZN(n26360));
    NANDX1 U13489 (.A1(n13143), .A2(N1663), .ZN(N26361));
    NOR2X1 U13490 (.A1(N4341), .A2(N5420), .ZN(n26362));
    INVX1 U13491 (.I(N8988), .ZN(N26363));
    INVX1 U13492 (.I(n24709), .ZN(n26364));
    NANDX1 U13493 (.A1(n20796), .A2(n15999), .ZN(N26365));
    NOR2X1 U13494 (.A1(n14301), .A2(n14458), .ZN(n26366));
    NOR2X1 U13495 (.A1(N7322), .A2(n21113), .ZN(N26367));
    NOR2X1 U13496 (.A1(N7072), .A2(n20399), .ZN(n26368));
    INVX1 U13497 (.I(n18714), .ZN(N26369));
    NANDX1 U13498 (.A1(n17449), .A2(N7653), .ZN(n26370));
    INVX1 U13499 (.I(N5676), .ZN(n26371));
    NANDX1 U13500 (.A1(n17784), .A2(n18656), .ZN(N26372));
    INVX1 U13501 (.I(N8214), .ZN(n26373));
    NOR2X1 U13502 (.A1(n20753), .A2(n13634), .ZN(N26374));
    NOR2X1 U13503 (.A1(n18508), .A2(N12586), .ZN(N26375));
    NOR2X1 U13504 (.A1(n24809), .A2(n22149), .ZN(n26376));
    NOR2X1 U13505 (.A1(n14567), .A2(n25217), .ZN(n26377));
    NOR2X1 U13506 (.A1(n17467), .A2(N7036), .ZN(N26378));
    INVX1 U13507 (.I(N2527), .ZN(n26379));
    INVX1 U13508 (.I(n18082), .ZN(n26380));
    NANDX1 U13509 (.A1(n21589), .A2(n18908), .ZN(n26381));
    NANDX1 U13510 (.A1(n18009), .A2(n24554), .ZN(n26382));
    NANDX1 U13511 (.A1(N7009), .A2(N5603), .ZN(n26383));
    NANDX1 U13512 (.A1(N12189), .A2(n13817), .ZN(N26384));
    NOR2X1 U13513 (.A1(N7439), .A2(N1948), .ZN(N26385));
    NANDX1 U13514 (.A1(n14714), .A2(N3301), .ZN(N26386));
    NANDX1 U13515 (.A1(n14020), .A2(n14218), .ZN(N26387));
    NANDX1 U13516 (.A1(n17354), .A2(N2700), .ZN(n26388));
    NANDX1 U13517 (.A1(N9318), .A2(N9736), .ZN(n26389));
    NOR2X1 U13518 (.A1(N612), .A2(N12611), .ZN(n26390));
    INVX1 U13519 (.I(n20466), .ZN(n26391));
    NANDX1 U13520 (.A1(n23067), .A2(N6765), .ZN(n26392));
    INVX1 U13521 (.I(N10886), .ZN(n26393));
    NANDX1 U13522 (.A1(N11250), .A2(n16489), .ZN(n26394));
    NOR2X1 U13523 (.A1(n23438), .A2(N4803), .ZN(n26395));
    NANDX1 U13524 (.A1(n19644), .A2(n21020), .ZN(n26396));
    NANDX1 U13525 (.A1(n23125), .A2(n13088), .ZN(N26397));
    NOR2X1 U13526 (.A1(N410), .A2(N1803), .ZN(n26398));
    NANDX1 U13527 (.A1(n17763), .A2(N4503), .ZN(N26399));
    INVX1 U13528 (.I(N1578), .ZN(N26400));
    NOR2X1 U13529 (.A1(N6618), .A2(n16459), .ZN(n26401));
    INVX1 U13530 (.I(N10777), .ZN(N26402));
    NANDX1 U13531 (.A1(N1848), .A2(n22611), .ZN(N26403));
    NANDX1 U13532 (.A1(N6089), .A2(N7995), .ZN(n26404));
    INVX1 U13533 (.I(n17338), .ZN(n26405));
    NANDX1 U13534 (.A1(n15060), .A2(N4041), .ZN(N26406));
    NANDX1 U13535 (.A1(N11710), .A2(N12452), .ZN(n26407));
    NANDX1 U13536 (.A1(n16021), .A2(N10074), .ZN(N26408));
    NOR2X1 U13537 (.A1(n22075), .A2(N10483), .ZN(N26409));
    NOR2X1 U13538 (.A1(N3217), .A2(n17013), .ZN(N26410));
    NANDX1 U13539 (.A1(n23757), .A2(n18590), .ZN(n26411));
    INVX1 U13540 (.I(N4872), .ZN(n26412));
    NOR2X1 U13541 (.A1(N6654), .A2(n15649), .ZN(N26413));
    NOR2X1 U13542 (.A1(n22771), .A2(N1525), .ZN(n26414));
    INVX1 U13543 (.I(N3358), .ZN(n26415));
    INVX1 U13544 (.I(n22381), .ZN(n26416));
    INVX1 U13545 (.I(N11537), .ZN(n26417));
    NOR2X1 U13546 (.A1(N2272), .A2(N4087), .ZN(n26418));
    NOR2X1 U13547 (.A1(n14723), .A2(N6424), .ZN(n26419));
    NOR2X1 U13548 (.A1(n13565), .A2(N10617), .ZN(n26420));
    NANDX1 U13549 (.A1(N12815), .A2(n16612), .ZN(n26421));
    NOR2X1 U13550 (.A1(N4326), .A2(n15877), .ZN(n26422));
    INVX1 U13551 (.I(N11683), .ZN(n26423));
    INVX1 U13552 (.I(N8885), .ZN(n26424));
    INVX1 U13553 (.I(N2336), .ZN(n26425));
    NANDX1 U13554 (.A1(n22770), .A2(n25106), .ZN(n26426));
    INVX1 U13555 (.I(N2724), .ZN(n26427));
    INVX1 U13556 (.I(n13112), .ZN(n26428));
    NOR2X1 U13557 (.A1(n15462), .A2(n24649), .ZN(N26429));
    NOR2X1 U13558 (.A1(n17733), .A2(n17503), .ZN(n26430));
    NOR2X1 U13559 (.A1(n21223), .A2(N12695), .ZN(n26431));
    NOR2X1 U13560 (.A1(n23555), .A2(n23311), .ZN(N26432));
    INVX1 U13561 (.I(N10868), .ZN(n26433));
    NOR2X1 U13562 (.A1(n21839), .A2(N3961), .ZN(N26434));
    NOR2X1 U13563 (.A1(N350), .A2(N4411), .ZN(N26435));
    NOR2X1 U13564 (.A1(n23504), .A2(N3175), .ZN(N26436));
    NANDX1 U13565 (.A1(N71), .A2(N442), .ZN(n26437));
    NOR2X1 U13566 (.A1(N3664), .A2(n17436), .ZN(n26438));
    NANDX1 U13567 (.A1(N5543), .A2(N5805), .ZN(n26439));
    INVX1 U13568 (.I(n18959), .ZN(N26440));
    NOR2X1 U13569 (.A1(N7910), .A2(N10960), .ZN(n26441));
    NOR2X1 U13570 (.A1(N3630), .A2(n23654), .ZN(N26442));
    NANDX1 U13571 (.A1(n15953), .A2(n21462), .ZN(n26443));
    NANDX1 U13572 (.A1(n15588), .A2(n24649), .ZN(n26444));
    NOR2X1 U13573 (.A1(n19548), .A2(N6978), .ZN(n26445));
    NOR2X1 U13574 (.A1(n23958), .A2(n21723), .ZN(N26446));
    NANDX1 U13575 (.A1(n15901), .A2(n13301), .ZN(n26447));
    INVX1 U13576 (.I(N5110), .ZN(n26448));
    NANDX1 U13577 (.A1(N8015), .A2(n22545), .ZN(n26449));
    NOR2X1 U13578 (.A1(n13558), .A2(N2848), .ZN(n26450));
    NOR2X1 U13579 (.A1(N7014), .A2(N11997), .ZN(n26451));
    NOR2X1 U13580 (.A1(n17973), .A2(N3209), .ZN(N26452));
    NOR2X1 U13581 (.A1(N4892), .A2(N4919), .ZN(N26453));
    NOR2X1 U13582 (.A1(n15121), .A2(n22708), .ZN(N26454));
    INVX1 U13583 (.I(N3035), .ZN(n26455));
    INVX1 U13584 (.I(n23806), .ZN(n26456));
    NANDX1 U13585 (.A1(n14573), .A2(N11029), .ZN(n26457));
    NANDX1 U13586 (.A1(N4584), .A2(N1427), .ZN(n26458));
    INVX1 U13587 (.I(n20168), .ZN(n26459));
    NANDX1 U13588 (.A1(n15820), .A2(N2680), .ZN(n26460));
    INVX1 U13589 (.I(N9287), .ZN(N26461));
    NOR2X1 U13590 (.A1(n20696), .A2(n18434), .ZN(n26462));
    INVX1 U13591 (.I(n21460), .ZN(n26463));
    NOR2X1 U13592 (.A1(N4489), .A2(n24668), .ZN(n26464));
    NANDX1 U13593 (.A1(n23651), .A2(N4084), .ZN(n26465));
    INVX1 U13594 (.I(n13269), .ZN(n26466));
    INVX1 U13595 (.I(N12369), .ZN(N26467));
    NOR2X1 U13596 (.A1(N12619), .A2(N10672), .ZN(n26468));
    NANDX1 U13597 (.A1(N1689), .A2(n21701), .ZN(n26469));
    INVX1 U13598 (.I(n20543), .ZN(N26470));
    NOR2X1 U13599 (.A1(n18382), .A2(n15208), .ZN(n26471));
    NANDX1 U13600 (.A1(n22969), .A2(N6655), .ZN(n26472));
    INVX1 U13601 (.I(N6754), .ZN(n26473));
    NOR2X1 U13602 (.A1(N5971), .A2(n13955), .ZN(n26474));
    INVX1 U13603 (.I(N1929), .ZN(N26475));
    NOR2X1 U13604 (.A1(N2664), .A2(n15364), .ZN(n26476));
    NANDX1 U13605 (.A1(n15082), .A2(n19448), .ZN(N26477));
    NOR2X1 U13606 (.A1(N2849), .A2(N9504), .ZN(N26478));
    NOR2X1 U13607 (.A1(N7920), .A2(N10891), .ZN(n26479));
    NANDX1 U13608 (.A1(n23002), .A2(N1347), .ZN(N26480));
    INVX1 U13609 (.I(N7582), .ZN(n26481));
    INVX1 U13610 (.I(N962), .ZN(n26482));
    NOR2X1 U13611 (.A1(N362), .A2(n19392), .ZN(N26483));
    INVX1 U13612 (.I(N7017), .ZN(n26484));
    INVX1 U13613 (.I(n18951), .ZN(n26485));
    NOR2X1 U13614 (.A1(n24908), .A2(n21673), .ZN(n26486));
    NOR2X1 U13615 (.A1(n15604), .A2(n23150), .ZN(n26487));
    NOR2X1 U13616 (.A1(N5465), .A2(N7332), .ZN(n26488));
    INVX1 U13617 (.I(n13680), .ZN(n26489));
    NANDX1 U13618 (.A1(N710), .A2(N11952), .ZN(N26490));
    INVX1 U13619 (.I(n22899), .ZN(n26491));
    NOR2X1 U13620 (.A1(N11424), .A2(n20398), .ZN(N26492));
    NANDX1 U13621 (.A1(N490), .A2(N2478), .ZN(n26493));
    INVX1 U13622 (.I(n15721), .ZN(N26494));
    INVX1 U13623 (.I(n23974), .ZN(n26495));
    INVX1 U13624 (.I(N3904), .ZN(N26496));
    NANDX1 U13625 (.A1(n17315), .A2(N11623), .ZN(n26497));
    INVX1 U13626 (.I(N5488), .ZN(n26498));
    INVX1 U13627 (.I(n15511), .ZN(N26499));
    NANDX1 U13628 (.A1(N5440), .A2(n23793), .ZN(N26500));
    INVX1 U13629 (.I(N12771), .ZN(n26501));
    NOR2X1 U13630 (.A1(n17771), .A2(N1163), .ZN(n26502));
    NANDX1 U13631 (.A1(n18490), .A2(N8485), .ZN(N26503));
    NANDX1 U13632 (.A1(N4597), .A2(N8676), .ZN(n26504));
    NANDX1 U13633 (.A1(n17553), .A2(n23436), .ZN(N26505));
    NOR2X1 U13634 (.A1(n15663), .A2(n13654), .ZN(n26506));
    NOR2X1 U13635 (.A1(n14134), .A2(N12032), .ZN(n26507));
    NOR2X1 U13636 (.A1(N8390), .A2(n18115), .ZN(n26508));
    INVX1 U13637 (.I(N7050), .ZN(n26509));
    INVX1 U13638 (.I(N1497), .ZN(n26510));
    NOR2X1 U13639 (.A1(N7959), .A2(n21207), .ZN(n26511));
    NOR2X1 U13640 (.A1(n23282), .A2(N8475), .ZN(n26512));
    NOR2X1 U13641 (.A1(N4318), .A2(n23907), .ZN(n26513));
    NANDX1 U13642 (.A1(n22808), .A2(n21160), .ZN(N26514));
    NOR2X1 U13643 (.A1(N1902), .A2(n18603), .ZN(N26515));
    NANDX1 U13644 (.A1(N8222), .A2(n16536), .ZN(n26516));
    NANDX1 U13645 (.A1(N12652), .A2(n18958), .ZN(n26517));
    NANDX1 U13646 (.A1(n15554), .A2(n19757), .ZN(N26518));
    INVX1 U13647 (.I(n23943), .ZN(n26519));
    NOR2X1 U13648 (.A1(N9056), .A2(n19760), .ZN(n26520));
    INVX1 U13649 (.I(N10553), .ZN(N26521));
    INVX1 U13650 (.I(n18427), .ZN(N26522));
    INVX1 U13651 (.I(n18242), .ZN(N26523));
    NANDX1 U13652 (.A1(N3499), .A2(N1547), .ZN(N26524));
    INVX1 U13653 (.I(n16174), .ZN(n26525));
    NOR2X1 U13654 (.A1(n20866), .A2(N599), .ZN(n26526));
    NOR2X1 U13655 (.A1(N11536), .A2(n19201), .ZN(n26527));
    NANDX1 U13656 (.A1(n19757), .A2(n24505), .ZN(N26528));
    INVX1 U13657 (.I(N6907), .ZN(N26529));
    INVX1 U13658 (.I(N6868), .ZN(n26530));
    INVX1 U13659 (.I(N982), .ZN(N26531));
    INVX1 U13660 (.I(N9668), .ZN(n26532));
    NOR2X1 U13661 (.A1(n20043), .A2(N3925), .ZN(n26533));
    INVX1 U13662 (.I(n19363), .ZN(N26534));
    INVX1 U13663 (.I(n19781), .ZN(N26535));
    INVX1 U13664 (.I(N5288), .ZN(n26536));
    INVX1 U13665 (.I(n17886), .ZN(N26537));
    INVX1 U13666 (.I(N11580), .ZN(n26538));
    INVX1 U13667 (.I(N5854), .ZN(n26539));
    NOR2X1 U13668 (.A1(n23425), .A2(N10873), .ZN(N26540));
    NANDX1 U13669 (.A1(n17123), .A2(n14080), .ZN(N26541));
    NANDX1 U13670 (.A1(n16125), .A2(n24412), .ZN(n26542));
    NOR2X1 U13671 (.A1(n22852), .A2(N5777), .ZN(n26543));
    INVX1 U13672 (.I(n23834), .ZN(n26544));
    NANDX1 U13673 (.A1(n21107), .A2(N450), .ZN(n26545));
    INVX1 U13674 (.I(n25032), .ZN(n26546));
    NANDX1 U13675 (.A1(N8203), .A2(N12078), .ZN(n26547));
    INVX1 U13676 (.I(n22590), .ZN(n26548));
    NOR2X1 U13677 (.A1(n23873), .A2(n14973), .ZN(n26549));
    NOR2X1 U13678 (.A1(n24220), .A2(N12297), .ZN(n26550));
    INVX1 U13679 (.I(N8699), .ZN(N26551));
    INVX1 U13680 (.I(N7229), .ZN(n26552));
    INVX1 U13681 (.I(n16109), .ZN(N26553));
    NOR2X1 U13682 (.A1(N9252), .A2(n21002), .ZN(n26554));
    NANDX1 U13683 (.A1(n20696), .A2(N7119), .ZN(n26555));
    NOR2X1 U13684 (.A1(N6634), .A2(N5450), .ZN(n26556));
    NANDX1 U13685 (.A1(N2238), .A2(n20169), .ZN(n26557));
    NOR2X1 U13686 (.A1(n16037), .A2(N10740), .ZN(N26558));
    NOR2X1 U13687 (.A1(n16882), .A2(n21091), .ZN(n26559));
    INVX1 U13688 (.I(n23015), .ZN(n26560));
    INVX1 U13689 (.I(n18162), .ZN(n26561));
    INVX1 U13690 (.I(N6947), .ZN(N26562));
    INVX1 U13691 (.I(n21105), .ZN(N26563));
    NANDX1 U13692 (.A1(n18212), .A2(n17101), .ZN(n26564));
    NOR2X1 U13693 (.A1(n23089), .A2(n12906), .ZN(n26565));
    NOR2X1 U13694 (.A1(n18588), .A2(n21890), .ZN(n26566));
    NOR2X1 U13695 (.A1(n14474), .A2(N11149), .ZN(n26567));
    INVX1 U13696 (.I(N8692), .ZN(n26568));
    NANDX1 U13697 (.A1(N11209), .A2(N3358), .ZN(n26569));
    INVX1 U13698 (.I(N1743), .ZN(N26570));
    NANDX1 U13699 (.A1(n21173), .A2(n18625), .ZN(N26571));
    INVX1 U13700 (.I(n24363), .ZN(n26572));
    NANDX1 U13701 (.A1(N6683), .A2(n17022), .ZN(N26573));
    NOR2X1 U13702 (.A1(N2397), .A2(N10746), .ZN(N26574));
    NANDX1 U13703 (.A1(N6809), .A2(n17725), .ZN(N26575));
    NOR2X1 U13704 (.A1(N4702), .A2(n15311), .ZN(n26576));
    NANDX1 U13705 (.A1(n23078), .A2(n22666), .ZN(N26577));
    INVX1 U13706 (.I(n25416), .ZN(n26578));
    NANDX1 U13707 (.A1(N3599), .A2(n23154), .ZN(n26579));
    NOR2X1 U13708 (.A1(n23807), .A2(N8860), .ZN(n26580));
    NANDX1 U13709 (.A1(N2143), .A2(n24873), .ZN(n26581));
    NOR2X1 U13710 (.A1(N12084), .A2(n17995), .ZN(n26582));
    NANDX1 U13711 (.A1(N10944), .A2(n22899), .ZN(n26583));
    INVX1 U13712 (.I(n16733), .ZN(n26584));
    NANDX1 U13713 (.A1(N8581), .A2(n16246), .ZN(n26585));
    NOR2X1 U13714 (.A1(n15389), .A2(N8469), .ZN(n26586));
    NOR2X1 U13715 (.A1(n20091), .A2(n23779), .ZN(n26587));
    NANDX1 U13716 (.A1(N6434), .A2(N9711), .ZN(n26588));
    NANDX1 U13717 (.A1(n20617), .A2(n21348), .ZN(n26589));
    NOR2X1 U13718 (.A1(n18269), .A2(N4942), .ZN(n26590));
    NANDX1 U13719 (.A1(n15896), .A2(n17395), .ZN(n26591));
    NANDX1 U13720 (.A1(n15266), .A2(n18444), .ZN(N26592));
    INVX1 U13721 (.I(n22028), .ZN(N26593));
    NOR2X1 U13722 (.A1(N3081), .A2(N8192), .ZN(N26594));
    NOR2X1 U13723 (.A1(n19813), .A2(n24009), .ZN(n26595));
    NOR2X1 U13724 (.A1(N10557), .A2(N2844), .ZN(n26596));
    NOR2X1 U13725 (.A1(N7793), .A2(N1571), .ZN(n26597));
    INVX1 U13726 (.I(n20339), .ZN(n26598));
    NANDX1 U13727 (.A1(N4192), .A2(N4547), .ZN(n26599));
    NANDX1 U13728 (.A1(n13576), .A2(N392), .ZN(n26600));
    NANDX1 U13729 (.A1(n20612), .A2(N5333), .ZN(n26601));
    NOR2X1 U13730 (.A1(N11006), .A2(N11496), .ZN(n26602));
    INVX1 U13731 (.I(n15039), .ZN(N26603));
    NOR2X1 U13732 (.A1(n17437), .A2(N11565), .ZN(n26604));
    NANDX1 U13733 (.A1(n20517), .A2(n19756), .ZN(n26605));
    NANDX1 U13734 (.A1(N3596), .A2(N7030), .ZN(n26606));
    INVX1 U13735 (.I(n14152), .ZN(n26607));
    NANDX1 U13736 (.A1(N727), .A2(N10712), .ZN(n26608));
    NOR2X1 U13737 (.A1(n23987), .A2(N5548), .ZN(N26609));
    NOR2X1 U13738 (.A1(n16946), .A2(N10095), .ZN(n26610));
    INVX1 U13739 (.I(N5019), .ZN(N26611));
    INVX1 U13740 (.I(N10774), .ZN(n26612));
    NANDX1 U13741 (.A1(n18857), .A2(N8053), .ZN(n26613));
    NOR2X1 U13742 (.A1(N4850), .A2(N7851), .ZN(n26614));
    INVX1 U13743 (.I(n23556), .ZN(n26615));
    NANDX1 U13744 (.A1(N1002), .A2(n23473), .ZN(n26616));
    NANDX1 U13745 (.A1(N9526), .A2(N10785), .ZN(n26617));
    NOR2X1 U13746 (.A1(n16555), .A2(n22612), .ZN(n26618));
    NANDX1 U13747 (.A1(n15196), .A2(N12106), .ZN(n26619));
    NANDX1 U13748 (.A1(n15408), .A2(N10590), .ZN(N26620));
    NOR2X1 U13749 (.A1(N748), .A2(N2033), .ZN(n26621));
    NANDX1 U13750 (.A1(N3385), .A2(n21322), .ZN(n26622));
    INVX1 U13751 (.I(N2926), .ZN(n26623));
    INVX1 U13752 (.I(N12080), .ZN(n26624));
    NANDX1 U13753 (.A1(N10119), .A2(N5697), .ZN(N26625));
    NANDX1 U13754 (.A1(n25058), .A2(N3750), .ZN(n26626));
    INVX1 U13755 (.I(n14828), .ZN(n26627));
    INVX1 U13756 (.I(n19488), .ZN(n26628));
    INVX1 U13757 (.I(n15542), .ZN(N26629));
    NANDX1 U13758 (.A1(N4173), .A2(N12651), .ZN(N26630));
    INVX1 U13759 (.I(N8137), .ZN(N26631));
    NOR2X1 U13760 (.A1(N11793), .A2(n23544), .ZN(n26632));
    NANDX1 U13761 (.A1(N6900), .A2(n13059), .ZN(n26633));
    INVX1 U13762 (.I(N870), .ZN(n26634));
    NANDX1 U13763 (.A1(N10733), .A2(n19595), .ZN(n26635));
    NOR2X1 U13764 (.A1(n20950), .A2(n20442), .ZN(n26636));
    INVX1 U13765 (.I(n19836), .ZN(N26637));
    NOR2X1 U13766 (.A1(n15477), .A2(n19392), .ZN(n26638));
    NOR2X1 U13767 (.A1(N393), .A2(N8717), .ZN(n26639));
    NOR2X1 U13768 (.A1(n19880), .A2(n21837), .ZN(N26640));
    NANDX1 U13769 (.A1(n15297), .A2(N507), .ZN(n26641));
    INVX1 U13770 (.I(N795), .ZN(n26642));
    NANDX1 U13771 (.A1(n14122), .A2(N1355), .ZN(n26643));
    INVX1 U13772 (.I(N1501), .ZN(N26644));
    NOR2X1 U13773 (.A1(N8510), .A2(n16415), .ZN(n26645));
    NANDX1 U13774 (.A1(n13720), .A2(n15915), .ZN(n26646));
    NOR2X1 U13775 (.A1(n21855), .A2(N131), .ZN(n26647));
    NANDX1 U13776 (.A1(N4234), .A2(n19966), .ZN(n26648));
    INVX1 U13777 (.I(n19710), .ZN(N26649));
    NOR2X1 U13778 (.A1(N9249), .A2(n20102), .ZN(n26650));
    NOR2X1 U13779 (.A1(n18390), .A2(N3247), .ZN(n26651));
    INVX1 U13780 (.I(n17570), .ZN(n26652));
    NANDX1 U13781 (.A1(n22450), .A2(N6936), .ZN(n26653));
    INVX1 U13782 (.I(N5590), .ZN(n26654));
    NANDX1 U13783 (.A1(n20691), .A2(n15312), .ZN(n26655));
    NOR2X1 U13784 (.A1(n17712), .A2(n23821), .ZN(N26656));
    NOR2X1 U13785 (.A1(n15603), .A2(N807), .ZN(n26657));
    INVX1 U13786 (.I(n21855), .ZN(n26658));
    NOR2X1 U13787 (.A1(n21321), .A2(N11815), .ZN(N26659));
    INVX1 U13788 (.I(n15784), .ZN(N26660));
    INVX1 U13789 (.I(N9869), .ZN(n26661));
    NANDX1 U13790 (.A1(N11658), .A2(n18738), .ZN(N26662));
    NANDX1 U13791 (.A1(N4545), .A2(n21984), .ZN(n26663));
    NOR2X1 U13792 (.A1(N10883), .A2(n15024), .ZN(n26664));
    NOR2X1 U13793 (.A1(n17818), .A2(n23128), .ZN(n26665));
    NANDX1 U13794 (.A1(N2141), .A2(n18316), .ZN(n26666));
    NANDX1 U13795 (.A1(n13467), .A2(n24796), .ZN(n26667));
    INVX1 U13796 (.I(N4472), .ZN(N26668));
    NOR2X1 U13797 (.A1(N9462), .A2(N11392), .ZN(n26669));
    INVX1 U13798 (.I(N6620), .ZN(n26670));
    INVX1 U13799 (.I(N598), .ZN(n26671));
    NOR2X1 U13800 (.A1(N11762), .A2(n14239), .ZN(N26672));
    INVX1 U13801 (.I(n18936), .ZN(n26673));
    INVX1 U13802 (.I(N2922), .ZN(n26674));
    NANDX1 U13803 (.A1(n19208), .A2(n24905), .ZN(n26675));
    INVX1 U13804 (.I(N4588), .ZN(n26676));
    INVX1 U13805 (.I(n13297), .ZN(n26677));
    NOR2X1 U13806 (.A1(N820), .A2(n19555), .ZN(n26678));
    INVX1 U13807 (.I(n19136), .ZN(n26679));
    NOR2X1 U13808 (.A1(n15548), .A2(n18429), .ZN(n26680));
    NOR2X1 U13809 (.A1(n20020), .A2(N10860), .ZN(N26681));
    NANDX1 U13810 (.A1(n20179), .A2(n25145), .ZN(n26682));
    NANDX1 U13811 (.A1(n16157), .A2(N241), .ZN(n26683));
    NANDX1 U13812 (.A1(n16686), .A2(N3247), .ZN(n26684));
    NOR2X1 U13813 (.A1(n24389), .A2(n17910), .ZN(n26685));
    INVX1 U13814 (.I(n25102), .ZN(n26686));
    INVX1 U13815 (.I(N12411), .ZN(n26687));
    NOR2X1 U13816 (.A1(N4971), .A2(N4373), .ZN(n26688));
    NOR2X1 U13817 (.A1(N4912), .A2(N5192), .ZN(n26689));
    INVX1 U13818 (.I(N6993), .ZN(n26690));
    INVX1 U13819 (.I(N1502), .ZN(n26691));
    NANDX1 U13820 (.A1(N6021), .A2(N275), .ZN(N26692));
    NOR2X1 U13821 (.A1(n16880), .A2(N8510), .ZN(n26693));
    NANDX1 U13822 (.A1(n16523), .A2(N12132), .ZN(n26694));
    INVX1 U13823 (.I(N5531), .ZN(n26695));
    INVX1 U13824 (.I(N10879), .ZN(n26696));
    NANDX1 U13825 (.A1(N11387), .A2(n24035), .ZN(n26697));
    NOR2X1 U13826 (.A1(n24395), .A2(n23635), .ZN(N26698));
    NOR2X1 U13827 (.A1(N71), .A2(n13399), .ZN(N26699));
    NANDX1 U13828 (.A1(N4443), .A2(N5227), .ZN(n26700));
    NOR2X1 U13829 (.A1(N9634), .A2(n16610), .ZN(N26701));
    NOR2X1 U13830 (.A1(n22729), .A2(n18111), .ZN(N26702));
    INVX1 U13831 (.I(n17517), .ZN(n26703));
    INVX1 U13832 (.I(n13109), .ZN(n26704));
    NOR2X1 U13833 (.A1(n15662), .A2(n16648), .ZN(N26705));
    NANDX1 U13834 (.A1(N2291), .A2(n25112), .ZN(N26706));
    INVX1 U13835 (.I(n14823), .ZN(n26707));
    INVX1 U13836 (.I(n17259), .ZN(n26708));
    NOR2X1 U13837 (.A1(n23291), .A2(n18442), .ZN(n26709));
    INVX1 U13838 (.I(n21423), .ZN(N26710));
    INVX1 U13839 (.I(n13940), .ZN(n26711));
    NOR2X1 U13840 (.A1(n15311), .A2(N7150), .ZN(N26712));
    NANDX1 U13841 (.A1(N1255), .A2(n16783), .ZN(n26713));
    NOR2X1 U13842 (.A1(n22732), .A2(N2777), .ZN(N26714));
    NOR2X1 U13843 (.A1(n15745), .A2(n20294), .ZN(n26715));
    NANDX1 U13844 (.A1(n17621), .A2(n17956), .ZN(n26716));
    NOR2X1 U13845 (.A1(n23037), .A2(n20908), .ZN(N26717));
    INVX1 U13846 (.I(n22646), .ZN(N26718));
    INVX1 U13847 (.I(n15723), .ZN(n26719));
    NOR2X1 U13848 (.A1(N9914), .A2(N5198), .ZN(n26720));
    INVX1 U13849 (.I(N2853), .ZN(N26721));
    NANDX1 U13850 (.A1(N4377), .A2(N11627), .ZN(n26722));
    NANDX1 U13851 (.A1(N2463), .A2(N1435), .ZN(n26723));
    NANDX1 U13852 (.A1(N5776), .A2(n16960), .ZN(n26724));
    NANDX1 U13853 (.A1(N195), .A2(n14189), .ZN(n26725));
    NANDX1 U13854 (.A1(N1493), .A2(N4432), .ZN(N26726));
    INVX1 U13855 (.I(n21175), .ZN(n26727));
    INVX1 U13856 (.I(n16300), .ZN(N26728));
    NANDX1 U13857 (.A1(N8354), .A2(N11705), .ZN(n26729));
    NOR2X1 U13858 (.A1(n19767), .A2(N4360), .ZN(n26730));
    NANDX1 U13859 (.A1(n16166), .A2(n14273), .ZN(n26731));
    NOR2X1 U13860 (.A1(n13390), .A2(N5893), .ZN(n26732));
    NOR2X1 U13861 (.A1(n17767), .A2(n17520), .ZN(n26733));
    INVX1 U13862 (.I(N8997), .ZN(n26734));
    INVX1 U13863 (.I(n18473), .ZN(n26735));
    NOR2X1 U13864 (.A1(N10411), .A2(n16212), .ZN(N26736));
    NOR2X1 U13865 (.A1(n24600), .A2(N5495), .ZN(n26737));
    INVX1 U13866 (.I(n17799), .ZN(n26738));
    NANDX1 U13867 (.A1(N899), .A2(N3116), .ZN(N26739));
    INVX1 U13868 (.I(N9450), .ZN(n26740));
    INVX1 U13869 (.I(n20612), .ZN(N26741));
    INVX1 U13870 (.I(n20004), .ZN(n26742));
    NANDX1 U13871 (.A1(N4304), .A2(N10667), .ZN(N26743));
    NOR2X1 U13872 (.A1(n23443), .A2(n24057), .ZN(n26744));
    NANDX1 U13873 (.A1(n24915), .A2(N5089), .ZN(N26745));
    NANDX1 U13874 (.A1(N11427), .A2(n14085), .ZN(n26746));
    INVX1 U13875 (.I(N4397), .ZN(N26747));
    NOR2X1 U13876 (.A1(N7319), .A2(N9376), .ZN(n26748));
    NOR2X1 U13877 (.A1(N6416), .A2(N3638), .ZN(n26749));
    NOR2X1 U13878 (.A1(n12982), .A2(n21747), .ZN(n26750));
    NANDX1 U13879 (.A1(n16098), .A2(n16384), .ZN(n26751));
    NANDX1 U13880 (.A1(n16335), .A2(N261), .ZN(n26752));
    NANDX1 U13881 (.A1(N10836), .A2(n13999), .ZN(n26753));
    NANDX1 U13882 (.A1(N10271), .A2(n16508), .ZN(n26754));
    NANDX1 U13883 (.A1(n23095), .A2(n24910), .ZN(n26755));
    NOR2X1 U13884 (.A1(n16951), .A2(n14096), .ZN(n26756));
    NOR2X1 U13885 (.A1(n19803), .A2(n22236), .ZN(N26757));
    NANDX1 U13886 (.A1(N11925), .A2(n18323), .ZN(n26758));
    INVX1 U13887 (.I(N7781), .ZN(n26759));
    NANDX1 U13888 (.A1(n15894), .A2(N8863), .ZN(N26760));
    NOR2X1 U13889 (.A1(N12138), .A2(n13881), .ZN(n26761));
    INVX1 U13890 (.I(n17289), .ZN(n26762));
    INVX1 U13891 (.I(N10953), .ZN(n26763));
    NOR2X1 U13892 (.A1(N7675), .A2(N10556), .ZN(n26764));
    NOR2X1 U13893 (.A1(N5575), .A2(n20826), .ZN(N26765));
    INVX1 U13894 (.I(n15685), .ZN(N26766));
    NANDX1 U13895 (.A1(N10728), .A2(N10937), .ZN(n26767));
    NANDX1 U13896 (.A1(n13592), .A2(n20654), .ZN(n26768));
    NANDX1 U13897 (.A1(n24595), .A2(n20496), .ZN(n26769));
    INVX1 U13898 (.I(n17415), .ZN(n26770));
    INVX1 U13899 (.I(N1408), .ZN(N26771));
    NOR2X1 U13900 (.A1(n23143), .A2(n24540), .ZN(n26772));
    NANDX1 U13901 (.A1(N9778), .A2(n12919), .ZN(n26773));
    NANDX1 U13902 (.A1(N1565), .A2(n15765), .ZN(n26774));
    INVX1 U13903 (.I(N7881), .ZN(n26775));
    INVX1 U13904 (.I(N8259), .ZN(N26776));
    NOR2X1 U13905 (.A1(n17781), .A2(n17853), .ZN(N26777));
    NANDX1 U13906 (.A1(N7963), .A2(n25038), .ZN(n26778));
    INVX1 U13907 (.I(N7668), .ZN(n26779));
    NANDX1 U13908 (.A1(N12831), .A2(N2819), .ZN(n26780));
    INVX1 U13909 (.I(N11924), .ZN(N26781));
    NOR2X1 U13910 (.A1(n13270), .A2(n18106), .ZN(n26782));
    INVX1 U13911 (.I(N3445), .ZN(n26783));
    NANDX1 U13912 (.A1(N5739), .A2(N2483), .ZN(N26784));
    NOR2X1 U13913 (.A1(N4285), .A2(N4169), .ZN(N26785));
    NANDX1 U13914 (.A1(N5849), .A2(n19933), .ZN(n26786));
    NANDX1 U13915 (.A1(n13729), .A2(n17869), .ZN(N26787));
    NANDX1 U13916 (.A1(n16423), .A2(n24418), .ZN(n26788));
    NOR2X1 U13917 (.A1(N4935), .A2(n21148), .ZN(N26789));
    NANDX1 U13918 (.A1(N4174), .A2(N3313), .ZN(N26790));
    NOR2X1 U13919 (.A1(n17005), .A2(n20401), .ZN(n26791));
    INVX1 U13920 (.I(n17696), .ZN(n26792));
    INVX1 U13921 (.I(n17987), .ZN(n26793));
    NANDX1 U13922 (.A1(N3847), .A2(n21431), .ZN(N26794));
    NANDX1 U13923 (.A1(n23856), .A2(N12681), .ZN(n26795));
    INVX1 U13924 (.I(N2638), .ZN(n26796));
    NOR2X1 U13925 (.A1(N6959), .A2(n22756), .ZN(n26797));
    NOR2X1 U13926 (.A1(n24377), .A2(n25252), .ZN(N26798));
    NANDX1 U13927 (.A1(n13320), .A2(n16172), .ZN(N26799));
    INVX1 U13928 (.I(n20115), .ZN(N26800));
    INVX1 U13929 (.I(N1244), .ZN(n26801));
    NANDX1 U13930 (.A1(n14048), .A2(n18827), .ZN(n26802));
    NANDX1 U13931 (.A1(n19820), .A2(n13725), .ZN(N26803));
    NOR2X1 U13932 (.A1(N781), .A2(n23743), .ZN(n26804));
    NANDX1 U13933 (.A1(N11079), .A2(N2088), .ZN(n26805));
    INVX1 U13934 (.I(N8167), .ZN(n26806));
    NANDX1 U13935 (.A1(n17329), .A2(n23950), .ZN(n26807));
    INVX1 U13936 (.I(N8675), .ZN(n26808));
    NOR2X1 U13937 (.A1(n14601), .A2(N8722), .ZN(N26809));
    NANDX1 U13938 (.A1(n14350), .A2(N1135), .ZN(n26810));
    NOR2X1 U13939 (.A1(n19290), .A2(N6733), .ZN(n26811));
    NOR2X1 U13940 (.A1(N3661), .A2(n22246), .ZN(n26812));
    NANDX1 U13941 (.A1(N6476), .A2(n15570), .ZN(n26813));
    INVX1 U13942 (.I(N793), .ZN(n26814));
    NANDX1 U13943 (.A1(N10251), .A2(N1573), .ZN(n26815));
    NOR2X1 U13944 (.A1(n18970), .A2(N1420), .ZN(N26816));
    NOR2X1 U13945 (.A1(n23617), .A2(n23856), .ZN(n26817));
    INVX1 U13946 (.I(n15443), .ZN(n26818));
    NOR2X1 U13947 (.A1(n13713), .A2(n24118), .ZN(n26819));
    NOR2X1 U13948 (.A1(N2811), .A2(N7337), .ZN(N26820));
    NANDX1 U13949 (.A1(N5929), .A2(n22741), .ZN(N26821));
    NANDX1 U13950 (.A1(n13986), .A2(n18241), .ZN(N26822));
    NANDX1 U13951 (.A1(N6414), .A2(N3752), .ZN(N26823));
    INVX1 U13952 (.I(n12890), .ZN(n26824));
    NANDX1 U13953 (.A1(n16766), .A2(n13682), .ZN(N26825));
    NOR2X1 U13954 (.A1(N1514), .A2(N4023), .ZN(n26826));
    NOR2X1 U13955 (.A1(n20483), .A2(N5442), .ZN(n26827));
    NOR2X1 U13956 (.A1(N7365), .A2(N3795), .ZN(N26828));
    INVX1 U13957 (.I(n22808), .ZN(n26829));
    INVX1 U13958 (.I(N8686), .ZN(N26830));
    NOR2X1 U13959 (.A1(n20109), .A2(N11496), .ZN(n26831));
    NANDX1 U13960 (.A1(N7168), .A2(N6192), .ZN(N26832));
    NANDX1 U13961 (.A1(n17902), .A2(N8945), .ZN(n26833));
    NANDX1 U13962 (.A1(N7152), .A2(n15359), .ZN(n26834));
    NOR2X1 U13963 (.A1(N4400), .A2(N2746), .ZN(n26835));
    NANDX1 U13964 (.A1(N9933), .A2(N5195), .ZN(n26836));
    INVX1 U13965 (.I(N214), .ZN(N26837));
    INVX1 U13966 (.I(N210), .ZN(n26838));
    NANDX1 U13967 (.A1(n14658), .A2(n24319), .ZN(n26839));
    INVX1 U13968 (.I(N7221), .ZN(n26840));
    NOR2X1 U13969 (.A1(n14133), .A2(n22086), .ZN(n26841));
    NOR2X1 U13970 (.A1(n24323), .A2(n16692), .ZN(n26842));
    NANDX1 U13971 (.A1(N5115), .A2(N12628), .ZN(n26843));
    NANDX1 U13972 (.A1(n22917), .A2(N5027), .ZN(N26844));
    NOR2X1 U13973 (.A1(N7955), .A2(N946), .ZN(N26845));
    NOR2X1 U13974 (.A1(N11015), .A2(N5345), .ZN(n26846));
    NOR2X1 U13975 (.A1(N7893), .A2(n15277), .ZN(n26847));
    NOR2X1 U13976 (.A1(N5421), .A2(n15490), .ZN(n26848));
    NANDX1 U13977 (.A1(n19900), .A2(n24953), .ZN(n26849));
    NANDX1 U13978 (.A1(N7484), .A2(n16279), .ZN(n26850));
    INVX1 U13979 (.I(N1272), .ZN(N26851));
    INVX1 U13980 (.I(N12688), .ZN(n26852));
    INVX1 U13981 (.I(n18000), .ZN(n26853));
    NOR2X1 U13982 (.A1(N9521), .A2(N11882), .ZN(N26854));
    NOR2X1 U13983 (.A1(n21487), .A2(N9297), .ZN(N26855));
    INVX1 U13984 (.I(n16896), .ZN(n26856));
    NOR2X1 U13985 (.A1(N11245), .A2(N2161), .ZN(N26857));
    NANDX1 U13986 (.A1(N5357), .A2(N4441), .ZN(n26858));
    INVX1 U13987 (.I(n20634), .ZN(n26859));
    NOR2X1 U13988 (.A1(n19114), .A2(n24891), .ZN(n26860));
    INVX1 U13989 (.I(n13511), .ZN(n26861));
    NOR2X1 U13990 (.A1(N757), .A2(n20994), .ZN(n26862));
    NOR2X1 U13991 (.A1(n16862), .A2(N11033), .ZN(n26863));
    INVX1 U13992 (.I(N4047), .ZN(N26864));
    NOR2X1 U13993 (.A1(n18599), .A2(n22194), .ZN(N26865));
    NANDX1 U13994 (.A1(n19249), .A2(n13196), .ZN(n26866));
    INVX1 U13995 (.I(N3043), .ZN(n26867));
    NOR2X1 U13996 (.A1(n17752), .A2(N9061), .ZN(n26868));
    NANDX1 U13997 (.A1(n19913), .A2(n14862), .ZN(n26869));
    NOR2X1 U13998 (.A1(n24353), .A2(N3053), .ZN(n26870));
    NANDX1 U13999 (.A1(n25036), .A2(N10934), .ZN(n26871));
    NANDX1 U14000 (.A1(n16908), .A2(n24444), .ZN(n26872));
    NANDX1 U14001 (.A1(N6433), .A2(N8703), .ZN(n26873));
    NANDX1 U14002 (.A1(N12062), .A2(n19735), .ZN(n26874));
    NANDX1 U14003 (.A1(n16108), .A2(N817), .ZN(n26875));
    INVX1 U14004 (.I(N12800), .ZN(n26876));
    NANDX1 U14005 (.A1(n22663), .A2(n14763), .ZN(n26877));
    NANDX1 U14006 (.A1(N203), .A2(N1523), .ZN(n26878));
    NOR2X1 U14007 (.A1(n23533), .A2(n25029), .ZN(n26879));
    NOR2X1 U14008 (.A1(N1660), .A2(N2888), .ZN(N26880));
    NOR2X1 U14009 (.A1(N4712), .A2(n15649), .ZN(n26881));
    NOR2X1 U14010 (.A1(n15645), .A2(n16567), .ZN(n26882));
    NOR2X1 U14011 (.A1(N3354), .A2(n19362), .ZN(n26883));
    NOR2X1 U14012 (.A1(N12056), .A2(n14810), .ZN(n26884));
    NANDX1 U14013 (.A1(n20559), .A2(n25128), .ZN(N26885));
    NANDX1 U14014 (.A1(n21375), .A2(N3040), .ZN(N26886));
    INVX1 U14015 (.I(N1560), .ZN(n26887));
    INVX1 U14016 (.I(N227), .ZN(n26888));
    INVX1 U14017 (.I(n14672), .ZN(n26889));
    NANDX1 U14018 (.A1(n21167), .A2(N1470), .ZN(n26890));
    INVX1 U14019 (.I(N3138), .ZN(n26891));
    NOR2X1 U14020 (.A1(N7201), .A2(N9461), .ZN(n26892));
    NANDX1 U14021 (.A1(N11618), .A2(n15318), .ZN(n26893));
    NANDX1 U14022 (.A1(n16952), .A2(N1349), .ZN(n26894));
    NOR2X1 U14023 (.A1(N10812), .A2(N8081), .ZN(N26895));
    NANDX1 U14024 (.A1(n14389), .A2(N1373), .ZN(N26896));
    NOR2X1 U14025 (.A1(n14014), .A2(N10772), .ZN(n26897));
    NOR2X1 U14026 (.A1(N5821), .A2(n21738), .ZN(n26898));
    INVX1 U14027 (.I(n20290), .ZN(N26899));
    NOR2X1 U14028 (.A1(N11865), .A2(n23729), .ZN(n26900));
    NANDX1 U14029 (.A1(N7529), .A2(n13967), .ZN(n26901));
    NOR2X1 U14030 (.A1(N10666), .A2(N5864), .ZN(n26902));
    NANDX1 U14031 (.A1(n20127), .A2(N2472), .ZN(N26903));
    NANDX1 U14032 (.A1(n24212), .A2(n17763), .ZN(N26904));
    NANDX1 U14033 (.A1(N58), .A2(N10906), .ZN(N26905));
    NOR2X1 U14034 (.A1(n22409), .A2(n16104), .ZN(n26906));
    NOR2X1 U14035 (.A1(n23781), .A2(n19396), .ZN(N26907));
    NANDX1 U14036 (.A1(N9050), .A2(n18560), .ZN(n26908));
    INVX1 U14037 (.I(n19555), .ZN(N26909));
    NOR2X1 U14038 (.A1(n21955), .A2(N4784), .ZN(n26910));
    INVX1 U14039 (.I(N8949), .ZN(n26911));
    NANDX1 U14040 (.A1(n16212), .A2(n22915), .ZN(N26912));
    NANDX1 U14041 (.A1(N1376), .A2(N3276), .ZN(N26913));
    INVX1 U14042 (.I(N10270), .ZN(n26914));
    INVX1 U14043 (.I(N8965), .ZN(n26915));
    NANDX1 U14044 (.A1(N12278), .A2(n24794), .ZN(n26916));
    NANDX1 U14045 (.A1(n23183), .A2(n14700), .ZN(n26917));
    NANDX1 U14046 (.A1(N2552), .A2(n18994), .ZN(n26918));
    NANDX1 U14047 (.A1(n21947), .A2(N568), .ZN(n26919));
    INVX1 U14048 (.I(n15004), .ZN(n26920));
    NOR2X1 U14049 (.A1(n24630), .A2(n23055), .ZN(N26921));
    NANDX1 U14050 (.A1(N3911), .A2(N6236), .ZN(n26922));
    NOR2X1 U14051 (.A1(n24213), .A2(n22447), .ZN(N26923));
    NOR2X1 U14052 (.A1(n24575), .A2(N12590), .ZN(N26924));
    NOR2X1 U14053 (.A1(n23430), .A2(n22859), .ZN(n26925));
    INVX1 U14054 (.I(n21162), .ZN(n26926));
    NOR2X1 U14055 (.A1(N3882), .A2(n20453), .ZN(n26927));
    INVX1 U14056 (.I(N1562), .ZN(n26928));
    NANDX1 U14057 (.A1(N1888), .A2(N4114), .ZN(n26929));
    NANDX1 U14058 (.A1(n20378), .A2(N558), .ZN(N26930));
    NANDX1 U14059 (.A1(n25453), .A2(n15562), .ZN(N26931));
    INVX1 U14060 (.I(n24580), .ZN(n26932));
    NOR2X1 U14061 (.A1(n18895), .A2(n17258), .ZN(n26933));
    NOR2X1 U14062 (.A1(N1025), .A2(N4737), .ZN(n26934));
    NANDX1 U14063 (.A1(n20340), .A2(n18079), .ZN(n26935));
    NOR2X1 U14064 (.A1(N3159), .A2(n16006), .ZN(n26936));
    NANDX1 U14065 (.A1(n20264), .A2(N11665), .ZN(n26937));
    INVX1 U14066 (.I(n24145), .ZN(n26938));
    NOR2X1 U14067 (.A1(n20325), .A2(n14475), .ZN(N26939));
    INVX1 U14068 (.I(n22212), .ZN(N26940));
    INVX1 U14069 (.I(n22443), .ZN(n26941));
    NANDX1 U14070 (.A1(N7913), .A2(n14919), .ZN(N26942));
    NOR2X1 U14071 (.A1(n23474), .A2(N9627), .ZN(n26943));
    NOR2X1 U14072 (.A1(n14123), .A2(N3019), .ZN(n26944));
    NANDX1 U14073 (.A1(n25277), .A2(n18313), .ZN(N26945));
    INVX1 U14074 (.I(N7874), .ZN(n26946));
    NOR2X1 U14075 (.A1(N11258), .A2(N3060), .ZN(n26947));
    NANDX1 U14076 (.A1(N1762), .A2(n21104), .ZN(n26948));
    NANDX1 U14077 (.A1(N2194), .A2(n23020), .ZN(n26949));
    INVX1 U14078 (.I(n23079), .ZN(N26950));
    NOR2X1 U14079 (.A1(n15993), .A2(N2608), .ZN(n26951));
    INVX1 U14080 (.I(N9078), .ZN(n26952));
    INVX1 U14081 (.I(n20406), .ZN(n26953));
    INVX1 U14082 (.I(n17504), .ZN(N26954));
    NOR2X1 U14083 (.A1(N3730), .A2(N1628), .ZN(N26955));
    NOR2X1 U14084 (.A1(N6620), .A2(n18916), .ZN(n26956));
    INVX1 U14085 (.I(N6395), .ZN(N26957));
    NANDX1 U14086 (.A1(n15752), .A2(n14268), .ZN(n26958));
    INVX1 U14087 (.I(N1508), .ZN(n26959));
    NANDX1 U14088 (.A1(N4451), .A2(n17539), .ZN(n26960));
    NANDX1 U14089 (.A1(n18558), .A2(n19732), .ZN(N26961));
    NOR2X1 U14090 (.A1(n20076), .A2(n17308), .ZN(n26962));
    NOR2X1 U14091 (.A1(n24836), .A2(N8684), .ZN(n26963));
    INVX1 U14092 (.I(N8411), .ZN(N26964));
    NOR2X1 U14093 (.A1(n15277), .A2(n14169), .ZN(n26965));
    NOR2X1 U14094 (.A1(n19023), .A2(N6666), .ZN(n26966));
    INVX1 U14095 (.I(n16419), .ZN(n26967));
    NOR2X1 U14096 (.A1(n23814), .A2(n13489), .ZN(n26968));
    NANDX1 U14097 (.A1(n24308), .A2(n18009), .ZN(n26969));
    NANDX1 U14098 (.A1(n23682), .A2(N8284), .ZN(n26970));
    INVX1 U14099 (.I(n16900), .ZN(N26971));
    NANDX1 U14100 (.A1(N8040), .A2(n24225), .ZN(n26972));
    INVX1 U14101 (.I(N7252), .ZN(N26973));
    INVX1 U14102 (.I(n14895), .ZN(n26974));
    NOR2X1 U14103 (.A1(N6900), .A2(n23578), .ZN(n26975));
    INVX1 U14104 (.I(N4079), .ZN(n26976));
    INVX1 U14105 (.I(N758), .ZN(n26977));
    INVX1 U14106 (.I(N1382), .ZN(n26978));
    NANDX1 U14107 (.A1(n13680), .A2(n20550), .ZN(n26979));
    NOR2X1 U14108 (.A1(n15732), .A2(n18861), .ZN(n26980));
    NOR2X1 U14109 (.A1(N1715), .A2(N6434), .ZN(n26981));
    INVX1 U14110 (.I(N1964), .ZN(n26982));
    NANDX1 U14111 (.A1(N2510), .A2(n19540), .ZN(n26983));
    INVX1 U14112 (.I(n17099), .ZN(N26984));
    NANDX1 U14113 (.A1(N9002), .A2(N415), .ZN(n26985));
    NANDX1 U14114 (.A1(n16568), .A2(N4077), .ZN(N26986));
    NANDX1 U14115 (.A1(N12236), .A2(N2152), .ZN(N26987));
    NOR2X1 U14116 (.A1(n16314), .A2(N264), .ZN(N26988));
    NOR2X1 U14117 (.A1(n23328), .A2(n15915), .ZN(N26989));
    NANDX1 U14118 (.A1(N11505), .A2(N10962), .ZN(n26990));
    NANDX1 U14119 (.A1(n16004), .A2(n18590), .ZN(N26991));
    NANDX1 U14120 (.A1(n17718), .A2(n25023), .ZN(N26992));
    NANDX1 U14121 (.A1(N8450), .A2(n18403), .ZN(N26993));
    INVX1 U14122 (.I(n16757), .ZN(n26994));
    NOR2X1 U14123 (.A1(N9739), .A2(N7601), .ZN(n26995));
    NOR2X1 U14124 (.A1(N10154), .A2(n19966), .ZN(n26996));
    NOR2X1 U14125 (.A1(n14230), .A2(N8671), .ZN(N26997));
    NANDX1 U14126 (.A1(N5150), .A2(n19591), .ZN(n26998));
    NOR2X1 U14127 (.A1(n19683), .A2(N5765), .ZN(N26999));
    NANDX1 U14128 (.A1(n24365), .A2(N11719), .ZN(n27000));
    NOR2X1 U14129 (.A1(N9825), .A2(N5905), .ZN(N27001));
    NOR2X1 U14130 (.A1(N2912), .A2(n13042), .ZN(N27002));
    NANDX1 U14131 (.A1(n16703), .A2(n14406), .ZN(n27003));
    INVX1 U14132 (.I(N9603), .ZN(N27004));
    NOR2X1 U14133 (.A1(n18388), .A2(N1551), .ZN(n27005));
    NOR2X1 U14134 (.A1(N486), .A2(n16770), .ZN(n27006));
    NANDX1 U14135 (.A1(N9220), .A2(N11822), .ZN(n27007));
    NANDX1 U14136 (.A1(n17890), .A2(N4840), .ZN(n27008));
    NANDX1 U14137 (.A1(N11978), .A2(N2938), .ZN(n27009));
    INVX1 U14138 (.I(N6511), .ZN(N27010));
    NOR2X1 U14139 (.A1(n19933), .A2(N6997), .ZN(n27011));
    NOR2X1 U14140 (.A1(N4255), .A2(n12901), .ZN(n27012));
    NANDX1 U14141 (.A1(n21436), .A2(N441), .ZN(N27013));
    NANDX1 U14142 (.A1(N12636), .A2(N3614), .ZN(N27014));
    NOR2X1 U14143 (.A1(N11007), .A2(N10659), .ZN(n27015));
    INVX1 U14144 (.I(N1325), .ZN(N27016));
    INVX1 U14145 (.I(N12749), .ZN(n27017));
    NOR2X1 U14146 (.A1(n17646), .A2(N10736), .ZN(n27018));
    NOR2X1 U14147 (.A1(N10847), .A2(N3124), .ZN(n27019));
    NANDX1 U14148 (.A1(n23466), .A2(N3869), .ZN(n27020));
    NOR2X1 U14149 (.A1(n19034), .A2(N10379), .ZN(N27021));
    NANDX1 U14150 (.A1(N2232), .A2(N6144), .ZN(n27022));
    NANDX1 U14151 (.A1(N6486), .A2(n19044), .ZN(N27023));
    INVX1 U14152 (.I(n16689), .ZN(N27024));
    NANDX1 U14153 (.A1(N8645), .A2(n18093), .ZN(N27025));
    INVX1 U14154 (.I(n13752), .ZN(n27026));
    INVX1 U14155 (.I(N11292), .ZN(N27027));
    NOR2X1 U14156 (.A1(n19191), .A2(n13232), .ZN(n27028));
    NOR2X1 U14157 (.A1(N550), .A2(n19646), .ZN(n27029));
    NOR2X1 U14158 (.A1(n19232), .A2(n19260), .ZN(n27030));
    NOR2X1 U14159 (.A1(N6020), .A2(N5991), .ZN(n27031));
    INVX1 U14160 (.I(N10015), .ZN(n27032));
    NANDX1 U14161 (.A1(N7671), .A2(n24103), .ZN(n27033));
    INVX1 U14162 (.I(n13814), .ZN(N27034));
    NOR2X1 U14163 (.A1(N11276), .A2(N7356), .ZN(N27035));
    INVX1 U14164 (.I(N2463), .ZN(N27036));
    INVX1 U14165 (.I(n13363), .ZN(n27037));
    NOR2X1 U14166 (.A1(n16240), .A2(N1613), .ZN(N27038));
    INVX1 U14167 (.I(n16299), .ZN(n27039));
    NANDX1 U14168 (.A1(N6607), .A2(N4028), .ZN(N27040));
    NANDX1 U14169 (.A1(N7156), .A2(N12441), .ZN(N27041));
    NANDX1 U14170 (.A1(n15155), .A2(N6198), .ZN(N27042));
    NANDX1 U14171 (.A1(N9942), .A2(N957), .ZN(n27043));
    NANDX1 U14172 (.A1(n19956), .A2(n14748), .ZN(n27044));
    NOR2X1 U14173 (.A1(N7324), .A2(N5269), .ZN(N27045));
    INVX1 U14174 (.I(n18107), .ZN(N27046));
    NANDX1 U14175 (.A1(n22203), .A2(n22825), .ZN(N27047));
    INVX1 U14176 (.I(N1076), .ZN(N27048));
    NANDX1 U14177 (.A1(n17096), .A2(N6083), .ZN(n27049));
    INVX1 U14178 (.I(N4512), .ZN(n27050));
    INVX1 U14179 (.I(N3190), .ZN(n27051));
    INVX1 U14180 (.I(n15176), .ZN(n27052));
    NOR2X1 U14181 (.A1(n21311), .A2(N2115), .ZN(n27053));
    NANDX1 U14182 (.A1(n25234), .A2(n22582), .ZN(n27054));
    INVX1 U14183 (.I(N9673), .ZN(n27055));
    INVX1 U14184 (.I(N5503), .ZN(n27056));
    INVX1 U14185 (.I(N1552), .ZN(n27057));
    INVX1 U14186 (.I(N11450), .ZN(N27058));
    INVX1 U14187 (.I(n21384), .ZN(n27059));
    INVX1 U14188 (.I(N899), .ZN(n27060));
    INVX1 U14189 (.I(N1377), .ZN(N27061));
    NOR2X1 U14190 (.A1(n22198), .A2(N830), .ZN(n27062));
    INVX1 U14191 (.I(n17048), .ZN(N27063));
    NANDX1 U14192 (.A1(N7816), .A2(n13926), .ZN(n27064));
    INVX1 U14193 (.I(N7701), .ZN(N27065));
    INVX1 U14194 (.I(n15465), .ZN(n27066));
    NANDX1 U14195 (.A1(N8751), .A2(N6030), .ZN(n27067));
    NOR2X1 U14196 (.A1(n20101), .A2(N6937), .ZN(n27068));
    INVX1 U14197 (.I(n18136), .ZN(n27069));
    NANDX1 U14198 (.A1(N5807), .A2(n19687), .ZN(n27070));
    NANDX1 U14199 (.A1(N6025), .A2(N4042), .ZN(N27071));
    NOR2X1 U14200 (.A1(N10078), .A2(N4941), .ZN(n27072));
    NOR2X1 U14201 (.A1(N222), .A2(N2381), .ZN(N27073));
    INVX1 U14202 (.I(N1051), .ZN(N27074));
    NANDX1 U14203 (.A1(n12986), .A2(N2945), .ZN(N27075));
    INVX1 U14204 (.I(n15679), .ZN(n27076));
    NOR2X1 U14205 (.A1(n21200), .A2(N8046), .ZN(n27077));
    INVX1 U14206 (.I(n13477), .ZN(N27078));
    INVX1 U14207 (.I(n21329), .ZN(N27079));
    INVX1 U14208 (.I(N162), .ZN(n27080));
    NOR2X1 U14209 (.A1(N7165), .A2(n18298), .ZN(n27081));
    INVX1 U14210 (.I(n12972), .ZN(n27082));
    NOR2X1 U14211 (.A1(n22943), .A2(n18996), .ZN(n27083));
    NOR2X1 U14212 (.A1(n15334), .A2(n17841), .ZN(n27084));
    NANDX1 U14213 (.A1(N308), .A2(N6831), .ZN(n27085));
    NOR2X1 U14214 (.A1(n21748), .A2(n22151), .ZN(n27086));
    INVX1 U14215 (.I(n23502), .ZN(n27087));
    NOR2X1 U14216 (.A1(N6292), .A2(n13678), .ZN(N27088));
    NOR2X1 U14217 (.A1(N1989), .A2(n21723), .ZN(n27089));
    INVX1 U14218 (.I(n15465), .ZN(N27090));
    NANDX1 U14219 (.A1(N10552), .A2(n20949), .ZN(N27091));
    NOR2X1 U14220 (.A1(n13314), .A2(n16881), .ZN(n27092));
    INVX1 U14221 (.I(n17282), .ZN(n27093));
    NOR2X1 U14222 (.A1(n13299), .A2(N3490), .ZN(N27094));
    NANDX1 U14223 (.A1(N7358), .A2(n18824), .ZN(n27095));
    NOR2X1 U14224 (.A1(N6357), .A2(N7899), .ZN(n27096));
    INVX1 U14225 (.I(N7736), .ZN(n27097));
    INVX1 U14226 (.I(N10968), .ZN(n27098));
    NOR2X1 U14227 (.A1(n16413), .A2(n13599), .ZN(n27099));
    NOR2X1 U14228 (.A1(N4589), .A2(n13026), .ZN(n27100));
    INVX1 U14229 (.I(n15079), .ZN(n27101));
    NANDX1 U14230 (.A1(N4845), .A2(N5631), .ZN(n27102));
    NOR2X1 U14231 (.A1(N291), .A2(n21847), .ZN(n27103));
    NANDX1 U14232 (.A1(n17172), .A2(n19625), .ZN(n27104));
    NOR2X1 U14233 (.A1(N10289), .A2(n21691), .ZN(n27105));
    NOR2X1 U14234 (.A1(N11170), .A2(N3546), .ZN(N27106));
    INVX1 U14235 (.I(N4389), .ZN(n27107));
    NANDX1 U14236 (.A1(n14409), .A2(N7476), .ZN(n27108));
    INVX1 U14237 (.I(N7320), .ZN(n27109));
    INVX1 U14238 (.I(N9971), .ZN(n27110));
    NANDX1 U14239 (.A1(n20810), .A2(n19827), .ZN(n27111));
    NOR2X1 U14240 (.A1(n22603), .A2(n20440), .ZN(n27112));
    INVX1 U14241 (.I(n13620), .ZN(n27113));
    NOR2X1 U14242 (.A1(N12296), .A2(n15189), .ZN(N27114));
    NOR2X1 U14243 (.A1(N8640), .A2(N7607), .ZN(n27115));
    INVX1 U14244 (.I(n17032), .ZN(n27116));
    NANDX1 U14245 (.A1(n19338), .A2(n13221), .ZN(n27117));
    NANDX1 U14246 (.A1(N5005), .A2(N5534), .ZN(N27118));
    NANDX1 U14247 (.A1(n23663), .A2(n15436), .ZN(n27119));
    NOR2X1 U14248 (.A1(N5636), .A2(N10608), .ZN(N27120));
    INVX1 U14249 (.I(N12847), .ZN(n27121));
    INVX1 U14250 (.I(n20229), .ZN(n27122));
    NOR2X1 U14251 (.A1(N3671), .A2(N11815), .ZN(n27123));
    NANDX1 U14252 (.A1(n12878), .A2(n18479), .ZN(n27124));
    INVX1 U14253 (.I(N12659), .ZN(n27125));
    INVX1 U14254 (.I(n22830), .ZN(n27126));
    INVX1 U14255 (.I(N2679), .ZN(n27127));
    NOR2X1 U14256 (.A1(n24818), .A2(n19711), .ZN(N27128));
    NANDX1 U14257 (.A1(n18654), .A2(n21699), .ZN(N27129));
    INVX1 U14258 (.I(n23658), .ZN(N27130));
    NANDX1 U14259 (.A1(N2000), .A2(N10587), .ZN(n27131));
    INVX1 U14260 (.I(n16679), .ZN(n27132));
    NOR2X1 U14261 (.A1(n16541), .A2(n13175), .ZN(N27133));
    INVX1 U14262 (.I(N384), .ZN(N27134));
    NOR2X1 U14263 (.A1(N487), .A2(N4054), .ZN(N27135));
    INVX1 U14264 (.I(n20011), .ZN(N27136));
    NANDX1 U14265 (.A1(N1459), .A2(N2150), .ZN(n27137));
    INVX1 U14266 (.I(N6731), .ZN(n27138));
    INVX1 U14267 (.I(n22894), .ZN(n27139));
    NANDX1 U14268 (.A1(N7448), .A2(n22210), .ZN(n27140));
    NANDX1 U14269 (.A1(n18454), .A2(N4129), .ZN(n27141));
    INVX1 U14270 (.I(n20183), .ZN(N27142));
    NOR2X1 U14271 (.A1(N4581), .A2(N10951), .ZN(n27143));
    NANDX1 U14272 (.A1(N10513), .A2(N2127), .ZN(n27144));
    NANDX1 U14273 (.A1(n15821), .A2(n15301), .ZN(n27145));
    NOR2X1 U14274 (.A1(N4973), .A2(N11969), .ZN(n27146));
    INVX1 U14275 (.I(n23296), .ZN(n27147));
    INVX1 U14276 (.I(N8226), .ZN(N27148));
    NOR2X1 U14277 (.A1(N10677), .A2(n24645), .ZN(n27149));
    NOR2X1 U14278 (.A1(n17407), .A2(N1657), .ZN(N27150));
    NANDX1 U14279 (.A1(n15584), .A2(N9104), .ZN(n27151));
    NOR2X1 U14280 (.A1(N7968), .A2(N2055), .ZN(n27152));
    INVX1 U14281 (.I(N10819), .ZN(n27153));
    INVX1 U14282 (.I(n14166), .ZN(n27154));
    NOR2X1 U14283 (.A1(n21956), .A2(n15803), .ZN(n27155));
    INVX1 U14284 (.I(n24082), .ZN(n27156));
    NANDX1 U14285 (.A1(n19268), .A2(N2648), .ZN(n27157));
    NANDX1 U14286 (.A1(n24240), .A2(N3384), .ZN(N27158));
    NANDX1 U14287 (.A1(N10801), .A2(N12602), .ZN(N27159));
    NANDX1 U14288 (.A1(n14293), .A2(N12046), .ZN(n27160));
    INVX1 U14289 (.I(n24910), .ZN(n27161));
    NOR2X1 U14290 (.A1(N7397), .A2(N7417), .ZN(n27162));
    NANDX1 U14291 (.A1(N5268), .A2(N900), .ZN(n27163));
    NOR2X1 U14292 (.A1(N7322), .A2(n24014), .ZN(n27164));
    NANDX1 U14293 (.A1(n18327), .A2(N12677), .ZN(n27165));
    NANDX1 U14294 (.A1(N3548), .A2(n17247), .ZN(N27166));
    INVX1 U14295 (.I(n16397), .ZN(n27167));
    NOR2X1 U14296 (.A1(n17233), .A2(N7812), .ZN(n27168));
    INVX1 U14297 (.I(N4738), .ZN(N27169));
    NOR2X1 U14298 (.A1(N8436), .A2(n15538), .ZN(n27170));
    NANDX1 U14299 (.A1(n15034), .A2(N4329), .ZN(n27171));
    NANDX1 U14300 (.A1(N9542), .A2(n18006), .ZN(N27172));
    INVX1 U14301 (.I(N5706), .ZN(n27173));
    NANDX1 U14302 (.A1(N3165), .A2(N10973), .ZN(n27174));
    NANDX1 U14303 (.A1(N8201), .A2(n18294), .ZN(n27175));
    NANDX1 U14304 (.A1(N12824), .A2(n25389), .ZN(n27176));
    NOR2X1 U14305 (.A1(N7342), .A2(N3434), .ZN(n27177));
    NOR2X1 U14306 (.A1(N5307), .A2(N8599), .ZN(n27178));
    NANDX1 U14307 (.A1(N11307), .A2(n16410), .ZN(n27179));
    NOR2X1 U14308 (.A1(N4812), .A2(n16373), .ZN(N27180));
    NANDX1 U14309 (.A1(N9118), .A2(n17704), .ZN(n27181));
    NOR2X1 U14310 (.A1(N2214), .A2(N5579), .ZN(n27182));
    INVX1 U14311 (.I(n20219), .ZN(n27183));
    NANDX1 U14312 (.A1(N10541), .A2(n20139), .ZN(n27184));
    INVX1 U14313 (.I(n21513), .ZN(n27185));
    NANDX1 U14314 (.A1(N11807), .A2(N3073), .ZN(n27186));
    NOR2X1 U14315 (.A1(n13398), .A2(N2959), .ZN(N27187));
    NANDX1 U14316 (.A1(n20739), .A2(n20662), .ZN(N27188));
    INVX1 U14317 (.I(n14814), .ZN(N27189));
    NOR2X1 U14318 (.A1(n24231), .A2(n14888), .ZN(n27190));
    NOR2X1 U14319 (.A1(n21559), .A2(n19700), .ZN(n27191));
    NOR2X1 U14320 (.A1(n13053), .A2(n17585), .ZN(N27192));
    NOR2X1 U14321 (.A1(n22617), .A2(n19798), .ZN(N27193));
    INVX1 U14322 (.I(N1951), .ZN(N27194));
    NANDX1 U14323 (.A1(n23529), .A2(N12491), .ZN(N27195));
    NANDX1 U14324 (.A1(N1633), .A2(n22772), .ZN(n27196));
    INVX1 U14325 (.I(N2207), .ZN(n27197));
    NANDX1 U14326 (.A1(N11542), .A2(n15604), .ZN(N27198));
    NOR2X1 U14327 (.A1(N4983), .A2(n25110), .ZN(n27199));
    NANDX1 U14328 (.A1(n19483), .A2(N3189), .ZN(N27200));
    NANDX1 U14329 (.A1(n18211), .A2(n18077), .ZN(n27201));
    NANDX1 U14330 (.A1(N3035), .A2(N1042), .ZN(N27202));
    NANDX1 U14331 (.A1(N4855), .A2(n18626), .ZN(N27203));
    INVX1 U14332 (.I(N1970), .ZN(N27204));
    NOR2X1 U14333 (.A1(n17856), .A2(N3920), .ZN(n27205));
    NANDX1 U14334 (.A1(n15883), .A2(N5178), .ZN(n27206));
    NANDX1 U14335 (.A1(N6283), .A2(N2447), .ZN(n27207));
    NANDX1 U14336 (.A1(n22759), .A2(n17058), .ZN(N27208));
    NANDX1 U14337 (.A1(N1628), .A2(N9125), .ZN(n27209));
    INVX1 U14338 (.I(N1235), .ZN(n27210));
    NOR2X1 U14339 (.A1(N12840), .A2(N4424), .ZN(n27211));
    INVX1 U14340 (.I(n19818), .ZN(N27212));
    INVX1 U14341 (.I(N7601), .ZN(n27213));
    INVX1 U14342 (.I(N12309), .ZN(n27214));
    INVX1 U14343 (.I(N2205), .ZN(n27215));
    INVX1 U14344 (.I(n16363), .ZN(N27216));
    NOR2X1 U14345 (.A1(N7120), .A2(N8717), .ZN(n27217));
    INVX1 U14346 (.I(N12089), .ZN(n27218));
    NANDX1 U14347 (.A1(N2039), .A2(n14976), .ZN(n27219));
    NANDX1 U14348 (.A1(N4485), .A2(N3042), .ZN(n27220));
    NOR2X1 U14349 (.A1(N10311), .A2(n16919), .ZN(n27221));
    INVX1 U14350 (.I(N8203), .ZN(N27222));
    NANDX1 U14351 (.A1(N8534), .A2(N7592), .ZN(n27223));
    INVX1 U14352 (.I(N1725), .ZN(N27224));
    NOR2X1 U14353 (.A1(N6199), .A2(n12992), .ZN(n27225));
    NOR2X1 U14354 (.A1(N3549), .A2(n25300), .ZN(n27226));
    NOR2X1 U14355 (.A1(n20024), .A2(N5229), .ZN(N27227));
    NOR2X1 U14356 (.A1(n24197), .A2(N1116), .ZN(N27228));
    NOR2X1 U14357 (.A1(n21058), .A2(n13205), .ZN(n27229));
    INVX1 U14358 (.I(n23096), .ZN(N27230));
    NANDX1 U14359 (.A1(n14822), .A2(n16348), .ZN(n27231));
    NANDX1 U14360 (.A1(n20494), .A2(N1156), .ZN(n27232));
    INVX1 U14361 (.I(N2291), .ZN(N27233));
    NOR2X1 U14362 (.A1(n24719), .A2(n25094), .ZN(n27234));
    NANDX1 U14363 (.A1(N11100), .A2(N1317), .ZN(n27235));
    NOR2X1 U14364 (.A1(n17298), .A2(n14308), .ZN(n27236));
    NANDX1 U14365 (.A1(N9615), .A2(n14106), .ZN(n27237));
    NOR2X1 U14366 (.A1(N4136), .A2(N8102), .ZN(N27238));
    NANDX1 U14367 (.A1(N2830), .A2(n23488), .ZN(n27239));
    NANDX1 U14368 (.A1(N12655), .A2(N11190), .ZN(n27240));
    NANDX1 U14369 (.A1(N10248), .A2(N2635), .ZN(n27241));
    INVX1 U14370 (.I(N1094), .ZN(N27242));
    NOR2X1 U14371 (.A1(n16635), .A2(N2249), .ZN(N27243));
    NOR2X1 U14372 (.A1(n18925), .A2(N375), .ZN(N27244));
    NOR2X1 U14373 (.A1(n18516), .A2(n17325), .ZN(n27245));
    NOR2X1 U14374 (.A1(N8600), .A2(N9775), .ZN(N27246));
    NANDX1 U14375 (.A1(n22908), .A2(n25097), .ZN(n27247));
    INVX1 U14376 (.I(N279), .ZN(N27248));
    INVX1 U14377 (.I(n16192), .ZN(n27249));
    INVX1 U14378 (.I(n23952), .ZN(n27250));
    NOR2X1 U14379 (.A1(N6365), .A2(N10099), .ZN(N27251));
    NOR2X1 U14380 (.A1(N6322), .A2(n16921), .ZN(n27252));
    NANDX1 U14381 (.A1(N8957), .A2(n13062), .ZN(N27253));
    NOR2X1 U14382 (.A1(n20348), .A2(N4194), .ZN(N27254));
    NOR2X1 U14383 (.A1(n20679), .A2(N11886), .ZN(n27255));
    INVX1 U14384 (.I(N5957), .ZN(n27256));
    NOR2X1 U14385 (.A1(n18035), .A2(N2333), .ZN(n27257));
    INVX1 U14386 (.I(n16577), .ZN(N27258));
    INVX1 U14387 (.I(n13942), .ZN(n27259));
    NOR2X1 U14388 (.A1(n16831), .A2(n14220), .ZN(n27260));
    NOR2X1 U14389 (.A1(n21790), .A2(n22600), .ZN(n27261));
    NOR2X1 U14390 (.A1(N4077), .A2(n17732), .ZN(n27262));
    NOR2X1 U14391 (.A1(n13288), .A2(n24054), .ZN(N27263));
    NANDX1 U14392 (.A1(N7244), .A2(n21778), .ZN(n27264));
    NANDX1 U14393 (.A1(n16564), .A2(N5391), .ZN(n27265));
    NANDX1 U14394 (.A1(n16900), .A2(N567), .ZN(n27266));
    INVX1 U14395 (.I(N6378), .ZN(n27267));
    NOR2X1 U14396 (.A1(N2397), .A2(n24413), .ZN(n27268));
    NOR2X1 U14397 (.A1(N4664), .A2(N4255), .ZN(n27269));
    INVX1 U14398 (.I(n18605), .ZN(n27270));
    NOR2X1 U14399 (.A1(N7997), .A2(N7323), .ZN(n27271));
    NOR2X1 U14400 (.A1(n18554), .A2(n18690), .ZN(n27272));
    NOR2X1 U14401 (.A1(n22630), .A2(n25189), .ZN(N27273));
    NANDX1 U14402 (.A1(n24685), .A2(n23740), .ZN(n27274));
    INVX1 U14403 (.I(N6427), .ZN(n27275));
    NOR2X1 U14404 (.A1(N5003), .A2(N11758), .ZN(n27276));
    INVX1 U14405 (.I(n13079), .ZN(N27277));
    NOR2X1 U14406 (.A1(n14740), .A2(n21808), .ZN(n27278));
    INVX1 U14407 (.I(n21262), .ZN(n27279));
    NOR2X1 U14408 (.A1(N11480), .A2(N7653), .ZN(n27280));
    NANDX1 U14409 (.A1(n15735), .A2(n24321), .ZN(n27281));
    INVX1 U14410 (.I(N10658), .ZN(n27282));
    INVX1 U14411 (.I(n21098), .ZN(n27283));
    INVX1 U14412 (.I(n14136), .ZN(N27284));
    NANDX1 U14413 (.A1(n21602), .A2(N32), .ZN(n27285));
    INVX1 U14414 (.I(n23707), .ZN(n27286));
    INVX1 U14415 (.I(N977), .ZN(n27287));
    NOR2X1 U14416 (.A1(N5640), .A2(N9760), .ZN(n27288));
    NOR2X1 U14417 (.A1(N6165), .A2(N12700), .ZN(n27289));
    NOR2X1 U14418 (.A1(n23589), .A2(N1937), .ZN(n27290));
    NOR2X1 U14419 (.A1(N10657), .A2(N11967), .ZN(n27291));
    NANDX1 U14420 (.A1(n22136), .A2(n19619), .ZN(N27292));
    INVX1 U14421 (.I(N12368), .ZN(n27293));
    INVX1 U14422 (.I(N10126), .ZN(n27294));
    NANDX1 U14423 (.A1(N2787), .A2(N5722), .ZN(N27295));
    NOR2X1 U14424 (.A1(n16923), .A2(N8774), .ZN(n27296));
    NOR2X1 U14425 (.A1(N5722), .A2(N11513), .ZN(n27297));
    NOR2X1 U14426 (.A1(N4935), .A2(N1258), .ZN(n27298));
    NANDX1 U14427 (.A1(n24845), .A2(n25287), .ZN(N27299));
    NANDX1 U14428 (.A1(N5507), .A2(N12484), .ZN(n27300));
    NANDX1 U14429 (.A1(n17864), .A2(N3189), .ZN(n27301));
    NANDX1 U14430 (.A1(N3018), .A2(n15155), .ZN(N27302));
    NOR2X1 U14431 (.A1(n25153), .A2(n23541), .ZN(n27303));
    INVX1 U14432 (.I(N787), .ZN(n27304));
    NOR2X1 U14433 (.A1(N12173), .A2(N12580), .ZN(n27305));
    NOR2X1 U14434 (.A1(N6662), .A2(N3500), .ZN(N27306));
    INVX1 U14435 (.I(n15435), .ZN(N27307));
    INVX1 U14436 (.I(N8209), .ZN(n27308));
    NOR2X1 U14437 (.A1(N4284), .A2(N1912), .ZN(n27309));
    NOR2X1 U14438 (.A1(N6140), .A2(N1254), .ZN(n27310));
    NANDX1 U14439 (.A1(N1089), .A2(n21030), .ZN(N27311));
    INVX1 U14440 (.I(n19517), .ZN(N27312));
    NANDX1 U14441 (.A1(N9964), .A2(n17959), .ZN(N27313));
    NOR2X1 U14442 (.A1(n13886), .A2(N9385), .ZN(n27314));
    NANDX1 U14443 (.A1(N11925), .A2(N11432), .ZN(N27315));
    INVX1 U14444 (.I(n20206), .ZN(n27316));
    NANDX1 U14445 (.A1(n21230), .A2(n17003), .ZN(n27317));
    NOR2X1 U14446 (.A1(n24729), .A2(N8259), .ZN(n27318));
    NOR2X1 U14447 (.A1(n18287), .A2(N5235), .ZN(n27319));
    NOR2X1 U14448 (.A1(n22570), .A2(N7146), .ZN(n27320));
    NOR2X1 U14449 (.A1(N3207), .A2(n22669), .ZN(n27321));
    INVX1 U14450 (.I(n18565), .ZN(N27322));
    INVX1 U14451 (.I(n20256), .ZN(N27323));
    NANDX1 U14452 (.A1(N9123), .A2(N4717), .ZN(n27324));
    NOR2X1 U14453 (.A1(N3067), .A2(n18603), .ZN(n27325));
    NANDX1 U14454 (.A1(n22163), .A2(n19295), .ZN(N27326));
    NANDX1 U14455 (.A1(N5311), .A2(n13998), .ZN(n27327));
    NOR2X1 U14456 (.A1(N1038), .A2(n19768), .ZN(n27328));
    NOR2X1 U14457 (.A1(n14534), .A2(N2524), .ZN(n27329));
    INVX1 U14458 (.I(N7318), .ZN(N27330));
    INVX1 U14459 (.I(N1042), .ZN(n27331));
    INVX1 U14460 (.I(N3672), .ZN(n27332));
    NOR2X1 U14461 (.A1(N10630), .A2(N839), .ZN(N27333));
    INVX1 U14462 (.I(n17963), .ZN(n27334));
    NANDX1 U14463 (.A1(N5998), .A2(n19310), .ZN(N27335));
    INVX1 U14464 (.I(n24985), .ZN(n27336));
    INVX1 U14465 (.I(N8759), .ZN(n27337));
    NOR2X1 U14466 (.A1(n19338), .A2(N5419), .ZN(N27338));
    INVX1 U14467 (.I(N11493), .ZN(n27339));
    NANDX1 U14468 (.A1(n14642), .A2(N4786), .ZN(n27340));
    NOR2X1 U14469 (.A1(N8907), .A2(n17112), .ZN(N27341));
    INVX1 U14470 (.I(N199), .ZN(n27342));
    NANDX1 U14471 (.A1(n25423), .A2(N7957), .ZN(N27343));
    INVX1 U14472 (.I(N7344), .ZN(N27344));
    NANDX1 U14473 (.A1(N3512), .A2(n17974), .ZN(N27345));
    INVX1 U14474 (.I(N3525), .ZN(n27346));
    INVX1 U14475 (.I(n23306), .ZN(n27347));
    NOR2X1 U14476 (.A1(n18511), .A2(N3497), .ZN(N27348));
    INVX1 U14477 (.I(n20391), .ZN(n27349));
    NOR2X1 U14478 (.A1(N4624), .A2(n14226), .ZN(N27350));
    NOR2X1 U14479 (.A1(N5268), .A2(n14486), .ZN(N27351));
    NANDX1 U14480 (.A1(N8677), .A2(n19272), .ZN(N27352));
    NANDX1 U14481 (.A1(n17584), .A2(n25151), .ZN(n27353));
    NOR2X1 U14482 (.A1(N6550), .A2(N4354), .ZN(n27354));
    NOR2X1 U14483 (.A1(N3274), .A2(n24370), .ZN(n27355));
    INVX1 U14484 (.I(N3669), .ZN(N27356));
    INVX1 U14485 (.I(N4886), .ZN(n27357));
    NANDX1 U14486 (.A1(n20174), .A2(N4087), .ZN(n27358));
    INVX1 U14487 (.I(n18463), .ZN(N27359));
    NANDX1 U14488 (.A1(n23510), .A2(N5003), .ZN(n27360));
    NOR2X1 U14489 (.A1(n24533), .A2(N9626), .ZN(n27361));
    NOR2X1 U14490 (.A1(n19742), .A2(N3662), .ZN(n27362));
    INVX1 U14491 (.I(n14447), .ZN(N27363));
    NANDX1 U14492 (.A1(n17501), .A2(N12724), .ZN(N27364));
    NOR2X1 U14493 (.A1(N5917), .A2(N3604), .ZN(n27365));
    INVX1 U14494 (.I(n24540), .ZN(n27366));
    INVX1 U14495 (.I(N3009), .ZN(N27367));
    NOR2X1 U14496 (.A1(N6819), .A2(N6678), .ZN(n27368));
    NOR2X1 U14497 (.A1(N472), .A2(n14618), .ZN(n27369));
    NOR2X1 U14498 (.A1(N4558), .A2(n20361), .ZN(n27370));
    NOR2X1 U14499 (.A1(N1652), .A2(n18369), .ZN(N27371));
    INVX1 U14500 (.I(N7904), .ZN(N27372));
    NANDX1 U14501 (.A1(n22889), .A2(N2879), .ZN(n27373));
    NANDX1 U14502 (.A1(N1048), .A2(N1108), .ZN(n27374));
    INVX1 U14503 (.I(N2154), .ZN(N27375));
    NOR2X1 U14504 (.A1(n16344), .A2(n20842), .ZN(n27376));
    NANDX1 U14505 (.A1(n19947), .A2(n20578), .ZN(n27377));
    NANDX1 U14506 (.A1(N3119), .A2(n23586), .ZN(n27378));
    NANDX1 U14507 (.A1(n24207), .A2(n19031), .ZN(n27379));
    NANDX1 U14508 (.A1(n24678), .A2(N8146), .ZN(n27380));
    NOR2X1 U14509 (.A1(N3733), .A2(N3005), .ZN(N27381));
    NANDX1 U14510 (.A1(n19654), .A2(N10141), .ZN(n27382));
    NANDX1 U14511 (.A1(N2055), .A2(n16307), .ZN(N27383));
    NOR2X1 U14512 (.A1(n19204), .A2(N5480), .ZN(n27384));
    INVX1 U14513 (.I(N9079), .ZN(N27385));
    NOR2X1 U14514 (.A1(N3001), .A2(n16455), .ZN(N27386));
    NANDX1 U14515 (.A1(N12610), .A2(n18514), .ZN(n27387));
    NANDX1 U14516 (.A1(N7685), .A2(N5341), .ZN(N27388));
    INVX1 U14517 (.I(n20039), .ZN(n27389));
    NOR2X1 U14518 (.A1(n24748), .A2(N2335), .ZN(N27390));
    NANDX1 U14519 (.A1(N12691), .A2(N10481), .ZN(n27391));
    INVX1 U14520 (.I(n16424), .ZN(n27392));
    NANDX1 U14521 (.A1(n16475), .A2(n24845), .ZN(n27393));
    NANDX1 U14522 (.A1(N4618), .A2(n15668), .ZN(n27394));
    NOR2X1 U14523 (.A1(N4418), .A2(n23639), .ZN(N27395));
    NANDX1 U14524 (.A1(n19535), .A2(N7215), .ZN(n27396));
    INVX1 U14525 (.I(n22535), .ZN(n27397));
    INVX1 U14526 (.I(n23790), .ZN(N27398));
    NANDX1 U14527 (.A1(n16681), .A2(n21212), .ZN(n27399));
    NOR2X1 U14528 (.A1(N10789), .A2(n21752), .ZN(N27400));
    INVX1 U14529 (.I(n18168), .ZN(n27401));
    NANDX1 U14530 (.A1(n17235), .A2(N5405), .ZN(n27402));
    NANDX1 U14531 (.A1(n16483), .A2(N10266), .ZN(n27403));
    NOR2X1 U14532 (.A1(N7503), .A2(n15508), .ZN(n27404));
    INVX1 U14533 (.I(N8663), .ZN(n27405));
    INVX1 U14534 (.I(N5922), .ZN(n27406));
    NOR2X1 U14535 (.A1(n13311), .A2(N4058), .ZN(n27407));
    INVX1 U14536 (.I(N7343), .ZN(n27408));
    NANDX1 U14537 (.A1(N10688), .A2(n18645), .ZN(N27409));
    NOR2X1 U14538 (.A1(N8975), .A2(n17054), .ZN(N27410));
    NOR2X1 U14539 (.A1(N4684), .A2(N11916), .ZN(n27411));
    NOR2X1 U14540 (.A1(n15203), .A2(N1314), .ZN(n27412));
    INVX1 U14541 (.I(n13736), .ZN(n27413));
    INVX1 U14542 (.I(n15551), .ZN(N27414));
    INVX1 U14543 (.I(N12567), .ZN(N27415));
    NOR2X1 U14544 (.A1(N12833), .A2(n20070), .ZN(n27416));
    INVX1 U14545 (.I(N3087), .ZN(n27417));
    NANDX1 U14546 (.A1(n24714), .A2(N9009), .ZN(N27418));
    NOR2X1 U14547 (.A1(N12522), .A2(n13066), .ZN(n27419));
    NOR2X1 U14548 (.A1(N8632), .A2(n13106), .ZN(n27420));
    NOR2X1 U14549 (.A1(N1774), .A2(N11313), .ZN(n27421));
    NOR2X1 U14550 (.A1(N7596), .A2(n14967), .ZN(n27422));
    INVX1 U14551 (.I(n19511), .ZN(n27423));
    NOR2X1 U14552 (.A1(n13853), .A2(N9593), .ZN(N27424));
    INVX1 U14553 (.I(n16356), .ZN(n27425));
    NANDX1 U14554 (.A1(n18371), .A2(N1542), .ZN(n27426));
    NOR2X1 U14555 (.A1(n18684), .A2(N3142), .ZN(n27427));
    INVX1 U14556 (.I(N9003), .ZN(n27428));
    NANDX1 U14557 (.A1(N4808), .A2(n22484), .ZN(n27429));
    NOR2X1 U14558 (.A1(N11702), .A2(N9504), .ZN(N27430));
    NANDX1 U14559 (.A1(N8471), .A2(N6903), .ZN(n27431));
    INVX1 U14560 (.I(N4696), .ZN(N27432));
    NOR2X1 U14561 (.A1(n19023), .A2(N9894), .ZN(n27433));
    NANDX1 U14562 (.A1(N8488), .A2(N8544), .ZN(n27434));
    NOR2X1 U14563 (.A1(n15433), .A2(N11164), .ZN(N27435));
    NOR2X1 U14564 (.A1(n18253), .A2(N2017), .ZN(n27436));
    NANDX1 U14565 (.A1(N11122), .A2(n17828), .ZN(N27437));
    NANDX1 U14566 (.A1(n18573), .A2(N9737), .ZN(n27438));
    NOR2X1 U14567 (.A1(n16343), .A2(N4732), .ZN(n27439));
    NOR2X1 U14568 (.A1(n13325), .A2(n23006), .ZN(n27440));
    NANDX1 U14569 (.A1(N11596), .A2(N3341), .ZN(N27441));
    NOR2X1 U14570 (.A1(n18498), .A2(N11051), .ZN(n27442));
    NOR2X1 U14571 (.A1(n15942), .A2(N4572), .ZN(N27443));
    NOR2X1 U14572 (.A1(n20981), .A2(n13059), .ZN(n27444));
    INVX1 U14573 (.I(n20029), .ZN(n27445));
    NANDX1 U14574 (.A1(n22979), .A2(n17436), .ZN(N27446));
    INVX1 U14575 (.I(n13763), .ZN(N27447));
    NOR2X1 U14576 (.A1(N9898), .A2(n20358), .ZN(n27448));
    NANDX1 U14577 (.A1(N2969), .A2(N4592), .ZN(n27449));
    INVX1 U14578 (.I(N8079), .ZN(N27450));
    NOR2X1 U14579 (.A1(N4722), .A2(n21403), .ZN(N27451));
    NANDX1 U14580 (.A1(N7399), .A2(n21766), .ZN(n27452));
    NOR2X1 U14581 (.A1(N7315), .A2(n14762), .ZN(n27453));
    INVX1 U14582 (.I(n23158), .ZN(n27454));
    INVX1 U14583 (.I(n14556), .ZN(n27455));
    NANDX1 U14584 (.A1(N680), .A2(n16382), .ZN(n27456));
    NOR2X1 U14585 (.A1(N9476), .A2(N8138), .ZN(N27457));
    NANDX1 U14586 (.A1(N1409), .A2(N6915), .ZN(N27458));
    NOR2X1 U14587 (.A1(N10696), .A2(n16812), .ZN(n27459));
    INVX1 U14588 (.I(n15807), .ZN(N27460));
    INVX1 U14589 (.I(N966), .ZN(N27461));
    NANDX1 U14590 (.A1(n16627), .A2(N10289), .ZN(n27462));
    NOR2X1 U14591 (.A1(N1295), .A2(N5883), .ZN(n27463));
    NOR2X1 U14592 (.A1(n23061), .A2(N4817), .ZN(n27464));
    NOR2X1 U14593 (.A1(N12320), .A2(n14802), .ZN(n27465));
    NANDX1 U14594 (.A1(N6288), .A2(n18125), .ZN(N27466));
    INVX1 U14595 (.I(n21237), .ZN(n27467));
    NANDX1 U14596 (.A1(n15385), .A2(n19480), .ZN(N27468));
    NANDX1 U14597 (.A1(n14373), .A2(n20889), .ZN(N27469));
    NOR2X1 U14598 (.A1(N1621), .A2(n20352), .ZN(N27470));
    NANDX1 U14599 (.A1(n23497), .A2(N10657), .ZN(N27471));
    NANDX1 U14600 (.A1(n24463), .A2(n17744), .ZN(n27472));
    INVX1 U14601 (.I(n23519), .ZN(n27473));
    NOR2X1 U14602 (.A1(N8138), .A2(n18170), .ZN(n27474));
    NOR2X1 U14603 (.A1(N5696), .A2(n22986), .ZN(N27475));
    NANDX1 U14604 (.A1(N6783), .A2(N1053), .ZN(N27476));
    NANDX1 U14605 (.A1(N1838), .A2(N7946), .ZN(n27477));
    NANDX1 U14606 (.A1(N11843), .A2(N5718), .ZN(n27478));
    NANDX1 U14607 (.A1(N5820), .A2(N11627), .ZN(n27479));
    NANDX1 U14608 (.A1(N1206), .A2(n13219), .ZN(n27480));
    NANDX1 U14609 (.A1(N10326), .A2(N6120), .ZN(N27481));
    INVX1 U14610 (.I(n20982), .ZN(n27482));
    NOR2X1 U14611 (.A1(N3837), .A2(N1991), .ZN(n27483));
    NANDX1 U14612 (.A1(n16124), .A2(n20310), .ZN(n27484));
    INVX1 U14613 (.I(N8791), .ZN(N27485));
    NOR2X1 U14614 (.A1(n17011), .A2(n20544), .ZN(n27486));
    NOR2X1 U14615 (.A1(n23793), .A2(N10365), .ZN(N27487));
    INVX1 U14616 (.I(n14398), .ZN(n27488));
    NANDX1 U14617 (.A1(N4978), .A2(N738), .ZN(n27489));
    NOR2X1 U14618 (.A1(n18332), .A2(N6558), .ZN(N27490));
    NOR2X1 U14619 (.A1(n20555), .A2(n22033), .ZN(N27491));
    NOR2X1 U14620 (.A1(n13167), .A2(N6856), .ZN(n27492));
    INVX1 U14621 (.I(N3774), .ZN(N27493));
    INVX1 U14622 (.I(N322), .ZN(N27494));
    NOR2X1 U14623 (.A1(n18595), .A2(N3500), .ZN(N27495));
    NOR2X1 U14624 (.A1(n13402), .A2(n14815), .ZN(n27496));
    INVX1 U14625 (.I(n23271), .ZN(N27497));
    NANDX1 U14626 (.A1(n19371), .A2(n23718), .ZN(n27498));
    NANDX1 U14627 (.A1(N4233), .A2(n19494), .ZN(n27499));
    NOR2X1 U14628 (.A1(N11310), .A2(n24471), .ZN(n27500));
    NOR2X1 U14629 (.A1(N9834), .A2(n17300), .ZN(n27501));
    NOR2X1 U14630 (.A1(n23022), .A2(N12353), .ZN(N27502));
    NANDX1 U14631 (.A1(N9657), .A2(N17), .ZN(n27503));
    INVX1 U14632 (.I(n16680), .ZN(N27504));
    NANDX1 U14633 (.A1(n15637), .A2(N5769), .ZN(N27505));
    NOR2X1 U14634 (.A1(N8730), .A2(N9268), .ZN(n27506));
    NOR2X1 U14635 (.A1(N10899), .A2(n24082), .ZN(n27507));
    INVX1 U14636 (.I(N8667), .ZN(n27508));
    NANDX1 U14637 (.A1(n22671), .A2(n21152), .ZN(n27509));
    INVX1 U14638 (.I(N1401), .ZN(n27510));
    INVX1 U14639 (.I(n23368), .ZN(n27511));
    NANDX1 U14640 (.A1(n14112), .A2(n20651), .ZN(n27512));
    INVX1 U14641 (.I(n20179), .ZN(n27513));
    NANDX1 U14642 (.A1(N8830), .A2(N7029), .ZN(n27514));
    INVX1 U14643 (.I(N7254), .ZN(n27515));
    NANDX1 U14644 (.A1(n15699), .A2(n23934), .ZN(n27516));
    INVX1 U14645 (.I(N5834), .ZN(n27517));
    INVX1 U14646 (.I(n20116), .ZN(n27518));
    INVX1 U14647 (.I(n13468), .ZN(n27519));
    INVX1 U14648 (.I(N2997), .ZN(n27520));
    INVX1 U14649 (.I(N2388), .ZN(n27521));
    NANDX1 U14650 (.A1(N8755), .A2(n25058), .ZN(n27522));
    INVX1 U14651 (.I(N10074), .ZN(n27523));
    NOR2X1 U14652 (.A1(n25494), .A2(N7939), .ZN(n27524));
    NANDX1 U14653 (.A1(N2871), .A2(n17357), .ZN(n27525));
    NANDX1 U14654 (.A1(n23049), .A2(N5113), .ZN(n27526));
    INVX1 U14655 (.I(n18846), .ZN(n27527));
    INVX1 U14656 (.I(n18594), .ZN(n27528));
    NANDX1 U14657 (.A1(n15014), .A2(n17025), .ZN(N27529));
    NOR2X1 U14658 (.A1(N9615), .A2(n21224), .ZN(N27530));
    INVX1 U14659 (.I(N1713), .ZN(N27531));
    NANDX1 U14660 (.A1(N2806), .A2(N4710), .ZN(n27532));
    INVX1 U14661 (.I(n19463), .ZN(n27533));
    NOR2X1 U14662 (.A1(N7526), .A2(n19018), .ZN(n27534));
    NOR2X1 U14663 (.A1(n17599), .A2(N8741), .ZN(n27535));
    NOR2X1 U14664 (.A1(N36), .A2(N11173), .ZN(n27536));
    NANDX1 U14665 (.A1(n17392), .A2(n13683), .ZN(n27537));
    NOR2X1 U14666 (.A1(N11273), .A2(n25022), .ZN(n27538));
    NOR2X1 U14667 (.A1(N10588), .A2(n18113), .ZN(N27539));
    NANDX1 U14668 (.A1(n14369), .A2(N9635), .ZN(n27540));
    INVX1 U14669 (.I(n23984), .ZN(n27541));
    NANDX1 U14670 (.A1(N6064), .A2(N194), .ZN(N27542));
    INVX1 U14671 (.I(N8869), .ZN(n27543));
    NOR2X1 U14672 (.A1(n16354), .A2(N2829), .ZN(n27544));
    NANDX1 U14673 (.A1(n23879), .A2(N10614), .ZN(n27545));
    NOR2X1 U14674 (.A1(N4744), .A2(n19354), .ZN(n27546));
    NANDX1 U14675 (.A1(n19049), .A2(n19294), .ZN(n27547));
    NANDX1 U14676 (.A1(n25208), .A2(n21744), .ZN(N27548));
    INVX1 U14677 (.I(n25248), .ZN(n27549));
    NOR2X1 U14678 (.A1(N3764), .A2(N10333), .ZN(N27550));
    INVX1 U14679 (.I(N11275), .ZN(N27551));
    INVX1 U14680 (.I(N1045), .ZN(n27552));
    NANDX1 U14681 (.A1(N11951), .A2(n20671), .ZN(n27553));
    INVX1 U14682 (.I(N912), .ZN(n27554));
    NANDX1 U14683 (.A1(N6088), .A2(n20085), .ZN(N27555));
    INVX1 U14684 (.I(n23187), .ZN(n27556));
    NANDX1 U14685 (.A1(N1979), .A2(N8298), .ZN(n27557));
    INVX1 U14686 (.I(n20992), .ZN(n27558));
    INVX1 U14687 (.I(n24127), .ZN(N27559));
    NANDX1 U14688 (.A1(n24481), .A2(N4869), .ZN(n27560));
    INVX1 U14689 (.I(n20723), .ZN(n27561));
    NANDX1 U14690 (.A1(n13989), .A2(N5252), .ZN(n27562));
    NANDX1 U14691 (.A1(n13090), .A2(n22163), .ZN(N27563));
    NOR2X1 U14692 (.A1(N1057), .A2(n23207), .ZN(n27564));
    INVX1 U14693 (.I(N1775), .ZN(n27565));
    INVX1 U14694 (.I(n22228), .ZN(n27566));
    NANDX1 U14695 (.A1(n19894), .A2(n17084), .ZN(n27567));
    NANDX1 U14696 (.A1(n23496), .A2(n14768), .ZN(N27568));
    INVX1 U14697 (.I(n14242), .ZN(N27569));
    NANDX1 U14698 (.A1(n21738), .A2(n24002), .ZN(N27570));
    NANDX1 U14699 (.A1(n20362), .A2(n13037), .ZN(n27571));
    NOR2X1 U14700 (.A1(n13998), .A2(N1778), .ZN(n27572));
    NANDX1 U14701 (.A1(N7312), .A2(n15767), .ZN(n27573));
    NOR2X1 U14702 (.A1(N7427), .A2(n17624), .ZN(n27574));
    NANDX1 U14703 (.A1(n18816), .A2(n18680), .ZN(n27575));
    NANDX1 U14704 (.A1(N7091), .A2(n20454), .ZN(N27576));
    NOR2X1 U14705 (.A1(n18086), .A2(n23139), .ZN(n27577));
    NANDX1 U14706 (.A1(N9667), .A2(n23445), .ZN(n27578));
    NANDX1 U14707 (.A1(n24434), .A2(N5911), .ZN(N27579));
    NANDX1 U14708 (.A1(n21997), .A2(N2146), .ZN(N27580));
    INVX1 U14709 (.I(n24746), .ZN(n27581));
    INVX1 U14710 (.I(n16712), .ZN(n27582));
    INVX1 U14711 (.I(n25273), .ZN(n27583));
    NOR2X1 U14712 (.A1(N12190), .A2(n21353), .ZN(n27584));
    NANDX1 U14713 (.A1(N3157), .A2(n17547), .ZN(n27585));
    NANDX1 U14714 (.A1(N5055), .A2(N10861), .ZN(N27586));
    NOR2X1 U14715 (.A1(n18927), .A2(N6719), .ZN(N27587));
    INVX1 U14716 (.I(N3207), .ZN(n27588));
    INVX1 U14717 (.I(n18217), .ZN(n27589));
    NOR2X1 U14718 (.A1(n23239), .A2(n16159), .ZN(N27590));
    INVX1 U14719 (.I(n22170), .ZN(N27591));
    NOR2X1 U14720 (.A1(N3491), .A2(N7432), .ZN(n27592));
    NOR2X1 U14721 (.A1(n21436), .A2(n20946), .ZN(n27593));
    NOR2X1 U14722 (.A1(N1414), .A2(n21917), .ZN(n27594));
    NOR2X1 U14723 (.A1(N8671), .A2(n22875), .ZN(n27595));
    NANDX1 U14724 (.A1(N9230), .A2(n14799), .ZN(n27596));
    INVX1 U14725 (.I(n13142), .ZN(n27597));
    NANDX1 U14726 (.A1(N3357), .A2(n24501), .ZN(n27598));
    NANDX1 U14727 (.A1(N10075), .A2(n19579), .ZN(n27599));
    NANDX1 U14728 (.A1(N9376), .A2(N12293), .ZN(n27600));
    INVX1 U14729 (.I(N7112), .ZN(n27601));
    INVX1 U14730 (.I(N10946), .ZN(n27602));
    NANDX1 U14731 (.A1(N2554), .A2(N3205), .ZN(N27603));
    NANDX1 U14732 (.A1(N4304), .A2(n24640), .ZN(n27604));
    NOR2X1 U14733 (.A1(N6097), .A2(n14821), .ZN(n27605));
    NOR2X1 U14734 (.A1(N7661), .A2(n23491), .ZN(n27606));
    NANDX1 U14735 (.A1(N8112), .A2(n21488), .ZN(n27607));
    NOR2X1 U14736 (.A1(N11840), .A2(N9127), .ZN(n27608));
    NOR2X1 U14737 (.A1(N3964), .A2(n22395), .ZN(n27609));
    NANDX1 U14738 (.A1(n14038), .A2(N5239), .ZN(n27610));
    INVX1 U14739 (.I(N12182), .ZN(N27611));
    INVX1 U14740 (.I(n13128), .ZN(N27612));
    INVX1 U14741 (.I(N9249), .ZN(N27613));
    INVX1 U14742 (.I(N608), .ZN(N27614));
    INVX1 U14743 (.I(N4814), .ZN(n27615));
    INVX1 U14744 (.I(N4874), .ZN(n27616));
    NOR2X1 U14745 (.A1(n13316), .A2(N10970), .ZN(n27617));
    NOR2X1 U14746 (.A1(N8190), .A2(N7398), .ZN(N27618));
    INVX1 U14747 (.I(N436), .ZN(n27619));
    INVX1 U14748 (.I(N1514), .ZN(n27620));
    NANDX1 U14749 (.A1(n16117), .A2(n24910), .ZN(n27621));
    NANDX1 U14750 (.A1(n20081), .A2(N10571), .ZN(N27622));
    NOR2X1 U14751 (.A1(n22886), .A2(n15809), .ZN(n27623));
    INVX1 U14752 (.I(N9565), .ZN(n27624));
    NANDX1 U14753 (.A1(N9551), .A2(N6394), .ZN(n27625));
    NOR2X1 U14754 (.A1(n22392), .A2(N7001), .ZN(N27626));
    INVX1 U14755 (.I(n15973), .ZN(N27627));
    INVX1 U14756 (.I(N65), .ZN(N27628));
    NOR2X1 U14757 (.A1(N12709), .A2(n25304), .ZN(N27629));
    NOR2X1 U14758 (.A1(n20898), .A2(N7200), .ZN(N27630));
    INVX1 U14759 (.I(N10102), .ZN(n27631));
    INVX1 U14760 (.I(N12039), .ZN(N27632));
    NANDX1 U14761 (.A1(N2091), .A2(N215), .ZN(N27633));
    NOR2X1 U14762 (.A1(n22171), .A2(n25055), .ZN(n27634));
    NOR2X1 U14763 (.A1(N8323), .A2(N4129), .ZN(N27635));
    NOR2X1 U14764 (.A1(n17887), .A2(N735), .ZN(N27636));
    NANDX1 U14765 (.A1(n24280), .A2(n20858), .ZN(n27637));
    INVX1 U14766 (.I(n20049), .ZN(n27638));
    NANDX1 U14767 (.A1(n21793), .A2(n19441), .ZN(n27639));
    NANDX1 U14768 (.A1(N4982), .A2(N6647), .ZN(n27640));
    NOR2X1 U14769 (.A1(n21212), .A2(n16313), .ZN(n27641));
    INVX1 U14770 (.I(N6235), .ZN(n27642));
    NOR2X1 U14771 (.A1(N894), .A2(N7042), .ZN(n27643));
    NANDX1 U14772 (.A1(N2984), .A2(N7256), .ZN(n27644));
    NANDX1 U14773 (.A1(n13923), .A2(n21078), .ZN(n27645));
    INVX1 U14774 (.I(n22245), .ZN(N27646));
    NOR2X1 U14775 (.A1(n19665), .A2(N3397), .ZN(N27647));
    NANDX1 U14776 (.A1(n14325), .A2(n16445), .ZN(N27648));
    NOR2X1 U14777 (.A1(N8912), .A2(N10991), .ZN(N27649));
    NANDX1 U14778 (.A1(n19472), .A2(n19199), .ZN(N27650));
    INVX1 U14779 (.I(n13221), .ZN(n27651));
    NANDX1 U14780 (.A1(N5017), .A2(N8930), .ZN(n27652));
    INVX1 U14781 (.I(n19936), .ZN(N27653));
    NOR2X1 U14782 (.A1(N6335), .A2(n20829), .ZN(N27654));
    NOR2X1 U14783 (.A1(N2363), .A2(N12580), .ZN(N27655));
    NANDX1 U14784 (.A1(N8459), .A2(N1000), .ZN(n27656));
    NANDX1 U14785 (.A1(N3241), .A2(N12012), .ZN(n27657));
    INVX1 U14786 (.I(n22905), .ZN(n27658));
    NANDX1 U14787 (.A1(N5751), .A2(N495), .ZN(n27659));
    NOR2X1 U14788 (.A1(n15814), .A2(n23677), .ZN(N27660));
    INVX1 U14789 (.I(N8229), .ZN(n27661));
    NANDX1 U14790 (.A1(n25307), .A2(n19795), .ZN(N27662));
    NANDX1 U14791 (.A1(n14418), .A2(n24811), .ZN(n27663));
    NANDX1 U14792 (.A1(n19841), .A2(n19244), .ZN(N27664));
    INVX1 U14793 (.I(N673), .ZN(N27665));
    NANDX1 U14794 (.A1(N6735), .A2(n17305), .ZN(n27666));
    NANDX1 U14795 (.A1(n13731), .A2(N261), .ZN(n27667));
    INVX1 U14796 (.I(n16302), .ZN(n27668));
    NOR2X1 U14797 (.A1(N6465), .A2(N7345), .ZN(n27669));
    NANDX1 U14798 (.A1(n21873), .A2(n13095), .ZN(n27670));
    NANDX1 U14799 (.A1(n16991), .A2(n17676), .ZN(N27671));
    NANDX1 U14800 (.A1(n23099), .A2(n14672), .ZN(N27672));
    NOR2X1 U14801 (.A1(N11671), .A2(N8965), .ZN(n27673));
    NANDX1 U14802 (.A1(N587), .A2(N8273), .ZN(n27674));
    INVX1 U14803 (.I(N9195), .ZN(N27675));
    INVX1 U14804 (.I(N1979), .ZN(N27676));
    NANDX1 U14805 (.A1(N8390), .A2(N8714), .ZN(n27677));
    NOR2X1 U14806 (.A1(n13075), .A2(N11212), .ZN(n27678));
    INVX1 U14807 (.I(n18760), .ZN(n27679));
    NOR2X1 U14808 (.A1(N11508), .A2(n13992), .ZN(n27680));
    INVX1 U14809 (.I(n15449), .ZN(N27681));
    INVX1 U14810 (.I(n25488), .ZN(N27682));
    NOR2X1 U14811 (.A1(N1850), .A2(N6429), .ZN(n27683));
    NANDX1 U14812 (.A1(n13716), .A2(n21100), .ZN(n27684));
    NANDX1 U14813 (.A1(n25386), .A2(n18832), .ZN(N27685));
    INVX1 U14814 (.I(n14740), .ZN(N27686));
    NOR2X1 U14815 (.A1(N10233), .A2(n23935), .ZN(n27687));
    INVX1 U14816 (.I(N12212), .ZN(n27688));
    NANDX1 U14817 (.A1(n15044), .A2(N9693), .ZN(N27689));
    INVX1 U14818 (.I(N2617), .ZN(n27690));
    NANDX1 U14819 (.A1(N9781), .A2(N10144), .ZN(n27691));
    INVX1 U14820 (.I(N10056), .ZN(n27692));
    NOR2X1 U14821 (.A1(n24076), .A2(N3), .ZN(N27693));
    INVX1 U14822 (.I(N12829), .ZN(n27694));
    NANDX1 U14823 (.A1(n13881), .A2(n19257), .ZN(n27695));
    NANDX1 U14824 (.A1(N2094), .A2(N3623), .ZN(n27696));
    INVX1 U14825 (.I(n16247), .ZN(n27697));
    NANDX1 U14826 (.A1(N2329), .A2(N5485), .ZN(n27698));
    NANDX1 U14827 (.A1(N12562), .A2(n18187), .ZN(N27699));
    NOR2X1 U14828 (.A1(n13541), .A2(n18292), .ZN(n27700));
    NOR2X1 U14829 (.A1(n23233), .A2(N8834), .ZN(N27701));
    NANDX1 U14830 (.A1(n18634), .A2(n18615), .ZN(n27702));
    INVX1 U14831 (.I(n19085), .ZN(n27703));
    NANDX1 U14832 (.A1(N985), .A2(n17658), .ZN(N27704));
    INVX1 U14833 (.I(n13016), .ZN(n27705));
    INVX1 U14834 (.I(N3631), .ZN(n27706));
    NANDX1 U14835 (.A1(n13009), .A2(N4122), .ZN(n27707));
    NANDX1 U14836 (.A1(N5399), .A2(n16705), .ZN(N27708));
    NANDX1 U14837 (.A1(n16621), .A2(N7801), .ZN(n27709));
    INVX1 U14838 (.I(n18212), .ZN(n27710));
    NANDX1 U14839 (.A1(n20939), .A2(N956), .ZN(N27711));
    NANDX1 U14840 (.A1(n13728), .A2(n13013), .ZN(n27712));
    NOR2X1 U14841 (.A1(N11330), .A2(n16454), .ZN(N27713));
    NANDX1 U14842 (.A1(n18712), .A2(N4536), .ZN(n27714));
    NOR2X1 U14843 (.A1(N10647), .A2(n19790), .ZN(n27715));
    INVX1 U14844 (.I(n16855), .ZN(N27716));
    NANDX1 U14845 (.A1(N7291), .A2(N9253), .ZN(n27717));
    NOR2X1 U14846 (.A1(N9068), .A2(n13374), .ZN(n27718));
    INVX1 U14847 (.I(n14466), .ZN(N27719));
    NOR2X1 U14848 (.A1(N12488), .A2(N5584), .ZN(N27720));
    NOR2X1 U14849 (.A1(n15241), .A2(n23796), .ZN(N27721));
    NANDX1 U14850 (.A1(n24947), .A2(n24751), .ZN(N27722));
    INVX1 U14851 (.I(N1941), .ZN(n27723));
    NOR2X1 U14852 (.A1(N2339), .A2(n13270), .ZN(n27724));
    INVX1 U14853 (.I(N4638), .ZN(n27725));
    INVX1 U14854 (.I(N10785), .ZN(n27726));
    NANDX1 U14855 (.A1(N5893), .A2(N5072), .ZN(n27727));
    NOR2X1 U14856 (.A1(n22747), .A2(N1142), .ZN(N27728));
    NOR2X1 U14857 (.A1(N6497), .A2(n12875), .ZN(N27729));
    NOR2X1 U14858 (.A1(N8638), .A2(n16862), .ZN(n27730));
    NOR2X1 U14859 (.A1(n16251), .A2(N3847), .ZN(N27731));
    NANDX1 U14860 (.A1(N6163), .A2(N7855), .ZN(n27732));
    NOR2X1 U14861 (.A1(N5204), .A2(n21570), .ZN(N27733));
    NANDX1 U14862 (.A1(N1412), .A2(n23510), .ZN(n27734));
    NANDX1 U14863 (.A1(N3750), .A2(N45), .ZN(N27735));
    NANDX1 U14864 (.A1(n22657), .A2(N9561), .ZN(n27736));
    INVX1 U14865 (.I(N11943), .ZN(n27737));
    INVX1 U14866 (.I(n14977), .ZN(N27738));
    INVX1 U14867 (.I(N1466), .ZN(n27739));
    NANDX1 U14868 (.A1(N2419), .A2(n22232), .ZN(n27740));
    NANDX1 U14869 (.A1(n24639), .A2(n19638), .ZN(n27741));
    NANDX1 U14870 (.A1(n21552), .A2(n24656), .ZN(n27742));
    NANDX1 U14871 (.A1(N1585), .A2(n19586), .ZN(n27743));
    INVX1 U14872 (.I(N5413), .ZN(N27744));
    NOR2X1 U14873 (.A1(n19925), .A2(n22759), .ZN(n27745));
    NANDX1 U14874 (.A1(N6700), .A2(n15631), .ZN(n27746));
    NOR2X1 U14875 (.A1(n21014), .A2(N482), .ZN(n27747));
    INVX1 U14876 (.I(N5072), .ZN(N27748));
    INVX1 U14877 (.I(N5351), .ZN(n27749));
    NOR2X1 U14878 (.A1(N11093), .A2(N8886), .ZN(n27750));
    NANDX1 U14879 (.A1(n15978), .A2(N72), .ZN(N27751));
    NOR2X1 U14880 (.A1(N8235), .A2(n24710), .ZN(N27752));
    NANDX1 U14881 (.A1(N6121), .A2(N9528), .ZN(n27753));
    INVX1 U14882 (.I(n22124), .ZN(n27754));
    INVX1 U14883 (.I(n23399), .ZN(n27755));
    NANDX1 U14884 (.A1(N5293), .A2(N11453), .ZN(N27756));
    INVX1 U14885 (.I(N2549), .ZN(N27757));
    NOR2X1 U14886 (.A1(N10368), .A2(n18180), .ZN(n27758));
    NOR2X1 U14887 (.A1(N5879), .A2(N7429), .ZN(n27759));
    INVX1 U14888 (.I(n25220), .ZN(n27760));
    NANDX1 U14889 (.A1(N7163), .A2(N9009), .ZN(n27761));
    INVX1 U14890 (.I(N4817), .ZN(N27762));
    INVX1 U14891 (.I(N8152), .ZN(n27763));
    NOR2X1 U14892 (.A1(N4788), .A2(N5154), .ZN(N27764));
    INVX1 U14893 (.I(n23717), .ZN(n27765));
    NOR2X1 U14894 (.A1(n16661), .A2(N2027), .ZN(n27766));
    INVX1 U14895 (.I(n16540), .ZN(n27767));
    INVX1 U14896 (.I(n17142), .ZN(n27768));
    INVX1 U14897 (.I(N144), .ZN(N27769));
    NOR2X1 U14898 (.A1(n13149), .A2(n15332), .ZN(N27770));
    NANDX1 U14899 (.A1(n20096), .A2(n23736), .ZN(n27771));
    NANDX1 U14900 (.A1(n16292), .A2(n14316), .ZN(n27772));
    NOR2X1 U14901 (.A1(N8605), .A2(n21479), .ZN(n27773));
    INVX1 U14902 (.I(N779), .ZN(n27774));
    INVX1 U14903 (.I(N6347), .ZN(N27775));
    NOR2X1 U14904 (.A1(N8718), .A2(n25404), .ZN(n27776));
    NOR2X1 U14905 (.A1(N1581), .A2(n23618), .ZN(n27777));
    NOR2X1 U14906 (.A1(N7009), .A2(N143), .ZN(N27778));
    INVX1 U14907 (.I(n23549), .ZN(n27779));
    NANDX1 U14908 (.A1(n16697), .A2(N8646), .ZN(N27780));
    INVX1 U14909 (.I(N12004), .ZN(n27781));
    NANDX1 U14910 (.A1(N7346), .A2(N6446), .ZN(n27782));
    INVX1 U14911 (.I(n19849), .ZN(N27783));
    INVX1 U14912 (.I(n21447), .ZN(n27784));
    INVX1 U14913 (.I(N9841), .ZN(n27785));
    INVX1 U14914 (.I(n18909), .ZN(N27786));
    NANDX1 U14915 (.A1(n19597), .A2(N8469), .ZN(N27787));
    NANDX1 U14916 (.A1(N3024), .A2(n17186), .ZN(N27788));
    INVX1 U14917 (.I(N5875), .ZN(N27789));
    INVX1 U14918 (.I(N786), .ZN(N27790));
    INVX1 U14919 (.I(n14543), .ZN(n27791));
    NOR2X1 U14920 (.A1(N8323), .A2(N1357), .ZN(N27792));
    NANDX1 U14921 (.A1(n25019), .A2(N10003), .ZN(n27793));
    NOR2X1 U14922 (.A1(N11521), .A2(N9332), .ZN(N27794));
    INVX1 U14923 (.I(N6734), .ZN(n27795));
    NOR2X1 U14924 (.A1(N12006), .A2(N2268), .ZN(n27796));
    INVX1 U14925 (.I(N9436), .ZN(n27797));
    NOR2X1 U14926 (.A1(n18017), .A2(N2842), .ZN(N27798));
    INVX1 U14927 (.I(N12112), .ZN(n27799));
    NOR2X1 U14928 (.A1(n22531), .A2(n15135), .ZN(n27800));
    INVX1 U14929 (.I(n25201), .ZN(n27801));
    NOR2X1 U14930 (.A1(n13565), .A2(N484), .ZN(n27802));
    INVX1 U14931 (.I(n16876), .ZN(n27803));
    NOR2X1 U14932 (.A1(n15634), .A2(n18232), .ZN(N27804));
    INVX1 U14933 (.I(n15150), .ZN(N27805));
    NOR2X1 U14934 (.A1(N7561), .A2(N1168), .ZN(n27806));
    NOR2X1 U14935 (.A1(n13988), .A2(n22172), .ZN(N27807));
    NANDX1 U14936 (.A1(N491), .A2(n24439), .ZN(n27808));
    NOR2X1 U14937 (.A1(N9926), .A2(n25314), .ZN(N27809));
    INVX1 U14938 (.I(N1535), .ZN(n27810));
    NOR2X1 U14939 (.A1(n22179), .A2(N1612), .ZN(N27811));
    NOR2X1 U14940 (.A1(N580), .A2(N7642), .ZN(n27812));
    INVX1 U14941 (.I(n24626), .ZN(N27813));
    NOR2X1 U14942 (.A1(N8589), .A2(N6435), .ZN(n27814));
    INVX1 U14943 (.I(n13038), .ZN(n27815));
    INVX1 U14944 (.I(N8347), .ZN(n27816));
    NANDX1 U14945 (.A1(N11716), .A2(n14117), .ZN(n27817));
    NOR2X1 U14946 (.A1(N1651), .A2(N3716), .ZN(N27818));
    INVX1 U14947 (.I(n23822), .ZN(n27819));
    NOR2X1 U14948 (.A1(N9859), .A2(N11526), .ZN(n27820));
    NANDX1 U14949 (.A1(n19784), .A2(N11338), .ZN(n27821));
    NANDX1 U14950 (.A1(N10086), .A2(n19679), .ZN(n27822));
    NOR2X1 U14951 (.A1(N11697), .A2(n25048), .ZN(n27823));
    NOR2X1 U14952 (.A1(N8106), .A2(N7651), .ZN(n27824));
    NANDX1 U14953 (.A1(n18080), .A2(n16239), .ZN(n27825));
    NOR2X1 U14954 (.A1(n19427), .A2(N3775), .ZN(n27826));
    INVX1 U14955 (.I(n16542), .ZN(n27827));
    NANDX1 U14956 (.A1(N1587), .A2(n19426), .ZN(N27828));
    INVX1 U14957 (.I(n17508), .ZN(N27829));
    NOR2X1 U14958 (.A1(n18808), .A2(n15827), .ZN(N27830));
    NOR2X1 U14959 (.A1(N3164), .A2(N1851), .ZN(n27831));
    INVX1 U14960 (.I(N11715), .ZN(n27832));
    INVX1 U14961 (.I(N10052), .ZN(N27833));
    NANDX1 U14962 (.A1(n21634), .A2(N8453), .ZN(n27834));
    NANDX1 U14963 (.A1(N9947), .A2(N7433), .ZN(N27835));
    NANDX1 U14964 (.A1(n17597), .A2(n19807), .ZN(n27836));
    NOR2X1 U14965 (.A1(N8333), .A2(n13113), .ZN(N27837));
    NOR2X1 U14966 (.A1(N875), .A2(N2984), .ZN(n27838));
    INVX1 U14967 (.I(N3702), .ZN(n27839));
    INVX1 U14968 (.I(N4872), .ZN(n27840));
    INVX1 U14969 (.I(N10846), .ZN(N27841));
    NOR2X1 U14970 (.A1(n20717), .A2(n15440), .ZN(N27842));
    NANDX1 U14971 (.A1(n23880), .A2(n17290), .ZN(n27843));
    NANDX1 U14972 (.A1(n24363), .A2(N8013), .ZN(N27844));
    NANDX1 U14973 (.A1(n20660), .A2(N4144), .ZN(n27845));
    NANDX1 U14974 (.A1(N6190), .A2(N2858), .ZN(n27846));
    INVX1 U14975 (.I(N11057), .ZN(n27847));
    NOR2X1 U14976 (.A1(n20127), .A2(n22771), .ZN(N27848));
    NANDX1 U14977 (.A1(n22007), .A2(n17178), .ZN(N27849));
    NOR2X1 U14978 (.A1(n24991), .A2(N2624), .ZN(N27850));
    NANDX1 U14979 (.A1(N7097), .A2(N7495), .ZN(n27851));
    INVX1 U14980 (.I(n17942), .ZN(n27852));
    NOR2X1 U14981 (.A1(N11059), .A2(N7879), .ZN(n27853));
    INVX1 U14982 (.I(n23706), .ZN(N27854));
    INVX1 U14983 (.I(N9643), .ZN(n27855));
    INVX1 U14984 (.I(n21949), .ZN(N27856));
    NOR2X1 U14985 (.A1(N6492), .A2(n14861), .ZN(n27857));
    NANDX1 U14986 (.A1(N12681), .A2(n17718), .ZN(n27858));
    NANDX1 U14987 (.A1(N12505), .A2(N1438), .ZN(n27859));
    NANDX1 U14988 (.A1(N9773), .A2(N7760), .ZN(n27860));
    NANDX1 U14989 (.A1(N1449), .A2(n14956), .ZN(N27861));
    NANDX1 U14990 (.A1(N4072), .A2(n14622), .ZN(n27862));
    NANDX1 U14991 (.A1(N335), .A2(n16196), .ZN(n27863));
    INVX1 U14992 (.I(n24608), .ZN(n27864));
    INVX1 U14993 (.I(N2626), .ZN(n27865));
    NOR2X1 U14994 (.A1(n25457), .A2(N5330), .ZN(n27866));
    NOR2X1 U14995 (.A1(N11289), .A2(N1776), .ZN(n27867));
    NANDX1 U14996 (.A1(n17780), .A2(n16636), .ZN(N27868));
    NOR2X1 U14997 (.A1(N4958), .A2(n23122), .ZN(n27869));
    NOR2X1 U14998 (.A1(n17462), .A2(n24559), .ZN(n27870));
    INVX1 U14999 (.I(n16002), .ZN(n27871));
    INVX1 U15000 (.I(n21550), .ZN(n27872));
    INVX1 U15001 (.I(N10539), .ZN(N27873));
    NOR2X1 U15002 (.A1(N10290), .A2(n25160), .ZN(n27874));
    NANDX1 U15003 (.A1(N10624), .A2(N4621), .ZN(n27875));
    NOR2X1 U15004 (.A1(n23999), .A2(N6372), .ZN(n27876));
    NOR2X1 U15005 (.A1(n24667), .A2(n20597), .ZN(n27877));
    NOR2X1 U15006 (.A1(N9476), .A2(N6383), .ZN(n27878));
    INVX1 U15007 (.I(n13864), .ZN(N27879));
    NOR2X1 U15008 (.A1(n17717), .A2(n19489), .ZN(n27880));
    INVX1 U15009 (.I(N4104), .ZN(n27881));
    NANDX1 U15010 (.A1(n24116), .A2(n17430), .ZN(n27882));
    NANDX1 U15011 (.A1(N3383), .A2(n13013), .ZN(N27883));
    NANDX1 U15012 (.A1(N9601), .A2(n23551), .ZN(n27884));
    INVX1 U15013 (.I(n19890), .ZN(n27885));
    NANDX1 U15014 (.A1(n22137), .A2(n19281), .ZN(N27886));
    INVX1 U15015 (.I(N10450), .ZN(N27887));
    NANDX1 U15016 (.A1(n22969), .A2(n15658), .ZN(n27888));
    NOR2X1 U15017 (.A1(N6831), .A2(n14963), .ZN(n27889));
    NOR2X1 U15018 (.A1(N1981), .A2(n16043), .ZN(N27890));
    NANDX1 U15019 (.A1(n14910), .A2(n22527), .ZN(n27891));
    INVX1 U15020 (.I(n21564), .ZN(n27892));
    NANDX1 U15021 (.A1(n24201), .A2(N8945), .ZN(n27893));
    NANDX1 U15022 (.A1(n14460), .A2(N12327), .ZN(N27894));
    NOR2X1 U15023 (.A1(N767), .A2(n21927), .ZN(n27895));
    INVX1 U15024 (.I(N3834), .ZN(N27896));
    NOR2X1 U15025 (.A1(n16092), .A2(n14738), .ZN(n27897));
    NOR2X1 U15026 (.A1(N7186), .A2(n13955), .ZN(n27898));
    NANDX1 U15027 (.A1(n18922), .A2(n18380), .ZN(n27899));
    NANDX1 U15028 (.A1(N250), .A2(N7840), .ZN(N27900));
    INVX1 U15029 (.I(N2230), .ZN(n27901));
    NANDX1 U15030 (.A1(N7379), .A2(N5907), .ZN(n27902));
    NOR2X1 U15031 (.A1(n19181), .A2(N1968), .ZN(N27903));
    NANDX1 U15032 (.A1(N6647), .A2(N10912), .ZN(n27904));
    INVX1 U15033 (.I(n21107), .ZN(n27905));
    NOR2X1 U15034 (.A1(n24194), .A2(n21873), .ZN(N27906));
    INVX1 U15035 (.I(n17077), .ZN(N27907));
    NANDX1 U15036 (.A1(N2281), .A2(n21936), .ZN(n27908));
    NOR2X1 U15037 (.A1(N1140), .A2(N3619), .ZN(n27909));
    INVX1 U15038 (.I(n20814), .ZN(n27910));
    NOR2X1 U15039 (.A1(n13580), .A2(n20695), .ZN(n27911));
    NOR2X1 U15040 (.A1(n21419), .A2(n24528), .ZN(n27912));
    NANDX1 U15041 (.A1(n19799), .A2(n20675), .ZN(n27913));
    NOR2X1 U15042 (.A1(N3972), .A2(N3121), .ZN(n27914));
    INVX1 U15043 (.I(n14774), .ZN(N27915));
    NOR2X1 U15044 (.A1(n13147), .A2(n18630), .ZN(n27916));
    NANDX1 U15045 (.A1(n25153), .A2(n17321), .ZN(n27917));
    INVX1 U15046 (.I(n22352), .ZN(N27918));
    NANDX1 U15047 (.A1(n19253), .A2(n24632), .ZN(n27919));
    NANDX1 U15048 (.A1(N498), .A2(n14539), .ZN(n27920));
    NOR2X1 U15049 (.A1(n21199), .A2(n24121), .ZN(n27921));
    NANDX1 U15050 (.A1(N9276), .A2(N8081), .ZN(N27922));
    INVX1 U15051 (.I(N5193), .ZN(n27923));
    INVX1 U15052 (.I(n14941), .ZN(n27924));
    NOR2X1 U15053 (.A1(N2279), .A2(N939), .ZN(n27925));
    NANDX1 U15054 (.A1(N5399), .A2(n14406), .ZN(n27926));
    NOR2X1 U15055 (.A1(N3933), .A2(N2050), .ZN(n27927));
    NOR2X1 U15056 (.A1(n23574), .A2(n15971), .ZN(n27928));
    NOR2X1 U15057 (.A1(N2850), .A2(N12820), .ZN(n27929));
    NANDX1 U15058 (.A1(N10870), .A2(N11949), .ZN(n27930));
    NOR2X1 U15059 (.A1(N11367), .A2(N985), .ZN(N27931));
    NOR2X1 U15060 (.A1(N7064), .A2(n25105), .ZN(N27932));
    INVX1 U15061 (.I(N5107), .ZN(n27933));
    INVX1 U15062 (.I(n23173), .ZN(n27934));
    NANDX1 U15063 (.A1(N3558), .A2(N1379), .ZN(N27935));
    NANDX1 U15064 (.A1(n20106), .A2(n16587), .ZN(n27936));
    INVX1 U15065 (.I(n14272), .ZN(n27937));
    INVX1 U15066 (.I(n15092), .ZN(n27938));
    NOR2X1 U15067 (.A1(n21810), .A2(N3988), .ZN(n27939));
    NANDX1 U15068 (.A1(N12278), .A2(n24474), .ZN(n27940));
    NOR2X1 U15069 (.A1(n25097), .A2(N5889), .ZN(N27941));
    NANDX1 U15070 (.A1(N311), .A2(n18134), .ZN(N27942));
    INVX1 U15071 (.I(N1295), .ZN(n27943));
    NANDX1 U15072 (.A1(N458), .A2(n15168), .ZN(N27944));
    INVX1 U15073 (.I(N5564), .ZN(n27945));
    NANDX1 U15074 (.A1(n17123), .A2(N4631), .ZN(n27946));
    INVX1 U15075 (.I(N7269), .ZN(N27947));
    NOR2X1 U15076 (.A1(n24049), .A2(n23856), .ZN(n27948));
    NOR2X1 U15077 (.A1(N12818), .A2(n18113), .ZN(N27949));
    INVX1 U15078 (.I(n19789), .ZN(n27950));
    NANDX1 U15079 (.A1(N7890), .A2(N10562), .ZN(n27951));
    NOR2X1 U15080 (.A1(N6862), .A2(n18454), .ZN(n27952));
    NOR2X1 U15081 (.A1(N12750), .A2(N11713), .ZN(n27953));
    NANDX1 U15082 (.A1(n19651), .A2(N5107), .ZN(N27954));
    NOR2X1 U15083 (.A1(N2815), .A2(N5564), .ZN(N27955));
    INVX1 U15084 (.I(n22267), .ZN(n27956));
    NOR2X1 U15085 (.A1(n20985), .A2(N2655), .ZN(n27957));
    INVX1 U15086 (.I(n24928), .ZN(N27958));
    NOR2X1 U15087 (.A1(n25019), .A2(N12242), .ZN(N27959));
    INVX1 U15088 (.I(n13830), .ZN(n27960));
    INVX1 U15089 (.I(n15157), .ZN(n27961));
    NANDX1 U15090 (.A1(N8113), .A2(n18344), .ZN(n27962));
    NOR2X1 U15091 (.A1(N7442), .A2(n19539), .ZN(n27963));
    NANDX1 U15092 (.A1(N393), .A2(N9095), .ZN(n27964));
    NOR2X1 U15093 (.A1(N874), .A2(n24464), .ZN(N27965));
    NANDX1 U15094 (.A1(N5980), .A2(N4393), .ZN(n27966));
    NOR2X1 U15095 (.A1(N312), .A2(n13759), .ZN(N27967));
    INVX1 U15096 (.I(n14477), .ZN(n27968));
    NOR2X1 U15097 (.A1(n22187), .A2(N7770), .ZN(n27969));
    NOR2X1 U15098 (.A1(n20878), .A2(n21556), .ZN(n27970));
    NOR2X1 U15099 (.A1(n17921), .A2(N9883), .ZN(n27971));
    INVX1 U15100 (.I(n21845), .ZN(n27972));
    NOR2X1 U15101 (.A1(N6111), .A2(n14687), .ZN(n27973));
    NOR2X1 U15102 (.A1(n13553), .A2(n22993), .ZN(N27974));
    NANDX1 U15103 (.A1(N2713), .A2(n20855), .ZN(n27975));
    NANDX1 U15104 (.A1(n17856), .A2(N8584), .ZN(N27976));
    INVX1 U15105 (.I(n23836), .ZN(N27977));
    NANDX1 U15106 (.A1(n15506), .A2(n12915), .ZN(n27978));
    NOR2X1 U15107 (.A1(N9537), .A2(N1889), .ZN(n27979));
    NOR2X1 U15108 (.A1(N6221), .A2(n23928), .ZN(n27980));
    NANDX1 U15109 (.A1(N1596), .A2(n19981), .ZN(n27981));
    NANDX1 U15110 (.A1(N8285), .A2(n18631), .ZN(n27982));
    NANDX1 U15111 (.A1(n18897), .A2(N9512), .ZN(n27983));
    NANDX1 U15112 (.A1(N8081), .A2(n14782), .ZN(N27984));
    NOR2X1 U15113 (.A1(n19841), .A2(N4568), .ZN(n27985));
    NANDX1 U15114 (.A1(n15194), .A2(n17123), .ZN(N27986));
    INVX1 U15115 (.I(n23777), .ZN(n27987));
    NOR2X1 U15116 (.A1(N1019), .A2(N19), .ZN(N27988));
    INVX1 U15117 (.I(n13933), .ZN(n27989));
    INVX1 U15118 (.I(N12437), .ZN(N27990));
    NANDX1 U15119 (.A1(n17798), .A2(N7426), .ZN(n27991));
    NOR2X1 U15120 (.A1(N3238), .A2(n23291), .ZN(n27992));
    NOR2X1 U15121 (.A1(N12623), .A2(n20343), .ZN(n27993));
    NOR2X1 U15122 (.A1(N8773), .A2(n13738), .ZN(N27994));
    NOR2X1 U15123 (.A1(n25304), .A2(N10586), .ZN(n27995));
    INVX1 U15124 (.I(N4383), .ZN(n27996));
    NOR2X1 U15125 (.A1(n22518), .A2(N445), .ZN(n27997));
    NOR2X1 U15126 (.A1(N2906), .A2(n14362), .ZN(n27998));
    NANDX1 U15127 (.A1(N1533), .A2(N4148), .ZN(n27999));
    NOR2X1 U15128 (.A1(n18703), .A2(n18080), .ZN(N28000));
    NANDX1 U15129 (.A1(N5638), .A2(N11436), .ZN(N28001));
    NOR2X1 U15130 (.A1(N1831), .A2(n14449), .ZN(n28002));
    NOR2X1 U15131 (.A1(n13889), .A2(N708), .ZN(N28003));
    NANDX1 U15132 (.A1(N8730), .A2(n19867), .ZN(n28004));
    NOR2X1 U15133 (.A1(N11235), .A2(n23036), .ZN(N28005));
    NOR2X1 U15134 (.A1(n21820), .A2(n15483), .ZN(n28006));
    NOR2X1 U15135 (.A1(n15512), .A2(N1266), .ZN(N28007));
    NOR2X1 U15136 (.A1(n24397), .A2(n18441), .ZN(n28008));
    INVX1 U15137 (.I(n20325), .ZN(n28009));
    NOR2X1 U15138 (.A1(N9639), .A2(N5038), .ZN(n28010));
    INVX1 U15139 (.I(n16486), .ZN(n28011));
    NANDX1 U15140 (.A1(n21849), .A2(N2419), .ZN(N28012));
    NANDX1 U15141 (.A1(n23679), .A2(N5635), .ZN(n28013));
    NANDX1 U15142 (.A1(N833), .A2(n20612), .ZN(n28014));
    INVX1 U15143 (.I(N9562), .ZN(n28015));
    INVX1 U15144 (.I(n16994), .ZN(n28016));
    NOR2X1 U15145 (.A1(N1277), .A2(n14530), .ZN(n28017));
    INVX1 U15146 (.I(N5528), .ZN(n28018));
    NOR2X1 U15147 (.A1(n21393), .A2(n21063), .ZN(n28019));
    NOR2X1 U15148 (.A1(n20288), .A2(n14002), .ZN(n28020));
    INVX1 U15149 (.I(N3878), .ZN(n28021));
    INVX1 U15150 (.I(N243), .ZN(n28022));
    NOR2X1 U15151 (.A1(n24683), .A2(n16728), .ZN(n28023));
    NOR2X1 U15152 (.A1(n21029), .A2(N7914), .ZN(n28024));
    INVX1 U15153 (.I(N7973), .ZN(n28025));
    NANDX1 U15154 (.A1(N392), .A2(N8806), .ZN(N28026));
    NANDX1 U15155 (.A1(n22690), .A2(n18367), .ZN(n28027));
    NANDX1 U15156 (.A1(N2949), .A2(N2429), .ZN(n28028));
    INVX1 U15157 (.I(n17478), .ZN(n28029));
    INVX1 U15158 (.I(n22242), .ZN(N28030));
    NOR2X1 U15159 (.A1(n18470), .A2(n17802), .ZN(n28031));
    NANDX1 U15160 (.A1(N2023), .A2(n20571), .ZN(N28032));
    NANDX1 U15161 (.A1(n20170), .A2(n17811), .ZN(N28033));
    INVX1 U15162 (.I(N3583), .ZN(n28034));
    NOR2X1 U15163 (.A1(n23573), .A2(N6536), .ZN(N28035));
    INVX1 U15164 (.I(n20254), .ZN(n28036));
    NANDX1 U15165 (.A1(n20490), .A2(n22569), .ZN(n28037));
    NOR2X1 U15166 (.A1(n18063), .A2(n19993), .ZN(N28038));
    NOR2X1 U15167 (.A1(N10928), .A2(N9929), .ZN(N28039));
    INVX1 U15168 (.I(N2124), .ZN(N28040));
    NANDX1 U15169 (.A1(N5866), .A2(n13471), .ZN(n28041));
    NANDX1 U15170 (.A1(N3056), .A2(n20708), .ZN(n28042));
    NOR2X1 U15171 (.A1(N7824), .A2(n22731), .ZN(n28043));
    NANDX1 U15172 (.A1(n14427), .A2(N6166), .ZN(n28044));
    INVX1 U15173 (.I(n21273), .ZN(n28045));
    NOR2X1 U15174 (.A1(N11854), .A2(N8111), .ZN(n28046));
    INVX1 U15175 (.I(n24371), .ZN(n28047));
    NANDX1 U15176 (.A1(n15376), .A2(N8127), .ZN(N28048));
    NANDX1 U15177 (.A1(N3628), .A2(N687), .ZN(n28049));
    NANDX1 U15178 (.A1(N299), .A2(N382), .ZN(n28050));
    NOR2X1 U15179 (.A1(N2956), .A2(n16775), .ZN(N28051));
    NANDX1 U15180 (.A1(N8821), .A2(n19013), .ZN(n28052));
    INVX1 U15181 (.I(N645), .ZN(n28053));
    NANDX1 U15182 (.A1(N2659), .A2(n22738), .ZN(N28054));
    NANDX1 U15183 (.A1(n16446), .A2(N11662), .ZN(n28055));
    NOR2X1 U15184 (.A1(N11309), .A2(N7432), .ZN(n28056));
    INVX1 U15185 (.I(n23163), .ZN(n28057));
    INVX1 U15186 (.I(N9946), .ZN(n28058));
    INVX1 U15187 (.I(n18405), .ZN(N28059));
    INVX1 U15188 (.I(N7693), .ZN(n28060));
    INVX1 U15189 (.I(n17716), .ZN(n28061));
    NANDX1 U15190 (.A1(n15790), .A2(N6782), .ZN(N28062));
    NANDX1 U15191 (.A1(n23175), .A2(N9738), .ZN(n28063));
    NOR2X1 U15192 (.A1(n20468), .A2(N7326), .ZN(n28064));
    NOR2X1 U15193 (.A1(N4408), .A2(N7970), .ZN(N28065));
    INVX1 U15194 (.I(N7067), .ZN(n28066));
    NANDX1 U15195 (.A1(n25284), .A2(N12280), .ZN(N28067));
    NOR2X1 U15196 (.A1(N6162), .A2(N12357), .ZN(N28068));
    INVX1 U15197 (.I(N11057), .ZN(n28069));
    INVX1 U15198 (.I(n17376), .ZN(n28070));
    NOR2X1 U15199 (.A1(N9583), .A2(n24548), .ZN(N28071));
    INVX1 U15200 (.I(N6044), .ZN(n28072));
    NOR2X1 U15201 (.A1(N4840), .A2(N3191), .ZN(N28073));
    NANDX1 U15202 (.A1(N11622), .A2(N3757), .ZN(N28074));
    INVX1 U15203 (.I(n21359), .ZN(N28075));
    NOR2X1 U15204 (.A1(N6380), .A2(N3182), .ZN(n28076));
    NOR2X1 U15205 (.A1(N10788), .A2(n25422), .ZN(n28077));
    NOR2X1 U15206 (.A1(N6622), .A2(n19394), .ZN(n28078));
    NOR2X1 U15207 (.A1(n18901), .A2(n25028), .ZN(n28079));
    NANDX1 U15208 (.A1(n20025), .A2(N1360), .ZN(N28080));
    INVX1 U15209 (.I(n18809), .ZN(n28081));
    NOR2X1 U15210 (.A1(n24589), .A2(N2890), .ZN(n28082));
    NANDX1 U15211 (.A1(N11713), .A2(n23203), .ZN(n28083));
    INVX1 U15212 (.I(n16553), .ZN(N28084));
    NOR2X1 U15213 (.A1(n15204), .A2(N2672), .ZN(N28085));
    NOR2X1 U15214 (.A1(N1116), .A2(N12798), .ZN(n28086));
    INVX1 U15215 (.I(N7496), .ZN(n28087));
    NANDX1 U15216 (.A1(n20960), .A2(n18283), .ZN(n28088));
    NANDX1 U15217 (.A1(n15742), .A2(n13672), .ZN(n28089));
    NOR2X1 U15218 (.A1(n24576), .A2(N7070), .ZN(n28090));
    NANDX1 U15219 (.A1(n14069), .A2(n15863), .ZN(n28091));
    NOR2X1 U15220 (.A1(N3386), .A2(N9169), .ZN(n28092));
    NOR2X1 U15221 (.A1(n16743), .A2(N12058), .ZN(n28093));
    NANDX1 U15222 (.A1(N2953), .A2(N9758), .ZN(n28094));
    NANDX1 U15223 (.A1(n19505), .A2(n24918), .ZN(n28095));
    INVX1 U15224 (.I(N10944), .ZN(n28096));
    NANDX1 U15225 (.A1(N3654), .A2(n23741), .ZN(n28097));
    NANDX1 U15226 (.A1(N11149), .A2(N2986), .ZN(n28098));
    NANDX1 U15227 (.A1(n18199), .A2(n21921), .ZN(N28099));
    NANDX1 U15228 (.A1(N6368), .A2(N9246), .ZN(N28100));
    NANDX1 U15229 (.A1(N2205), .A2(N10367), .ZN(n28101));
    NOR2X1 U15230 (.A1(n18067), .A2(N1614), .ZN(n28102));
    NANDX1 U15231 (.A1(N1734), .A2(n14634), .ZN(n28103));
    NOR2X1 U15232 (.A1(N2559), .A2(n22970), .ZN(n28104));
    INVX1 U15233 (.I(N1085), .ZN(n28105));
    NOR2X1 U15234 (.A1(N3838), .A2(n14770), .ZN(n28106));
    INVX1 U15235 (.I(n14781), .ZN(n28107));
    NOR2X1 U15236 (.A1(n16495), .A2(N1788), .ZN(N28108));
    NANDX1 U15237 (.A1(n16411), .A2(N4773), .ZN(n28109));
    INVX1 U15238 (.I(n23377), .ZN(n28110));
    NOR2X1 U15239 (.A1(n19894), .A2(n18512), .ZN(n28111));
    NANDX1 U15240 (.A1(N3812), .A2(N9484), .ZN(n28112));
    NOR2X1 U15241 (.A1(N1798), .A2(n16319), .ZN(n28113));
    NOR2X1 U15242 (.A1(n17440), .A2(n18052), .ZN(n28114));
    INVX1 U15243 (.I(n24322), .ZN(n28115));
    NANDX1 U15244 (.A1(N821), .A2(n22925), .ZN(n28116));
    NANDX1 U15245 (.A1(N11125), .A2(n15530), .ZN(N28117));
    NANDX1 U15246 (.A1(N12734), .A2(n19078), .ZN(n28118));
    INVX1 U15247 (.I(n17996), .ZN(N28119));
    NOR2X1 U15248 (.A1(n14077), .A2(n23174), .ZN(N28120));
    NOR2X1 U15249 (.A1(n23623), .A2(n21048), .ZN(n28121));
    NOR2X1 U15250 (.A1(N6782), .A2(N2825), .ZN(n28122));
    NANDX1 U15251 (.A1(N10593), .A2(N12308), .ZN(N28123));
    NANDX1 U15252 (.A1(N12391), .A2(N3124), .ZN(n28124));
    INVX1 U15253 (.I(n18598), .ZN(n28125));
    NANDX1 U15254 (.A1(N2172), .A2(N6186), .ZN(n28126));
    NANDX1 U15255 (.A1(n17263), .A2(N3608), .ZN(n28127));
    INVX1 U15256 (.I(n17155), .ZN(N28128));
    INVX1 U15257 (.I(n21317), .ZN(N28129));
    NANDX1 U15258 (.A1(N12712), .A2(n17414), .ZN(N28130));
    INVX1 U15259 (.I(N8075), .ZN(N28131));
    INVX1 U15260 (.I(n20052), .ZN(n28132));
    NOR2X1 U15261 (.A1(N7146), .A2(N4365), .ZN(n28133));
    NOR2X1 U15262 (.A1(n13928), .A2(N7189), .ZN(N28134));
    INVX1 U15263 (.I(n24520), .ZN(n28135));
    NANDX1 U15264 (.A1(N736), .A2(N176), .ZN(n28136));
    INVX1 U15265 (.I(n13825), .ZN(n28137));
    INVX1 U15266 (.I(N10098), .ZN(n28138));
    NOR2X1 U15267 (.A1(n24959), .A2(n18186), .ZN(n28139));
    NANDX1 U15268 (.A1(n17334), .A2(N2), .ZN(N28140));
    NOR2X1 U15269 (.A1(N10968), .A2(n21318), .ZN(n28141));
    INVX1 U15270 (.I(N12447), .ZN(n28142));
    NOR2X1 U15271 (.A1(n17979), .A2(N9289), .ZN(n28143));
    NOR2X1 U15272 (.A1(N1296), .A2(N6266), .ZN(n28144));
    NANDX1 U15273 (.A1(N5660), .A2(n18837), .ZN(N28145));
    NANDX1 U15274 (.A1(N1616), .A2(n20706), .ZN(n28146));
    NOR2X1 U15275 (.A1(n24150), .A2(n21441), .ZN(n28147));
    INVX1 U15276 (.I(N10035), .ZN(n28148));
    INVX1 U15277 (.I(n24559), .ZN(N28149));
    INVX1 U15278 (.I(n14527), .ZN(n28150));
    INVX1 U15279 (.I(N1584), .ZN(n28151));
    NOR2X1 U15280 (.A1(N4614), .A2(n15855), .ZN(N28152));
    NOR2X1 U15281 (.A1(n15581), .A2(N11670), .ZN(N28153));
    INVX1 U15282 (.I(n16795), .ZN(n28154));
    NOR2X1 U15283 (.A1(n15841), .A2(N582), .ZN(N28155));
    NOR2X1 U15284 (.A1(n17136), .A2(N6847), .ZN(n28156));
    INVX1 U15285 (.I(N11564), .ZN(N28157));
    NANDX1 U15286 (.A1(N9675), .A2(N1947), .ZN(n28158));
    NANDX1 U15287 (.A1(n15285), .A2(N594), .ZN(n28159));
    NANDX1 U15288 (.A1(n21070), .A2(n24898), .ZN(n28160));
    NOR2X1 U15289 (.A1(N8894), .A2(n22566), .ZN(n28161));
    NOR2X1 U15290 (.A1(n21676), .A2(n24149), .ZN(n28162));
    INVX1 U15291 (.I(N787), .ZN(n28163));
    INVX1 U15292 (.I(n20730), .ZN(n28164));
    NANDX1 U15293 (.A1(n14938), .A2(n18591), .ZN(n28165));
    NOR2X1 U15294 (.A1(n17372), .A2(N8929), .ZN(N28166));
    INVX1 U15295 (.I(n16558), .ZN(N28167));
    INVX1 U15296 (.I(n18124), .ZN(N28168));
    NANDX1 U15297 (.A1(n15164), .A2(n18305), .ZN(n28169));
    NANDX1 U15298 (.A1(N5878), .A2(N2456), .ZN(n28170));
    NANDX1 U15299 (.A1(n20742), .A2(N8048), .ZN(n28171));
    NANDX1 U15300 (.A1(N8905), .A2(n23403), .ZN(n28172));
    NANDX1 U15301 (.A1(N5968), .A2(n16549), .ZN(N28173));
    NOR2X1 U15302 (.A1(N4614), .A2(N9513), .ZN(n28174));
    NOR2X1 U15303 (.A1(N7882), .A2(n19010), .ZN(N28175));
    NANDX1 U15304 (.A1(n22820), .A2(N12099), .ZN(n28176));
    INVX1 U15305 (.I(n14689), .ZN(n28177));
    INVX1 U15306 (.I(n16966), .ZN(n28178));
    NOR2X1 U15307 (.A1(n13395), .A2(N9587), .ZN(n28179));
    NOR2X1 U15308 (.A1(n17326), .A2(n16659), .ZN(N28180));
    INVX1 U15309 (.I(n23204), .ZN(N28181));
    NANDX1 U15310 (.A1(N6402), .A2(N7211), .ZN(n28182));
    INVX1 U15311 (.I(N12871), .ZN(n28183));
    INVX1 U15312 (.I(n13830), .ZN(N28184));
    NOR2X1 U15313 (.A1(n22083), .A2(n19147), .ZN(n28185));
    NOR2X1 U15314 (.A1(N1194), .A2(n17427), .ZN(n28186));
    NANDX1 U15315 (.A1(n23346), .A2(N10935), .ZN(N28187));
    NOR2X1 U15316 (.A1(N9431), .A2(N11801), .ZN(N28188));
    INVX1 U15317 (.I(n24119), .ZN(N28189));
    NOR2X1 U15318 (.A1(N5378), .A2(n18631), .ZN(n28190));
    NANDX1 U15319 (.A1(n14965), .A2(n21550), .ZN(n28191));
    INVX1 U15320 (.I(n20391), .ZN(n28192));
    NANDX1 U15321 (.A1(n16320), .A2(N2771), .ZN(n28193));
    NANDX1 U15322 (.A1(n23530), .A2(n18701), .ZN(n28194));
    NOR2X1 U15323 (.A1(n14143), .A2(n21298), .ZN(n28195));
    NANDX1 U15324 (.A1(n24993), .A2(n14942), .ZN(N28196));
    NANDX1 U15325 (.A1(n14954), .A2(n21137), .ZN(n28197));
    INVX1 U15326 (.I(N12797), .ZN(n28198));
    NANDX1 U15327 (.A1(n18618), .A2(n22227), .ZN(n28199));
    INVX1 U15328 (.I(n18262), .ZN(N28200));
    NANDX1 U15329 (.A1(n17499), .A2(n23640), .ZN(n28201));
    INVX1 U15330 (.I(N4522), .ZN(n28202));
    INVX1 U15331 (.I(N1825), .ZN(n28203));
    NOR2X1 U15332 (.A1(n22260), .A2(N7641), .ZN(n28204));
    NOR2X1 U15333 (.A1(n25031), .A2(n22896), .ZN(n28205));
    NANDX1 U15334 (.A1(N6997), .A2(N17), .ZN(n28206));
    NANDX1 U15335 (.A1(N2792), .A2(N8408), .ZN(N28207));
    NOR2X1 U15336 (.A1(N6502), .A2(n22870), .ZN(n28208));
    NOR2X1 U15337 (.A1(N2136), .A2(n22028), .ZN(N28209));
    NOR2X1 U15338 (.A1(n22974), .A2(n15143), .ZN(N28210));
    NANDX1 U15339 (.A1(N4608), .A2(n22172), .ZN(n28211));
    INVX1 U15340 (.I(N10874), .ZN(N28212));
    INVX1 U15341 (.I(n17514), .ZN(N28213));
    INVX1 U15342 (.I(n25216), .ZN(n28214));
    NANDX1 U15343 (.A1(N1802), .A2(n21974), .ZN(n28215));
    NANDX1 U15344 (.A1(n15759), .A2(N10270), .ZN(N28216));
    NOR2X1 U15345 (.A1(n16512), .A2(N6034), .ZN(n28217));
    NOR2X1 U15346 (.A1(N5905), .A2(N8825), .ZN(n28218));
    NANDX1 U15347 (.A1(N9058), .A2(n15326), .ZN(n28219));
    NOR2X1 U15348 (.A1(N1663), .A2(N6229), .ZN(n28220));
    INVX1 U15349 (.I(N7064), .ZN(N28221));
    INVX1 U15350 (.I(n22402), .ZN(n28222));
    NANDX1 U15351 (.A1(n22577), .A2(n19072), .ZN(N28223));
    NOR2X1 U15352 (.A1(n22219), .A2(n16916), .ZN(N28224));
    NOR2X1 U15353 (.A1(N880), .A2(n16630), .ZN(N28225));
    NOR2X1 U15354 (.A1(N2681), .A2(N1869), .ZN(n28226));
    INVX1 U15355 (.I(N7207), .ZN(n28227));
    NANDX1 U15356 (.A1(N1961), .A2(n23719), .ZN(N28228));
    INVX1 U15357 (.I(N3883), .ZN(n28229));
    NOR2X1 U15358 (.A1(n15763), .A2(n25445), .ZN(N28230));
    INVX1 U15359 (.I(n19857), .ZN(N28231));
    NOR2X1 U15360 (.A1(n17879), .A2(N583), .ZN(n28232));
    INVX1 U15361 (.I(n13710), .ZN(n28233));
    NANDX1 U15362 (.A1(N11798), .A2(N11666), .ZN(n28234));
    NOR2X1 U15363 (.A1(n19637), .A2(N10127), .ZN(n28235));
    INVX1 U15364 (.I(n25321), .ZN(N28236));
    NANDX1 U15365 (.A1(N1990), .A2(n16448), .ZN(n28237));
    INVX1 U15366 (.I(n18940), .ZN(n28238));
    NOR2X1 U15367 (.A1(N2269), .A2(n14915), .ZN(N28239));
    INVX1 U15368 (.I(n18499), .ZN(N28240));
    INVX1 U15369 (.I(N657), .ZN(n28241));
    NOR2X1 U15370 (.A1(n20289), .A2(N5187), .ZN(n28242));
    NOR2X1 U15371 (.A1(n25273), .A2(n25043), .ZN(N28243));
    NANDX1 U15372 (.A1(N6417), .A2(N124), .ZN(n28244));
    NOR2X1 U15373 (.A1(n20126), .A2(n18676), .ZN(n28245));
    NOR2X1 U15374 (.A1(N6290), .A2(n23070), .ZN(n28246));
    NANDX1 U15375 (.A1(N5184), .A2(n24181), .ZN(N28247));
    INVX1 U15376 (.I(N8821), .ZN(n28248));
    NOR2X1 U15377 (.A1(N10897), .A2(n22268), .ZN(N28249));
    NANDX1 U15378 (.A1(N3710), .A2(n13305), .ZN(n28250));
    NANDX1 U15379 (.A1(N11698), .A2(N6301), .ZN(N28251));
    NANDX1 U15380 (.A1(N1122), .A2(n17450), .ZN(n28252));
    NANDX1 U15381 (.A1(N6309), .A2(n17309), .ZN(n28253));
    INVX1 U15382 (.I(N5849), .ZN(n28254));
    INVX1 U15383 (.I(N3697), .ZN(N28255));
    NANDX1 U15384 (.A1(n24738), .A2(n23823), .ZN(n28256));
    NANDX1 U15385 (.A1(N10965), .A2(n18880), .ZN(n28257));
    INVX1 U15386 (.I(N5597), .ZN(n28258));
    INVX1 U15387 (.I(n23931), .ZN(N28259));
    NOR2X1 U15388 (.A1(n21652), .A2(n13366), .ZN(n28260));
    INVX1 U15389 (.I(N7185), .ZN(N28261));
    NOR2X1 U15390 (.A1(N3420), .A2(n20489), .ZN(N28262));
    NANDX1 U15391 (.A1(N3886), .A2(n15558), .ZN(N28263));
    INVX1 U15392 (.I(N5007), .ZN(n28264));
    NANDX1 U15393 (.A1(n19761), .A2(N11315), .ZN(n28265));
    NOR2X1 U15394 (.A1(N5809), .A2(n17164), .ZN(N28266));
    NOR2X1 U15395 (.A1(N9505), .A2(N11903), .ZN(n28267));
    NOR2X1 U15396 (.A1(n22095), .A2(n14086), .ZN(N28268));
    NOR2X1 U15397 (.A1(N4240), .A2(n13836), .ZN(n28269));
    NANDX1 U15398 (.A1(n17071), .A2(N1032), .ZN(n28270));
    INVX1 U15399 (.I(N1988), .ZN(n28271));
    NOR2X1 U15400 (.A1(N9011), .A2(N9172), .ZN(n28272));
    INVX1 U15401 (.I(N1199), .ZN(n28273));
    INVX1 U15402 (.I(n25007), .ZN(N28274));
    NOR2X1 U15403 (.A1(n22754), .A2(N10524), .ZN(N28275));
    NOR2X1 U15404 (.A1(n19026), .A2(n19052), .ZN(n28276));
    NOR2X1 U15405 (.A1(n21375), .A2(n24860), .ZN(n28277));
    NANDX1 U15406 (.A1(N11796), .A2(n23132), .ZN(N28278));
    NANDX1 U15407 (.A1(n15723), .A2(n19725), .ZN(n28279));
    NANDX1 U15408 (.A1(N5112), .A2(n23964), .ZN(N28280));
    NANDX1 U15409 (.A1(n14367), .A2(N4300), .ZN(N28281));
    NOR2X1 U15410 (.A1(N12435), .A2(N6287), .ZN(n28282));
    INVX1 U15411 (.I(N10214), .ZN(N28283));
    NOR2X1 U15412 (.A1(N3365), .A2(N11412), .ZN(n28284));
    NOR2X1 U15413 (.A1(n17139), .A2(N5263), .ZN(N28285));
    NANDX1 U15414 (.A1(N2160), .A2(n15352), .ZN(N28286));
    NANDX1 U15415 (.A1(N9979), .A2(N22), .ZN(n28287));
    NOR2X1 U15416 (.A1(n23606), .A2(n16125), .ZN(N28288));
    NANDX1 U15417 (.A1(n21236), .A2(N7397), .ZN(n28289));
    NOR2X1 U15418 (.A1(n15458), .A2(N12753), .ZN(n28290));
    NOR2X1 U15419 (.A1(N2687), .A2(n20713), .ZN(N28291));
    NOR2X1 U15420 (.A1(N6987), .A2(n18471), .ZN(N28292));
    NOR2X1 U15421 (.A1(n13273), .A2(n19394), .ZN(N28293));
    INVX1 U15422 (.I(N6267), .ZN(n28294));
    NOR2X1 U15423 (.A1(N11731), .A2(n17689), .ZN(n28295));
    NOR2X1 U15424 (.A1(n16993), .A2(N860), .ZN(N28296));
    NANDX1 U15425 (.A1(n21112), .A2(n17327), .ZN(n28297));
    NANDX1 U15426 (.A1(N9902), .A2(N7202), .ZN(n28298));
    NOR2X1 U15427 (.A1(n14794), .A2(N8872), .ZN(n28299));
    NOR2X1 U15428 (.A1(n22190), .A2(N763), .ZN(N28300));
    INVX1 U15429 (.I(N9441), .ZN(n28301));
    NOR2X1 U15430 (.A1(n16049), .A2(N4651), .ZN(n28302));
    INVX1 U15431 (.I(N11803), .ZN(n28303));
    NANDX1 U15432 (.A1(N2276), .A2(n25075), .ZN(n28304));
    NOR2X1 U15433 (.A1(N2595), .A2(n20110), .ZN(n28305));
    NOR2X1 U15434 (.A1(N3093), .A2(N12296), .ZN(N28306));
    NOR2X1 U15435 (.A1(N8853), .A2(n13156), .ZN(n28307));
    NANDX1 U15436 (.A1(n18732), .A2(n19250), .ZN(n28308));
    INVX1 U15437 (.I(n17401), .ZN(n28309));
    INVX1 U15438 (.I(n20797), .ZN(n28310));
    NOR2X1 U15439 (.A1(N9820), .A2(n18702), .ZN(n28311));
    NOR2X1 U15440 (.A1(n24852), .A2(n20831), .ZN(n28312));
    NOR2X1 U15441 (.A1(N11384), .A2(N145), .ZN(n28313));
    NOR2X1 U15442 (.A1(N12321), .A2(N11947), .ZN(n28314));
    NOR2X1 U15443 (.A1(N3364), .A2(N288), .ZN(N28315));
    NOR2X1 U15444 (.A1(n20228), .A2(n20397), .ZN(N28316));
    NANDX1 U15445 (.A1(N12088), .A2(n21460), .ZN(n28317));
    NANDX1 U15446 (.A1(n20940), .A2(N9113), .ZN(n28318));
    INVX1 U15447 (.I(N2937), .ZN(N28319));
    NOR2X1 U15448 (.A1(n21394), .A2(n20338), .ZN(n28320));
    INVX1 U15449 (.I(n16688), .ZN(n28321));
    NANDX1 U15450 (.A1(N5434), .A2(n24157), .ZN(N28322));
    INVX1 U15451 (.I(N4783), .ZN(N28323));
    NANDX1 U15452 (.A1(N9533), .A2(n16166), .ZN(n28324));
    NOR2X1 U15453 (.A1(n18808), .A2(n17254), .ZN(n28325));
    NANDX1 U15454 (.A1(n14470), .A2(N9385), .ZN(n28326));
    NANDX1 U15455 (.A1(n15912), .A2(n18380), .ZN(N28327));
    INVX1 U15456 (.I(N9158), .ZN(n28328));
    NOR2X1 U15457 (.A1(N3289), .A2(n22871), .ZN(n28329));
    NANDX1 U15458 (.A1(N1170), .A2(n14407), .ZN(N28330));
    NOR2X1 U15459 (.A1(N7067), .A2(N10298), .ZN(N28331));
    INVX1 U15460 (.I(n13913), .ZN(N28332));
    INVX1 U15461 (.I(n17009), .ZN(N28333));
    INVX1 U15462 (.I(N3176), .ZN(n28334));
    NANDX1 U15463 (.A1(n24128), .A2(N11429), .ZN(n28335));
    NOR2X1 U15464 (.A1(N3560), .A2(N8594), .ZN(n28336));
    NANDX1 U15465 (.A1(N9581), .A2(N6474), .ZN(N28337));
    NANDX1 U15466 (.A1(N7734), .A2(n18911), .ZN(N28338));
    NOR2X1 U15467 (.A1(N611), .A2(n15010), .ZN(n28339));
    INVX1 U15468 (.I(n19846), .ZN(N28340));
    NANDX1 U15469 (.A1(n19769), .A2(n23285), .ZN(N28341));
    NANDX1 U15470 (.A1(N8673), .A2(N4159), .ZN(n28342));
    NANDX1 U15471 (.A1(N7738), .A2(n19640), .ZN(N28343));
    INVX1 U15472 (.I(N12258), .ZN(n28344));
    NOR2X1 U15473 (.A1(N11825), .A2(n15433), .ZN(n28345));
    NOR2X1 U15474 (.A1(n24721), .A2(N1359), .ZN(n28346));
    NOR2X1 U15475 (.A1(n17048), .A2(n24223), .ZN(n28347));
    INVX1 U15476 (.I(n15396), .ZN(n28348));
    INVX1 U15477 (.I(N11005), .ZN(n28349));
    NANDX1 U15478 (.A1(n12873), .A2(n24248), .ZN(n28350));
    NANDX1 U15479 (.A1(n16650), .A2(N6876), .ZN(N28351));
    NANDX1 U15480 (.A1(n23716), .A2(n15412), .ZN(n28352));
    INVX1 U15481 (.I(n20719), .ZN(n28353));
    NANDX1 U15482 (.A1(N11830), .A2(N10519), .ZN(n28354));
    NOR2X1 U15483 (.A1(n20237), .A2(n17268), .ZN(N28355));
    NOR2X1 U15484 (.A1(n20151), .A2(N3591), .ZN(n28356));
    INVX1 U15485 (.I(n19515), .ZN(N28357));
    NOR2X1 U15486 (.A1(N1671), .A2(N5397), .ZN(n28358));
    INVX1 U15487 (.I(n14661), .ZN(n28359));
    INVX1 U15488 (.I(N12787), .ZN(N28360));
    NANDX1 U15489 (.A1(n21880), .A2(N10414), .ZN(n28361));
    NOR2X1 U15490 (.A1(n20625), .A2(N11689), .ZN(N28362));
    INVX1 U15491 (.I(n16268), .ZN(n28363));
    NANDX1 U15492 (.A1(n25126), .A2(N6177), .ZN(n28364));
    NOR2X1 U15493 (.A1(n20342), .A2(n19028), .ZN(n28365));
    NANDX1 U15494 (.A1(n19628), .A2(N2882), .ZN(N28366));
    NOR2X1 U15495 (.A1(N11394), .A2(n24495), .ZN(N28367));
    INVX1 U15496 (.I(N3752), .ZN(n28368));
    INVX1 U15497 (.I(n13239), .ZN(N28369));
    NANDX1 U15498 (.A1(N976), .A2(N7403), .ZN(N28370));
    NANDX1 U15499 (.A1(n15636), .A2(n18278), .ZN(n28371));
    INVX1 U15500 (.I(n24258), .ZN(n28372));
    NOR2X1 U15501 (.A1(n18956), .A2(n23288), .ZN(N28373));
    NANDX1 U15502 (.A1(n19412), .A2(n24698), .ZN(n28374));
    NANDX1 U15503 (.A1(n15486), .A2(n13089), .ZN(n28375));
    NANDX1 U15504 (.A1(n19231), .A2(n22198), .ZN(N28376));
    NOR2X1 U15505 (.A1(n23572), .A2(N5092), .ZN(N28377));
    NOR2X1 U15506 (.A1(N11416), .A2(n16485), .ZN(N28378));
    INVX1 U15507 (.I(N5140), .ZN(n28379));
    NANDX1 U15508 (.A1(n21767), .A2(N7146), .ZN(n28380));
    INVX1 U15509 (.I(N11510), .ZN(n28381));
    NOR2X1 U15510 (.A1(n14357), .A2(N1644), .ZN(n28382));
    NANDX1 U15511 (.A1(n22899), .A2(n14669), .ZN(N28383));
    NANDX1 U15512 (.A1(N5121), .A2(N1223), .ZN(n28384));
    INVX1 U15513 (.I(n24532), .ZN(n28385));
    NOR2X1 U15514 (.A1(n15909), .A2(n14516), .ZN(n28386));
    NANDX1 U15515 (.A1(n14432), .A2(N8244), .ZN(n28387));
    NANDX1 U15516 (.A1(n20751), .A2(n20583), .ZN(N28388));
    NOR2X1 U15517 (.A1(n18718), .A2(N6497), .ZN(n28389));
    NOR2X1 U15518 (.A1(N4446), .A2(N11636), .ZN(n28390));
    NANDX1 U15519 (.A1(n14981), .A2(N7550), .ZN(N28391));
    NANDX1 U15520 (.A1(N988), .A2(N10866), .ZN(n28392));
    INVX1 U15521 (.I(n16901), .ZN(n28393));
    NOR2X1 U15522 (.A1(N3740), .A2(n20338), .ZN(N28394));
    INVX1 U15523 (.I(N8860), .ZN(N28395));
    INVX1 U15524 (.I(n18800), .ZN(n28396));
    NOR2X1 U15525 (.A1(N10745), .A2(n23476), .ZN(n28397));
    NOR2X1 U15526 (.A1(N1786), .A2(N1173), .ZN(N28398));
    NOR2X1 U15527 (.A1(n15024), .A2(N10691), .ZN(n28399));
    INVX1 U15528 (.I(n19084), .ZN(N28400));
    NOR2X1 U15529 (.A1(n24030), .A2(n17163), .ZN(n28401));
    INVX1 U15530 (.I(N10163), .ZN(N28402));
    NANDX1 U15531 (.A1(N868), .A2(N6480), .ZN(n28403));
    INVX1 U15532 (.I(n16126), .ZN(n28404));
    INVX1 U15533 (.I(n22575), .ZN(n28405));
    NANDX1 U15534 (.A1(n13070), .A2(N812), .ZN(n28406));
    NOR2X1 U15535 (.A1(n19540), .A2(n23941), .ZN(N28407));
    INVX1 U15536 (.I(N1605), .ZN(n28408));
    NANDX1 U15537 (.A1(N966), .A2(n13848), .ZN(n28409));
    NANDX1 U15538 (.A1(n17021), .A2(n15021), .ZN(n28410));
    NANDX1 U15539 (.A1(N6543), .A2(N209), .ZN(n28411));
    NANDX1 U15540 (.A1(n14394), .A2(n18385), .ZN(n28412));
    INVX1 U15541 (.I(n20324), .ZN(N28413));
    INVX1 U15542 (.I(N3938), .ZN(N28414));
    NOR2X1 U15543 (.A1(n19410), .A2(n24687), .ZN(N28415));
    NANDX1 U15544 (.A1(N10033), .A2(n16530), .ZN(N28416));
    INVX1 U15545 (.I(N6325), .ZN(n28417));
    NANDX1 U15546 (.A1(n24988), .A2(N11721), .ZN(n28418));
    INVX1 U15547 (.I(n23426), .ZN(n28419));
    NOR2X1 U15548 (.A1(n14009), .A2(N7288), .ZN(N28420));
    NANDX1 U15549 (.A1(n16624), .A2(n13554), .ZN(n28421));
    INVX1 U15550 (.I(N6142), .ZN(n28422));
    INVX1 U15551 (.I(n15239), .ZN(n28423));
    NANDX1 U15552 (.A1(N12018), .A2(N4130), .ZN(N28424));
    NOR2X1 U15553 (.A1(N5793), .A2(n24453), .ZN(N28425));
    INVX1 U15554 (.I(n24000), .ZN(n28426));
    NANDX1 U15555 (.A1(N451), .A2(n23184), .ZN(n28427));
    NOR2X1 U15556 (.A1(N10483), .A2(N2979), .ZN(N28428));
    INVX1 U15557 (.I(N5575), .ZN(n28429));
    NOR2X1 U15558 (.A1(N6547), .A2(n17296), .ZN(n28430));
    INVX1 U15559 (.I(n18740), .ZN(n28431));
    INVX1 U15560 (.I(N11023), .ZN(n28432));
    NANDX1 U15561 (.A1(n25183), .A2(N2144), .ZN(N28433));
    INVX1 U15562 (.I(N8377), .ZN(n28434));
    NANDX1 U15563 (.A1(N8385), .A2(n23615), .ZN(n28435));
    NOR2X1 U15564 (.A1(N9170), .A2(n16512), .ZN(n28436));
    NOR2X1 U15565 (.A1(n14962), .A2(N4231), .ZN(n28437));
    NANDX1 U15566 (.A1(N2227), .A2(n14054), .ZN(N28438));
    NANDX1 U15567 (.A1(n25411), .A2(n22441), .ZN(n28439));
    INVX1 U15568 (.I(n17157), .ZN(n28440));
    NANDX1 U15569 (.A1(n20530), .A2(n13000), .ZN(n28441));
    INVX1 U15570 (.I(N12323), .ZN(N28442));
    NANDX1 U15571 (.A1(n18053), .A2(n20328), .ZN(n28443));
    NANDX1 U15572 (.A1(n18577), .A2(n20008), .ZN(n28444));
    NANDX1 U15573 (.A1(n21423), .A2(n17153), .ZN(n28445));
    INVX1 U15574 (.I(N4305), .ZN(n28446));
    NANDX1 U15575 (.A1(N12403), .A2(n13475), .ZN(N28447));
    NANDX1 U15576 (.A1(N6845), .A2(n17204), .ZN(n28448));
    NANDX1 U15577 (.A1(N7829), .A2(n19431), .ZN(N28449));
    INVX1 U15578 (.I(n23533), .ZN(n28450));
    NOR2X1 U15579 (.A1(n13302), .A2(n12985), .ZN(n28451));
    NANDX1 U15580 (.A1(N6069), .A2(N8012), .ZN(n28452));
    NOR2X1 U15581 (.A1(n19652), .A2(N9102), .ZN(N28453));
    NANDX1 U15582 (.A1(N12202), .A2(n18197), .ZN(N28454));
    NOR2X1 U15583 (.A1(n19546), .A2(N1471), .ZN(n28455));
    NOR2X1 U15584 (.A1(N4235), .A2(n18623), .ZN(n28456));
    INVX1 U15585 (.I(N8539), .ZN(n28457));
    NOR2X1 U15586 (.A1(N3689), .A2(N10781), .ZN(n28458));
    INVX1 U15587 (.I(N10533), .ZN(n28459));
    NANDX1 U15588 (.A1(N8775), .A2(N7129), .ZN(n28460));
    INVX1 U15589 (.I(n25138), .ZN(n28461));
    NOR2X1 U15590 (.A1(n21825), .A2(N1705), .ZN(N28462));
    NOR2X1 U15591 (.A1(N10353), .A2(N7773), .ZN(n28463));
    INVX1 U15592 (.I(N11881), .ZN(N28464));
    INVX1 U15593 (.I(N12792), .ZN(n28465));
    NOR2X1 U15594 (.A1(N2891), .A2(n19757), .ZN(n28466));
    INVX1 U15595 (.I(n22437), .ZN(n28467));
    NANDX1 U15596 (.A1(N12781), .A2(n15439), .ZN(N28468));
    NOR2X1 U15597 (.A1(N4066), .A2(N12745), .ZN(n28469));
    NOR2X1 U15598 (.A1(N7754), .A2(n23526), .ZN(N28470));
    NANDX1 U15599 (.A1(N7054), .A2(N3544), .ZN(n28471));
    NANDX1 U15600 (.A1(N2950), .A2(N2992), .ZN(n28472));
    NOR2X1 U15601 (.A1(n22378), .A2(n13584), .ZN(N28473));
    NOR2X1 U15602 (.A1(n18057), .A2(n23936), .ZN(N28474));
    NOR2X1 U15603 (.A1(N10515), .A2(N10314), .ZN(n28475));
    INVX1 U15604 (.I(N12074), .ZN(n28476));
    INVX1 U15605 (.I(n24275), .ZN(n28477));
    INVX1 U15606 (.I(n16263), .ZN(n28478));
    NANDX1 U15607 (.A1(N2052), .A2(n17811), .ZN(n28479));
    NOR2X1 U15608 (.A1(N5166), .A2(N10644), .ZN(N28480));
    NOR2X1 U15609 (.A1(n19703), .A2(n18398), .ZN(n28481));
    INVX1 U15610 (.I(n15202), .ZN(N28482));
    NOR2X1 U15611 (.A1(N2991), .A2(N8243), .ZN(n28483));
    NANDX1 U15612 (.A1(n20252), .A2(n15190), .ZN(N28484));
    NOR2X1 U15613 (.A1(N8333), .A2(n23842), .ZN(n28485));
    INVX1 U15614 (.I(N6767), .ZN(n28486));
    NANDX1 U15615 (.A1(n20150), .A2(N5848), .ZN(n28487));
    NOR2X1 U15616 (.A1(n20992), .A2(n17118), .ZN(n28488));
    INVX1 U15617 (.I(N1817), .ZN(N28489));
    NOR2X1 U15618 (.A1(n19393), .A2(n18139), .ZN(n28490));
    INVX1 U15619 (.I(N8073), .ZN(n28491));
    INVX1 U15620 (.I(n13868), .ZN(N28492));
    NANDX1 U15621 (.A1(N6272), .A2(N6763), .ZN(n28493));
    NANDX1 U15622 (.A1(N10241), .A2(N9749), .ZN(n28494));
    NOR2X1 U15623 (.A1(N7252), .A2(N1415), .ZN(n28495));
    NOR2X1 U15624 (.A1(n22441), .A2(n18497), .ZN(n28496));
    NOR2X1 U15625 (.A1(n20780), .A2(N2630), .ZN(n28497));
    NANDX1 U15626 (.A1(n24311), .A2(N11548), .ZN(n28498));
    NOR2X1 U15627 (.A1(N9454), .A2(N7037), .ZN(n28499));
    INVX1 U15628 (.I(N7638), .ZN(n28500));
    INVX1 U15629 (.I(n18930), .ZN(n28501));
    INVX1 U15630 (.I(N4527), .ZN(N28502));
    NANDX1 U15631 (.A1(n23871), .A2(n16599), .ZN(n28503));
    NANDX1 U15632 (.A1(n19098), .A2(N11638), .ZN(N28504));
    INVX1 U15633 (.I(N2541), .ZN(N28505));
    NANDX1 U15634 (.A1(N4565), .A2(n14476), .ZN(n28506));
    NANDX1 U15635 (.A1(n20250), .A2(N9928), .ZN(n28507));
    NOR2X1 U15636 (.A1(n13244), .A2(N2481), .ZN(n28508));
    NANDX1 U15637 (.A1(N4641), .A2(N1800), .ZN(N28509));
    NANDX1 U15638 (.A1(n16188), .A2(n21237), .ZN(n28510));
    NANDX1 U15639 (.A1(N11992), .A2(N6787), .ZN(n28511));
    NOR2X1 U15640 (.A1(n23883), .A2(n14484), .ZN(n28512));
    NOR2X1 U15641 (.A1(N2907), .A2(n25405), .ZN(n28513));
    NANDX1 U15642 (.A1(N8273), .A2(n24691), .ZN(n28514));
    NANDX1 U15643 (.A1(n19911), .A2(n19507), .ZN(n28515));
    NANDX1 U15644 (.A1(n16287), .A2(n24072), .ZN(n28516));
    NOR2X1 U15645 (.A1(N8682), .A2(n18819), .ZN(N28517));
    INVX1 U15646 (.I(N9247), .ZN(N28518));
    NANDX1 U15647 (.A1(N7038), .A2(N8128), .ZN(N28519));
    INVX1 U15648 (.I(n23107), .ZN(n28520));
    INVX1 U15649 (.I(n16156), .ZN(n28521));
    INVX1 U15650 (.I(N1728), .ZN(n28522));
    INVX1 U15651 (.I(N3163), .ZN(n28523));
    NANDX1 U15652 (.A1(n15295), .A2(N6415), .ZN(N28524));
    INVX1 U15653 (.I(N6970), .ZN(N28525));
    NOR2X1 U15654 (.A1(N8641), .A2(n15242), .ZN(n28526));
    NANDX1 U15655 (.A1(n22989), .A2(n23920), .ZN(N28527));
    NOR2X1 U15656 (.A1(n14375), .A2(n14704), .ZN(n28528));
    NANDX1 U15657 (.A1(N9004), .A2(n23385), .ZN(n28529));
    NOR2X1 U15658 (.A1(n13560), .A2(n21400), .ZN(N28530));
    NANDX1 U15659 (.A1(N9365), .A2(n18295), .ZN(n28531));
    NOR2X1 U15660 (.A1(n21240), .A2(n24112), .ZN(n28532));
    NOR2X1 U15661 (.A1(n17616), .A2(N338), .ZN(N28533));
    INVX1 U15662 (.I(n20779), .ZN(N28534));
    INVX1 U15663 (.I(n15628), .ZN(N28535));
    NANDX1 U15664 (.A1(n22041), .A2(N11365), .ZN(N28536));
    NANDX1 U15665 (.A1(n19449), .A2(n15374), .ZN(n28537));
    NOR2X1 U15666 (.A1(n16935), .A2(n13792), .ZN(n28538));
    INVX1 U15667 (.I(N5807), .ZN(N28539));
    NOR2X1 U15668 (.A1(n20214), .A2(n14810), .ZN(n28540));
    NANDX1 U15669 (.A1(N3415), .A2(n17137), .ZN(N28541));
    INVX1 U15670 (.I(n18676), .ZN(N28542));
    INVX1 U15671 (.I(n18105), .ZN(N28543));
    NOR2X1 U15672 (.A1(N11007), .A2(n16715), .ZN(n28544));
    NOR2X1 U15673 (.A1(N3120), .A2(N5820), .ZN(n28545));
    INVX1 U15674 (.I(n23898), .ZN(n28546));
    NOR2X1 U15675 (.A1(n22051), .A2(n14356), .ZN(n28547));
    NOR2X1 U15676 (.A1(N7913), .A2(N11131), .ZN(n28548));
    NOR2X1 U15677 (.A1(n23286), .A2(n16448), .ZN(N28549));
    NANDX1 U15678 (.A1(N11575), .A2(n24313), .ZN(N28550));
    INVX1 U15679 (.I(N3336), .ZN(n28551));
    NOR2X1 U15680 (.A1(n20039), .A2(N7249), .ZN(N28552));
    NANDX1 U15681 (.A1(N11674), .A2(N7059), .ZN(n28553));
    NOR2X1 U15682 (.A1(N12673), .A2(n25163), .ZN(n28554));
    INVX1 U15683 (.I(N12447), .ZN(n28555));
    NANDX1 U15684 (.A1(n18873), .A2(n15566), .ZN(n28556));
    INVX1 U15685 (.I(N11026), .ZN(n28557));
    NOR2X1 U15686 (.A1(n14200), .A2(n21844), .ZN(N28558));
    NOR2X1 U15687 (.A1(N2743), .A2(N4254), .ZN(n28559));
    NOR2X1 U15688 (.A1(n21967), .A2(n16308), .ZN(n28560));
    INVX1 U15689 (.I(n21390), .ZN(n28561));
    NANDX1 U15690 (.A1(n21009), .A2(N1118), .ZN(N28562));
    NANDX1 U15691 (.A1(N3299), .A2(n21156), .ZN(N28563));
    NANDX1 U15692 (.A1(n14505), .A2(N7327), .ZN(n28564));
    INVX1 U15693 (.I(n18885), .ZN(n28565));
    NANDX1 U15694 (.A1(N11488), .A2(n20435), .ZN(n28566));
    NOR2X1 U15695 (.A1(n16630), .A2(N2573), .ZN(n28567));
    INVX1 U15696 (.I(n16360), .ZN(n28568));
    INVX1 U15697 (.I(N2774), .ZN(n28569));
    NANDX1 U15698 (.A1(n24210), .A2(N8626), .ZN(n28570));
    NANDX1 U15699 (.A1(n17232), .A2(n14377), .ZN(n28571));
    NOR2X1 U15700 (.A1(N8037), .A2(N11073), .ZN(n28572));
    NOR2X1 U15701 (.A1(n13454), .A2(n20849), .ZN(N28573));
    NANDX1 U15702 (.A1(n22207), .A2(n24148), .ZN(n28574));
    NOR2X1 U15703 (.A1(N12705), .A2(N1918), .ZN(n28575));
    NOR2X1 U15704 (.A1(N10262), .A2(n20802), .ZN(N28576));
    NANDX1 U15705 (.A1(N10517), .A2(N4502), .ZN(n28577));
    NANDX1 U15706 (.A1(N1644), .A2(N7075), .ZN(n28578));
    NOR2X1 U15707 (.A1(N6771), .A2(n23711), .ZN(N28579));
    NANDX1 U15708 (.A1(n14865), .A2(n22418), .ZN(N28580));
    NANDX1 U15709 (.A1(N11432), .A2(N2915), .ZN(n28581));
    NANDX1 U15710 (.A1(N7500), .A2(n25221), .ZN(n28582));
    NOR2X1 U15711 (.A1(n24958), .A2(n13173), .ZN(N28583));
    NANDX1 U15712 (.A1(n18031), .A2(N9877), .ZN(N28584));
    NANDX1 U15713 (.A1(N6758), .A2(n22581), .ZN(n28585));
    INVX1 U15714 (.I(n17081), .ZN(n28586));
    NOR2X1 U15715 (.A1(N12242), .A2(N10668), .ZN(n28587));
    NOR2X1 U15716 (.A1(n16743), .A2(n14236), .ZN(n28588));
    INVX1 U15717 (.I(N12585), .ZN(n28589));
    NANDX1 U15718 (.A1(n18076), .A2(N10793), .ZN(n28590));
    INVX1 U15719 (.I(N7439), .ZN(N28591));
    NANDX1 U15720 (.A1(n16780), .A2(N7638), .ZN(N28592));
    NANDX1 U15721 (.A1(N9432), .A2(n15137), .ZN(N28593));
    INVX1 U15722 (.I(N1925), .ZN(n28594));
    NANDX1 U15723 (.A1(N12282), .A2(N4034), .ZN(N28595));
    INVX1 U15724 (.I(n22158), .ZN(n28596));
    INVX1 U15725 (.I(n16916), .ZN(N28597));
    NOR2X1 U15726 (.A1(N7459), .A2(N8494), .ZN(N28598));
    NOR2X1 U15727 (.A1(N8468), .A2(N7930), .ZN(n28599));
    NOR2X1 U15728 (.A1(n25211), .A2(n22165), .ZN(n28600));
    INVX1 U15729 (.I(N1061), .ZN(n28601));
    NOR2X1 U15730 (.A1(N3382), .A2(N11854), .ZN(n28602));
    INVX1 U15731 (.I(N10820), .ZN(n28603));
    NOR2X1 U15732 (.A1(N7556), .A2(n18457), .ZN(N28604));
    NANDX1 U15733 (.A1(n16988), .A2(n22361), .ZN(N28605));
    NANDX1 U15734 (.A1(N7680), .A2(n14489), .ZN(n28606));
    NOR2X1 U15735 (.A1(N11713), .A2(n24648), .ZN(N28607));
    NANDX1 U15736 (.A1(N5268), .A2(n16061), .ZN(N28608));
    NANDX1 U15737 (.A1(N1494), .A2(n13323), .ZN(N28609));
    NANDX1 U15738 (.A1(N9962), .A2(N10020), .ZN(n28610));
    NANDX1 U15739 (.A1(n23940), .A2(N6682), .ZN(n28611));
    NOR2X1 U15740 (.A1(n25000), .A2(N9960), .ZN(N28612));
    NANDX1 U15741 (.A1(N119), .A2(N737), .ZN(N28613));
    NOR2X1 U15742 (.A1(N8448), .A2(n22562), .ZN(n28614));
    INVX1 U15743 (.I(N4936), .ZN(n28615));
    NOR2X1 U15744 (.A1(n14582), .A2(n14802), .ZN(n28616));
    INVX1 U15745 (.I(N3569), .ZN(n28617));
    NOR2X1 U15746 (.A1(N10974), .A2(N2714), .ZN(n28618));
    NANDX1 U15747 (.A1(N5009), .A2(N7542), .ZN(n28619));
    INVX1 U15748 (.I(N6503), .ZN(n28620));
    NANDX1 U15749 (.A1(N3273), .A2(n16464), .ZN(N28621));
    NOR2X1 U15750 (.A1(N11229), .A2(n14901), .ZN(n28622));
    INVX1 U15751 (.I(n18760), .ZN(N28623));
    NANDX1 U15752 (.A1(n25060), .A2(N4170), .ZN(N28624));
    NANDX1 U15753 (.A1(n14564), .A2(N399), .ZN(n28625));
    INVX1 U15754 (.I(N11624), .ZN(N28626));
    NOR2X1 U15755 (.A1(N5435), .A2(n14438), .ZN(n28627));
    INVX1 U15756 (.I(N9005), .ZN(n28628));
    INVX1 U15757 (.I(N10769), .ZN(n28629));
    NANDX1 U15758 (.A1(n13441), .A2(N2250), .ZN(n28630));
    NOR2X1 U15759 (.A1(n18450), .A2(N9792), .ZN(n28631));
    INVX1 U15760 (.I(n24952), .ZN(N28632));
    NOR2X1 U15761 (.A1(N12059), .A2(N4681), .ZN(n28633));
    NOR2X1 U15762 (.A1(N12055), .A2(N8349), .ZN(n28634));
    INVX1 U15763 (.I(N5312), .ZN(n28635));
    NANDX1 U15764 (.A1(n16997), .A2(N9481), .ZN(n28636));
    NOR2X1 U15765 (.A1(n20329), .A2(n24149), .ZN(n28637));
    INVX1 U15766 (.I(N6450), .ZN(N28638));
    INVX1 U15767 (.I(N9500), .ZN(n28639));
    NOR2X1 U15768 (.A1(n23969), .A2(n18504), .ZN(n28640));
    INVX1 U15769 (.I(n23505), .ZN(N28641));
    INVX1 U15770 (.I(n14331), .ZN(n28642));
    NANDX1 U15771 (.A1(N1918), .A2(N7278), .ZN(n28643));
    NANDX1 U15772 (.A1(N10704), .A2(n20997), .ZN(n28644));
    NANDX1 U15773 (.A1(n22762), .A2(n14445), .ZN(n28645));
    INVX1 U15774 (.I(N9315), .ZN(n28646));
    NOR2X1 U15775 (.A1(n23742), .A2(n14626), .ZN(N28647));
    NANDX1 U15776 (.A1(n15237), .A2(n12875), .ZN(N28648));
    NANDX1 U15777 (.A1(n24333), .A2(N11521), .ZN(n28649));
    NOR2X1 U15778 (.A1(N5280), .A2(n17057), .ZN(n28650));
    INVX1 U15779 (.I(N3702), .ZN(n28651));
    NANDX1 U15780 (.A1(N7704), .A2(N4592), .ZN(n28652));
    NOR2X1 U15781 (.A1(N9924), .A2(n18922), .ZN(n28653));
    INVX1 U15782 (.I(N11841), .ZN(n28654));
    NOR2X1 U15783 (.A1(N12588), .A2(n22544), .ZN(n28655));
    NOR2X1 U15784 (.A1(N5320), .A2(N8572), .ZN(n28656));
    NANDX1 U15785 (.A1(N390), .A2(n17886), .ZN(n28657));
    NANDX1 U15786 (.A1(n12900), .A2(n21279), .ZN(N28658));
    NOR2X1 U15787 (.A1(n16904), .A2(n22921), .ZN(n28659));
    NANDX1 U15788 (.A1(n15734), .A2(n23210), .ZN(n28660));
    INVX1 U15789 (.I(N9781), .ZN(N28661));
    NANDX1 U15790 (.A1(n15305), .A2(N2250), .ZN(n28662));
    NOR2X1 U15791 (.A1(N11776), .A2(N6841), .ZN(n28663));
    NOR2X1 U15792 (.A1(n21699), .A2(n14530), .ZN(n28664));
    NANDX1 U15793 (.A1(N8038), .A2(N3994), .ZN(n28665));
    INVX1 U15794 (.I(n19349), .ZN(N28666));
    NANDX1 U15795 (.A1(n16295), .A2(N2418), .ZN(n28667));
    INVX1 U15796 (.I(N5453), .ZN(n28668));
    INVX1 U15797 (.I(N5392), .ZN(n28669));
    NOR2X1 U15798 (.A1(n19118), .A2(n16964), .ZN(N28670));
    INVX1 U15799 (.I(n16536), .ZN(N28671));
    INVX1 U15800 (.I(n14254), .ZN(N28672));
    INVX1 U15801 (.I(n19043), .ZN(n28673));
    NANDX1 U15802 (.A1(N3504), .A2(N8845), .ZN(n28674));
    NANDX1 U15803 (.A1(n22557), .A2(N9388), .ZN(n28675));
    NOR2X1 U15804 (.A1(N4131), .A2(N5584), .ZN(N28676));
    NOR2X1 U15805 (.A1(n13751), .A2(N2389), .ZN(n28677));
    INVX1 U15806 (.I(n24726), .ZN(n28678));
    INVX1 U15807 (.I(n21172), .ZN(n28679));
    NANDX1 U15808 (.A1(n12923), .A2(n15602), .ZN(n28680));
    NANDX1 U15809 (.A1(N10762), .A2(N9761), .ZN(n28681));
    NANDX1 U15810 (.A1(N4377), .A2(N1222), .ZN(n28682));
    NOR2X1 U15811 (.A1(n20912), .A2(N5392), .ZN(N28683));
    NANDX1 U15812 (.A1(n23923), .A2(n24434), .ZN(n28684));
    NOR2X1 U15813 (.A1(n16194), .A2(n22046), .ZN(n28685));
    NANDX1 U15814 (.A1(n13249), .A2(N5931), .ZN(n28686));
    NANDX1 U15815 (.A1(N6147), .A2(N282), .ZN(n28687));
    NANDX1 U15816 (.A1(N8665), .A2(N2671), .ZN(n28688));
    NOR2X1 U15817 (.A1(N7888), .A2(n13176), .ZN(n28689));
    NANDX1 U15818 (.A1(N942), .A2(n14866), .ZN(n28690));
    NOR2X1 U15819 (.A1(N10680), .A2(N125), .ZN(n28691));
    INVX1 U15820 (.I(N2035), .ZN(n28692));
    INVX1 U15821 (.I(n17254), .ZN(n28693));
    NOR2X1 U15822 (.A1(N2949), .A2(n22645), .ZN(N28694));
    INVX1 U15823 (.I(N1369), .ZN(n28695));
    NANDX1 U15824 (.A1(N1735), .A2(n17562), .ZN(N28696));
    NOR2X1 U15825 (.A1(N8213), .A2(n19578), .ZN(n28697));
    NOR2X1 U15826 (.A1(N11079), .A2(N222), .ZN(n28698));
    INVX1 U15827 (.I(n13632), .ZN(n28699));
    NOR2X1 U15828 (.A1(N4537), .A2(n19865), .ZN(N28700));
    NOR2X1 U15829 (.A1(n17712), .A2(N10536), .ZN(n28701));
    NOR2X1 U15830 (.A1(n21345), .A2(n16807), .ZN(n28702));
    NOR2X1 U15831 (.A1(N10238), .A2(n18569), .ZN(n28703));
    NOR2X1 U15832 (.A1(N3506), .A2(n24591), .ZN(n28704));
    NOR2X1 U15833 (.A1(N6454), .A2(n21733), .ZN(n28705));
    NOR2X1 U15834 (.A1(n22092), .A2(N6575), .ZN(n28706));
    INVX1 U15835 (.I(n14152), .ZN(N28707));
    NOR2X1 U15836 (.A1(N703), .A2(n22497), .ZN(n28708));
    NOR2X1 U15837 (.A1(N11781), .A2(N11487), .ZN(n28709));
    INVX1 U15838 (.I(n25413), .ZN(n28710));
    INVX1 U15839 (.I(N7178), .ZN(n28711));
    INVX1 U15840 (.I(N3449), .ZN(n28712));
    INVX1 U15841 (.I(n19078), .ZN(N28713));
    NOR2X1 U15842 (.A1(N9499), .A2(n24653), .ZN(n28714));
    NOR2X1 U15843 (.A1(n19736), .A2(N6487), .ZN(N28715));
    NANDX1 U15844 (.A1(N12010), .A2(N5575), .ZN(n28716));
    INVX1 U15845 (.I(N7231), .ZN(n28717));
    NOR2X1 U15846 (.A1(N12338), .A2(N3821), .ZN(n28718));
    NANDX1 U15847 (.A1(N4828), .A2(N6740), .ZN(n28719));
    NANDX1 U15848 (.A1(N5530), .A2(N3734), .ZN(n28720));
    INVX1 U15849 (.I(N6078), .ZN(n28721));
    NANDX1 U15850 (.A1(n17062), .A2(n20258), .ZN(N28722));
    NOR2X1 U15851 (.A1(n24239), .A2(N3299), .ZN(N28723));
    NOR2X1 U15852 (.A1(N12393), .A2(N11144), .ZN(n28724));
    NOR2X1 U15853 (.A1(N10660), .A2(N10294), .ZN(N28725));
    NANDX1 U15854 (.A1(n19163), .A2(n16781), .ZN(n28726));
    INVX1 U15855 (.I(n19940), .ZN(n28727));
    INVX1 U15856 (.I(n15227), .ZN(N28728));
    INVX1 U15857 (.I(n12928), .ZN(n28729));
    NANDX1 U15858 (.A1(N5489), .A2(n24345), .ZN(n28730));
    INVX1 U15859 (.I(N12228), .ZN(n28731));
    INVX1 U15860 (.I(N4224), .ZN(n28732));
    NOR2X1 U15861 (.A1(N12639), .A2(N10302), .ZN(N28733));
    NANDX1 U15862 (.A1(n18469), .A2(N5057), .ZN(N28734));
    NANDX1 U15863 (.A1(n17205), .A2(n22625), .ZN(N28735));
    INVX1 U15864 (.I(n18366), .ZN(N28736));
    NANDX1 U15865 (.A1(n13922), .A2(n17793), .ZN(n28737));
    INVX1 U15866 (.I(n14399), .ZN(n28738));
    NOR2X1 U15867 (.A1(n24108), .A2(n19276), .ZN(n28739));
    NANDX1 U15868 (.A1(N9729), .A2(n23271), .ZN(n28740));
    NOR2X1 U15869 (.A1(N11424), .A2(N2868), .ZN(n28741));
    INVX1 U15870 (.I(n24537), .ZN(n28742));
    NANDX1 U15871 (.A1(N2810), .A2(N11523), .ZN(n28743));
    NOR2X1 U15872 (.A1(n18770), .A2(n12929), .ZN(n28744));
    NOR2X1 U15873 (.A1(n13216), .A2(N5895), .ZN(N28745));
    NANDX1 U15874 (.A1(n20789), .A2(n23100), .ZN(n28746));
    NANDX1 U15875 (.A1(n19436), .A2(N4731), .ZN(n28747));
    INVX1 U15876 (.I(N7855), .ZN(N28748));
    NOR2X1 U15877 (.A1(N164), .A2(N11021), .ZN(n28749));
    NOR2X1 U15878 (.A1(n13039), .A2(N4795), .ZN(n28750));
    NANDX1 U15879 (.A1(N11535), .A2(n16833), .ZN(N28751));
    INVX1 U15880 (.I(N11727), .ZN(N28752));
    NANDX1 U15881 (.A1(N4309), .A2(N10761), .ZN(n28753));
    NOR2X1 U15882 (.A1(N7118), .A2(n22283), .ZN(n28754));
    NOR2X1 U15883 (.A1(n14656), .A2(N9709), .ZN(N28755));
    NOR2X1 U15884 (.A1(n16639), .A2(n15604), .ZN(n28756));
    NANDX1 U15885 (.A1(N11926), .A2(N1969), .ZN(n28757));
    INVX1 U15886 (.I(N5859), .ZN(n28758));
    NANDX1 U15887 (.A1(n19218), .A2(N2481), .ZN(N28759));
    INVX1 U15888 (.I(N8149), .ZN(n28760));
    INVX1 U15889 (.I(N3997), .ZN(n28761));
    NOR2X1 U15890 (.A1(N7063), .A2(n21398), .ZN(n28762));
    INVX1 U15891 (.I(n23895), .ZN(n28763));
    INVX1 U15892 (.I(N7714), .ZN(n28764));
    INVX1 U15893 (.I(N2699), .ZN(N28765));
    NANDX1 U15894 (.A1(n25084), .A2(n24086), .ZN(n28766));
    NANDX1 U15895 (.A1(N1127), .A2(n13239), .ZN(n28767));
    NANDX1 U15896 (.A1(N7527), .A2(N4376), .ZN(n28768));
    INVX1 U15897 (.I(N12605), .ZN(n28769));
    NOR2X1 U15898 (.A1(N8838), .A2(n13485), .ZN(n28770));
    INVX1 U15899 (.I(N4304), .ZN(n28771));
    NOR2X1 U15900 (.A1(N2175), .A2(N11060), .ZN(n28772));
    NOR2X1 U15901 (.A1(n15675), .A2(n15056), .ZN(n28773));
    NOR2X1 U15902 (.A1(n22738), .A2(n25221), .ZN(n28774));
    INVX1 U15903 (.I(n21130), .ZN(N28775));
    INVX1 U15904 (.I(N3503), .ZN(n28776));
    NANDX1 U15905 (.A1(N3845), .A2(n21977), .ZN(n28777));
    NOR2X1 U15906 (.A1(n16698), .A2(N496), .ZN(N28778));
    NOR2X1 U15907 (.A1(N4435), .A2(N2994), .ZN(n28779));
    INVX1 U15908 (.I(n23080), .ZN(N28780));
    INVX1 U15909 (.I(N863), .ZN(n28781));
    INVX1 U15910 (.I(n18700), .ZN(n28782));
    INVX1 U15911 (.I(n16610), .ZN(n28783));
    INVX1 U15912 (.I(N10315), .ZN(N28784));
    INVX1 U15913 (.I(n22830), .ZN(n28785));
    INVX1 U15914 (.I(n23226), .ZN(n28786));
    NOR2X1 U15915 (.A1(n14233), .A2(n20461), .ZN(n28787));
    NANDX1 U15916 (.A1(N10022), .A2(N4857), .ZN(n28788));
    NANDX1 U15917 (.A1(n13525), .A2(N7344), .ZN(n28789));
    NOR2X1 U15918 (.A1(n24269), .A2(n23683), .ZN(N28790));
    NOR2X1 U15919 (.A1(n13532), .A2(N4415), .ZN(N28791));
    INVX1 U15920 (.I(n16526), .ZN(N28792));
    INVX1 U15921 (.I(n16375), .ZN(n28793));
    NOR2X1 U15922 (.A1(n19036), .A2(N7788), .ZN(n28794));
    INVX1 U15923 (.I(n22151), .ZN(n28795));
    NOR2X1 U15924 (.A1(n17086), .A2(N6963), .ZN(n28796));
    NOR2X1 U15925 (.A1(n14414), .A2(n21394), .ZN(n28797));
    INVX1 U15926 (.I(n15565), .ZN(n28798));
    NANDX1 U15927 (.A1(n24630), .A2(N5202), .ZN(N28799));
    NOR2X1 U15928 (.A1(n18254), .A2(n21488), .ZN(N28800));
    NANDX1 U15929 (.A1(n14365), .A2(n16115), .ZN(n28801));
    NOR2X1 U15930 (.A1(N12546), .A2(n16208), .ZN(N28802));
    INVX1 U15931 (.I(n16960), .ZN(n28803));
    NOR2X1 U15932 (.A1(n14527), .A2(N9631), .ZN(n28804));
    INVX1 U15933 (.I(n15412), .ZN(n28805));
    NANDX1 U15934 (.A1(n19394), .A2(n23765), .ZN(N28806));
    NANDX1 U15935 (.A1(N7056), .A2(n15349), .ZN(n28807));
    NANDX1 U15936 (.A1(n13501), .A2(n18530), .ZN(n28808));
    NOR2X1 U15937 (.A1(n17670), .A2(n22862), .ZN(n28809));
    NANDX1 U15938 (.A1(N5565), .A2(n16831), .ZN(n28810));
    NANDX1 U15939 (.A1(n23818), .A2(N1584), .ZN(N28811));
    INVX1 U15940 (.I(N12680), .ZN(N28812));
    NOR2X1 U15941 (.A1(N991), .A2(n13993), .ZN(n28813));
    NOR2X1 U15942 (.A1(n24494), .A2(N5450), .ZN(N28814));
    NOR2X1 U15943 (.A1(N2286), .A2(N3849), .ZN(n28815));
    INVX1 U15944 (.I(N6466), .ZN(N28816));
    INVX1 U15945 (.I(N941), .ZN(n28817));
    NOR2X1 U15946 (.A1(n12901), .A2(N7996), .ZN(N28818));
    NOR2X1 U15947 (.A1(N11481), .A2(n21497), .ZN(n28819));
    INVX1 U15948 (.I(n20223), .ZN(n28820));
    INVX1 U15949 (.I(n13500), .ZN(n28821));
    NANDX1 U15950 (.A1(N7996), .A2(n19099), .ZN(n28822));
    NANDX1 U15951 (.A1(n20581), .A2(n20682), .ZN(n28823));
    NANDX1 U15952 (.A1(N7758), .A2(N1646), .ZN(N28824));
    NANDX1 U15953 (.A1(N10519), .A2(n24320), .ZN(n28825));
    INVX1 U15954 (.I(n15968), .ZN(N28826));
    NOR2X1 U15955 (.A1(N12189), .A2(N8584), .ZN(N28827));
    NOR2X1 U15956 (.A1(N7422), .A2(n18634), .ZN(n28828));
    NOR2X1 U15957 (.A1(N918), .A2(N6032), .ZN(N28829));
    NOR2X1 U15958 (.A1(N9761), .A2(n17513), .ZN(N28830));
    INVX1 U15959 (.I(n14670), .ZN(n28831));
    NANDX1 U15960 (.A1(N8669), .A2(N2667), .ZN(n28832));
    NANDX1 U15961 (.A1(n16664), .A2(N10533), .ZN(n28833));
    NOR2X1 U15962 (.A1(N11742), .A2(N5713), .ZN(N28834));
    NANDX1 U15963 (.A1(N8267), .A2(N7358), .ZN(N28835));
    INVX1 U15964 (.I(n18785), .ZN(n28836));
    INVX1 U15965 (.I(n13221), .ZN(n28837));
    INVX1 U15966 (.I(N434), .ZN(n28838));
    NANDX1 U15967 (.A1(N6602), .A2(n24206), .ZN(n28839));
    NOR2X1 U15968 (.A1(n25236), .A2(N12183), .ZN(n28840));
    NANDX1 U15969 (.A1(n20035), .A2(N8156), .ZN(n28841));
    NANDX1 U15970 (.A1(N12045), .A2(n14393), .ZN(n28842));
    NANDX1 U15971 (.A1(n13046), .A2(n23061), .ZN(n28843));
    NOR2X1 U15972 (.A1(N2131), .A2(N2990), .ZN(n28844));
    NANDX1 U15973 (.A1(n24388), .A2(n14731), .ZN(n28845));
    INVX1 U15974 (.I(n16794), .ZN(n28846));
    NANDX1 U15975 (.A1(n14016), .A2(n20111), .ZN(n28847));
    INVX1 U15976 (.I(n23229), .ZN(n28848));
    NOR2X1 U15977 (.A1(n17336), .A2(n23662), .ZN(N28849));
    INVX1 U15978 (.I(N12706), .ZN(n28850));
    INVX1 U15979 (.I(n21141), .ZN(N28851));
    NOR2X1 U15980 (.A1(N9046), .A2(N6923), .ZN(N28852));
    NOR2X1 U15981 (.A1(N5969), .A2(n16735), .ZN(N28853));
    NOR2X1 U15982 (.A1(n20362), .A2(N1444), .ZN(n28854));
    INVX1 U15983 (.I(n17920), .ZN(n28855));
    INVX1 U15984 (.I(N11727), .ZN(n28856));
    NANDX1 U15985 (.A1(n18305), .A2(n24882), .ZN(n28857));
    NOR2X1 U15986 (.A1(n24963), .A2(n16173), .ZN(N28858));
    INVX1 U15987 (.I(N2245), .ZN(n28859));
    INVX1 U15988 (.I(N7525), .ZN(n28860));
    INVX1 U15989 (.I(n21648), .ZN(n28861));
    INVX1 U15990 (.I(n23632), .ZN(N28862));
    INVX1 U15991 (.I(N831), .ZN(N28863));
    INVX1 U15992 (.I(n16829), .ZN(n28864));
    NOR2X1 U15993 (.A1(n18308), .A2(n23751), .ZN(n28865));
    NOR2X1 U15994 (.A1(n24276), .A2(n14983), .ZN(N28866));
    NANDX1 U15995 (.A1(N7903), .A2(N5194), .ZN(n28867));
    NANDX1 U15996 (.A1(n14591), .A2(N11320), .ZN(n28868));
    NANDX1 U15997 (.A1(n24268), .A2(N4123), .ZN(N28869));
    INVX1 U15998 (.I(N11941), .ZN(n28870));
    NANDX1 U15999 (.A1(n23006), .A2(N148), .ZN(n28871));
    NOR2X1 U16000 (.A1(N11322), .A2(N7672), .ZN(N28872));
    NOR2X1 U16001 (.A1(N7468), .A2(n21299), .ZN(n28873));
    NANDX1 U16002 (.A1(N3155), .A2(N10898), .ZN(n28874));
    NANDX1 U16003 (.A1(N8751), .A2(N1702), .ZN(N28875));
    NOR2X1 U16004 (.A1(n21269), .A2(n13747), .ZN(n28876));
    NOR2X1 U16005 (.A1(n25019), .A2(N11111), .ZN(n28877));
    NANDX1 U16006 (.A1(N4710), .A2(n18071), .ZN(n28878));
    NANDX1 U16007 (.A1(n16030), .A2(N11255), .ZN(N28879));
    NANDX1 U16008 (.A1(N8920), .A2(n18088), .ZN(n28880));
    INVX1 U16009 (.I(N12502), .ZN(N28881));
    INVX1 U16010 (.I(n18686), .ZN(n28882));
    NOR2X1 U16011 (.A1(n15681), .A2(N855), .ZN(N28883));
    NOR2X1 U16012 (.A1(N11916), .A2(N10922), .ZN(n28884));
    NANDX1 U16013 (.A1(n15070), .A2(n21819), .ZN(n28885));
    INVX1 U16014 (.I(N12589), .ZN(n28886));
    NOR2X1 U16015 (.A1(n16574), .A2(N8355), .ZN(N28887));
    INVX1 U16016 (.I(n24379), .ZN(n28888));
    NANDX1 U16017 (.A1(N11643), .A2(N3352), .ZN(n28889));
    INVX1 U16018 (.I(N4212), .ZN(N28890));
    INVX1 U16019 (.I(N6146), .ZN(n28891));
    NANDX1 U16020 (.A1(n14745), .A2(n15065), .ZN(n28892));
    NOR2X1 U16021 (.A1(N7781), .A2(N2065), .ZN(n28893));
    NOR2X1 U16022 (.A1(n15235), .A2(N9161), .ZN(n28894));
    NANDX1 U16023 (.A1(n16089), .A2(N10821), .ZN(n28895));
    NOR2X1 U16024 (.A1(n15778), .A2(n16408), .ZN(n28896));
    INVX1 U16025 (.I(N12094), .ZN(n28897));
    NOR2X1 U16026 (.A1(n22735), .A2(N10112), .ZN(N28898));
    NANDX1 U16027 (.A1(N5587), .A2(n24914), .ZN(N28899));
    NANDX1 U16028 (.A1(N2226), .A2(N11054), .ZN(N28900));
    NANDX1 U16029 (.A1(N3575), .A2(N4033), .ZN(n28901));
    NANDX1 U16030 (.A1(n23990), .A2(N8267), .ZN(N28902));
    INVX1 U16031 (.I(n13553), .ZN(N28903));
    NANDX1 U16032 (.A1(n17261), .A2(N4385), .ZN(n28904));
    INVX1 U16033 (.I(n21263), .ZN(n28905));
    NANDX1 U16034 (.A1(n17965), .A2(N618), .ZN(n28906));
    NANDX1 U16035 (.A1(N10003), .A2(n16395), .ZN(n28907));
    NANDX1 U16036 (.A1(n20149), .A2(N2987), .ZN(n28908));
    NOR2X1 U16037 (.A1(n17381), .A2(N1866), .ZN(n28909));
    INVX1 U16038 (.I(N11736), .ZN(n28910));
    INVX1 U16039 (.I(N11978), .ZN(n28911));
    NANDX1 U16040 (.A1(N1098), .A2(N6762), .ZN(n28912));
    NANDX1 U16041 (.A1(N5131), .A2(N12730), .ZN(n28913));
    NANDX1 U16042 (.A1(N2165), .A2(N7940), .ZN(n28914));
    NANDX1 U16043 (.A1(N10288), .A2(n13968), .ZN(n28915));
    NOR2X1 U16044 (.A1(n22626), .A2(N9729), .ZN(n28916));
    NANDX1 U16045 (.A1(n15088), .A2(N10346), .ZN(N28917));
    NOR2X1 U16046 (.A1(n13859), .A2(N1238), .ZN(N28918));
    NOR2X1 U16047 (.A1(N8505), .A2(n18494), .ZN(n28919));
    NANDX1 U16048 (.A1(n14654), .A2(N9127), .ZN(n28920));
    NANDX1 U16049 (.A1(N887), .A2(N10403), .ZN(n28921));
    INVX1 U16050 (.I(N3615), .ZN(n28922));
    NOR2X1 U16051 (.A1(n21740), .A2(N9918), .ZN(n28923));
    NOR2X1 U16052 (.A1(n23237), .A2(n14708), .ZN(N28924));
    NOR2X1 U16053 (.A1(n19944), .A2(n21818), .ZN(n28925));
    INVX1 U16054 (.I(N8409), .ZN(N28926));
    INVX1 U16055 (.I(n18011), .ZN(n28927));
    INVX1 U16056 (.I(N7346), .ZN(N28928));
    INVX1 U16057 (.I(N6018), .ZN(N28929));
    NANDX1 U16058 (.A1(N10223), .A2(n21526), .ZN(n28930));
    NANDX1 U16059 (.A1(n18727), .A2(n14517), .ZN(N28931));
    NOR2X1 U16060 (.A1(n22148), .A2(N12412), .ZN(N28932));
    NANDX1 U16061 (.A1(n23034), .A2(n22814), .ZN(n28933));
    NANDX1 U16062 (.A1(N1147), .A2(N11850), .ZN(N28934));
    NOR2X1 U16063 (.A1(n25334), .A2(N6016), .ZN(N28935));
    INVX1 U16064 (.I(n14539), .ZN(N28936));
    INVX1 U16065 (.I(n17374), .ZN(n28937));
    NOR2X1 U16066 (.A1(N12001), .A2(N281), .ZN(n28938));
    INVX1 U16067 (.I(N4510), .ZN(n28939));
    NOR2X1 U16068 (.A1(N506), .A2(N874), .ZN(N28940));
    NOR2X1 U16069 (.A1(n20519), .A2(N11096), .ZN(N28941));
    NANDX1 U16070 (.A1(N6235), .A2(n18590), .ZN(n28942));
    NANDX1 U16071 (.A1(n14179), .A2(n15236), .ZN(n28943));
    NOR2X1 U16072 (.A1(n25125), .A2(N1535), .ZN(n28944));
    NOR2X1 U16073 (.A1(n14314), .A2(n16951), .ZN(n28945));
    INVX1 U16074 (.I(n14011), .ZN(n28946));
    INVX1 U16075 (.I(N6402), .ZN(N28947));
    NOR2X1 U16076 (.A1(n20088), .A2(n23017), .ZN(n28948));
    INVX1 U16077 (.I(N5439), .ZN(n28949));
    INVX1 U16078 (.I(n17863), .ZN(n28950));
    NOR2X1 U16079 (.A1(N2793), .A2(n13815), .ZN(n28951));
    NANDX1 U16080 (.A1(N3666), .A2(N4553), .ZN(n28952));
    NANDX1 U16081 (.A1(N3529), .A2(N2546), .ZN(n28953));
    NANDX1 U16082 (.A1(N10886), .A2(n18094), .ZN(n28954));
    NOR2X1 U16083 (.A1(n14889), .A2(n20550), .ZN(N28955));
    NANDX1 U16084 (.A1(n16424), .A2(n20318), .ZN(n28956));
    NANDX1 U16085 (.A1(N7872), .A2(n20704), .ZN(n28957));
    NANDX1 U16086 (.A1(n13422), .A2(N1603), .ZN(n28958));
    INVX1 U16087 (.I(N8007), .ZN(n28959));
    NANDX1 U16088 (.A1(n15341), .A2(N2214), .ZN(n28960));
    NOR2X1 U16089 (.A1(N7701), .A2(n15082), .ZN(N28961));
    INVX1 U16090 (.I(N10284), .ZN(n28962));
    NOR2X1 U16091 (.A1(n18127), .A2(n14836), .ZN(n28963));
    INVX1 U16092 (.I(n21655), .ZN(n28964));
    NOR2X1 U16093 (.A1(N6542), .A2(n21309), .ZN(n28965));
    NANDX1 U16094 (.A1(n12880), .A2(N10695), .ZN(n28966));
    INVX1 U16095 (.I(N7609), .ZN(N28967));
    NANDX1 U16096 (.A1(N2874), .A2(N5419), .ZN(n28968));
    NOR2X1 U16097 (.A1(n23577), .A2(n17239), .ZN(n28969));
    NANDX1 U16098 (.A1(n13947), .A2(N3765), .ZN(n28970));
    NANDX1 U16099 (.A1(N1831), .A2(n19106), .ZN(N28971));
    NANDX1 U16100 (.A1(n24733), .A2(n15574), .ZN(N28972));
    NOR2X1 U16101 (.A1(n13692), .A2(N355), .ZN(n28973));
    NANDX1 U16102 (.A1(N6317), .A2(N3959), .ZN(n28974));
    NOR2X1 U16103 (.A1(n16739), .A2(N10108), .ZN(n28975));
    NANDX1 U16104 (.A1(N12545), .A2(n23118), .ZN(N28976));
    INVX1 U16105 (.I(n23240), .ZN(n28977));
    INVX1 U16106 (.I(n25180), .ZN(n28978));
    NANDX1 U16107 (.A1(N8546), .A2(n19366), .ZN(n28979));
    NANDX1 U16108 (.A1(n20890), .A2(N11102), .ZN(n28980));
    NOR2X1 U16109 (.A1(N9334), .A2(N3635), .ZN(n28981));
    NANDX1 U16110 (.A1(n25435), .A2(n22740), .ZN(n28982));
    INVX1 U16111 (.I(n13433), .ZN(n28983));
    NOR2X1 U16112 (.A1(n23485), .A2(N1622), .ZN(n28984));
    INVX1 U16113 (.I(n18487), .ZN(N28985));
    INVX1 U16114 (.I(n20162), .ZN(n28986));
    INVX1 U16115 (.I(n13445), .ZN(n28987));
    NANDX1 U16116 (.A1(N7060), .A2(N487), .ZN(n28988));
    NANDX1 U16117 (.A1(n24632), .A2(N12494), .ZN(n28989));
    NOR2X1 U16118 (.A1(n13077), .A2(N615), .ZN(n28990));
    NOR2X1 U16119 (.A1(N6941), .A2(n15530), .ZN(n28991));
    NANDX1 U16120 (.A1(N6810), .A2(n16620), .ZN(N28992));
    NOR2X1 U16121 (.A1(N10444), .A2(n14928), .ZN(n28993));
    NOR2X1 U16122 (.A1(n21951), .A2(N12667), .ZN(N28994));
    NOR2X1 U16123 (.A1(n23530), .A2(n24920), .ZN(n28995));
    INVX1 U16124 (.I(n14231), .ZN(n28996));
    NANDX1 U16125 (.A1(n24818), .A2(n23160), .ZN(n28997));
    INVX1 U16126 (.I(N12760), .ZN(n28998));
    INVX1 U16127 (.I(n16099), .ZN(n28999));
    INVX1 U16128 (.I(N10881), .ZN(n29000));
    NOR2X1 U16129 (.A1(n14508), .A2(n21972), .ZN(N29001));
    NOR2X1 U16130 (.A1(n15122), .A2(n16107), .ZN(N29002));
    NOR2X1 U16131 (.A1(n19419), .A2(N5630), .ZN(N29003));
    NOR2X1 U16132 (.A1(N10536), .A2(n18756), .ZN(n29004));
    NANDX1 U16133 (.A1(n25463), .A2(N6312), .ZN(n29005));
    NOR2X1 U16134 (.A1(N1396), .A2(N7300), .ZN(n29006));
    NANDX1 U16135 (.A1(N813), .A2(n24179), .ZN(n29007));
    INVX1 U16136 (.I(n18716), .ZN(n29008));
    NANDX1 U16137 (.A1(n25164), .A2(N2253), .ZN(n29009));
    INVX1 U16138 (.I(n19393), .ZN(n29010));
    INVX1 U16139 (.I(N12765), .ZN(n29011));
    NANDX1 U16140 (.A1(n22347), .A2(N1770), .ZN(n29012));
    NANDX1 U16141 (.A1(n13917), .A2(N5659), .ZN(n29013));
    NOR2X1 U16142 (.A1(N12427), .A2(n25077), .ZN(n29014));
    NOR2X1 U16143 (.A1(n17747), .A2(N10111), .ZN(n29015));
    NOR2X1 U16144 (.A1(n22278), .A2(n24341), .ZN(n29016));
    NANDX1 U16145 (.A1(n23257), .A2(N234), .ZN(N29017));
    INVX1 U16146 (.I(n22264), .ZN(n29018));
    INVX1 U16147 (.I(n17284), .ZN(n29019));
    NOR2X1 U16148 (.A1(N8530), .A2(n15275), .ZN(N29020));
    NOR2X1 U16149 (.A1(n25052), .A2(n14794), .ZN(n29021));
    NANDX1 U16150 (.A1(N6669), .A2(N2056), .ZN(n29022));
    INVX1 U16151 (.I(n17784), .ZN(N29023));
    NANDX1 U16152 (.A1(N12599), .A2(N6198), .ZN(n29024));
    NOR2X1 U16153 (.A1(N4443), .A2(N7393), .ZN(n29025));
    NOR2X1 U16154 (.A1(n16187), .A2(n25139), .ZN(n29026));
    INVX1 U16155 (.I(N6913), .ZN(n29027));
    INVX1 U16156 (.I(N9812), .ZN(n29028));
    INVX1 U16157 (.I(N8436), .ZN(N29029));
    INVX1 U16158 (.I(N93), .ZN(n29030));
    NOR2X1 U16159 (.A1(n14129), .A2(n17376), .ZN(n29031));
    NOR2X1 U16160 (.A1(n22658), .A2(n21419), .ZN(n29032));
    NANDX1 U16161 (.A1(N10975), .A2(N10710), .ZN(n29033));
    INVX1 U16162 (.I(N6412), .ZN(N29034));
    NANDX1 U16163 (.A1(n23373), .A2(n24195), .ZN(n29035));
    INVX1 U16164 (.I(N10469), .ZN(n29036));
    INVX1 U16165 (.I(n17877), .ZN(n29037));
    INVX1 U16166 (.I(N1050), .ZN(n29038));
    NOR2X1 U16167 (.A1(n19866), .A2(n14956), .ZN(n29039));
    NANDX1 U16168 (.A1(n15546), .A2(N135), .ZN(n29040));
    NANDX1 U16169 (.A1(n22534), .A2(N8571), .ZN(n29041));
    NANDX1 U16170 (.A1(n22627), .A2(N2535), .ZN(N29042));
    INVX1 U16171 (.I(N3268), .ZN(n29043));
    NOR2X1 U16172 (.A1(n24116), .A2(n13454), .ZN(n29044));
    NANDX1 U16173 (.A1(N9589), .A2(n24163), .ZN(N29045));
    NOR2X1 U16174 (.A1(n16000), .A2(n14463), .ZN(n29046));
    NOR2X1 U16175 (.A1(N3460), .A2(N8587), .ZN(n29047));
    NOR2X1 U16176 (.A1(n22619), .A2(n15231), .ZN(n29048));
    INVX1 U16177 (.I(N12437), .ZN(n29049));
    INVX1 U16178 (.I(N10894), .ZN(n29050));
    INVX1 U16179 (.I(N9639), .ZN(n29051));
    NANDX1 U16180 (.A1(N2025), .A2(n23659), .ZN(n29052));
    INVX1 U16181 (.I(n24865), .ZN(N29053));
    NANDX1 U16182 (.A1(n23633), .A2(n16167), .ZN(N29054));
    INVX1 U16183 (.I(N1398), .ZN(n29055));
    NOR2X1 U16184 (.A1(n22293), .A2(n14852), .ZN(N29056));
    NANDX1 U16185 (.A1(n20649), .A2(N2280), .ZN(N29057));
    INVX1 U16186 (.I(n25416), .ZN(n29058));
    NOR2X1 U16187 (.A1(n12942), .A2(N3373), .ZN(N29059));
    INVX1 U16188 (.I(N11523), .ZN(N29060));
    NANDX1 U16189 (.A1(N3826), .A2(n13783), .ZN(n29061));
    INVX1 U16190 (.I(N12293), .ZN(N29062));
    INVX1 U16191 (.I(N3583), .ZN(n29063));
    INVX1 U16192 (.I(n14380), .ZN(n29064));
    INVX1 U16193 (.I(N8855), .ZN(n29065));
    NOR2X1 U16194 (.A1(N8007), .A2(N5573), .ZN(n29066));
    NOR2X1 U16195 (.A1(n24174), .A2(n18020), .ZN(N29067));
    NOR2X1 U16196 (.A1(n24373), .A2(n14811), .ZN(N29068));
    NOR2X1 U16197 (.A1(n25263), .A2(n24227), .ZN(n29069));
    INVX1 U16198 (.I(n13358), .ZN(N29070));
    NOR2X1 U16199 (.A1(N820), .A2(n15067), .ZN(n29071));
    INVX1 U16200 (.I(N3685), .ZN(n29072));
    NOR2X1 U16201 (.A1(N5538), .A2(n21780), .ZN(N29073));
    INVX1 U16202 (.I(n21501), .ZN(N29074));
    INVX1 U16203 (.I(N2810), .ZN(n29075));
    NANDX1 U16204 (.A1(n19268), .A2(n17189), .ZN(N29076));
    NANDX1 U16205 (.A1(N2620), .A2(n18305), .ZN(N29077));
    INVX1 U16206 (.I(N8192), .ZN(n29078));
    NOR2X1 U16207 (.A1(N3672), .A2(n14980), .ZN(n29079));
    NANDX1 U16208 (.A1(N2542), .A2(n18558), .ZN(N29080));
    NANDX1 U16209 (.A1(N2302), .A2(n17282), .ZN(N29081));
    NOR2X1 U16210 (.A1(N4427), .A2(N4688), .ZN(n29082));
    INVX1 U16211 (.I(N8261), .ZN(n29083));
    NANDX1 U16212 (.A1(n17112), .A2(N9347), .ZN(n29084));
    INVX1 U16213 (.I(n13389), .ZN(n29085));
    INVX1 U16214 (.I(N41), .ZN(N29086));
    NANDX1 U16215 (.A1(n15792), .A2(n13892), .ZN(n29087));
    NOR2X1 U16216 (.A1(N7479), .A2(N10885), .ZN(n29088));
    NANDX1 U16217 (.A1(n14551), .A2(n15885), .ZN(n29089));
    NANDX1 U16218 (.A1(N6598), .A2(n19556), .ZN(n29090));
    NANDX1 U16219 (.A1(N2327), .A2(N10865), .ZN(n29091));
    NOR2X1 U16220 (.A1(n16587), .A2(N1935), .ZN(N29092));
    NOR2X1 U16221 (.A1(n14925), .A2(n20631), .ZN(n29093));
    NANDX1 U16222 (.A1(N2851), .A2(N3390), .ZN(n29094));
    INVX1 U16223 (.I(n19962), .ZN(N29095));
    NOR2X1 U16224 (.A1(N11116), .A2(N7849), .ZN(N29096));
    NANDX1 U16225 (.A1(N11156), .A2(n18574), .ZN(n29097));
    INVX1 U16226 (.I(n13815), .ZN(n29098));
    INVX1 U16227 (.I(n15292), .ZN(n29099));
    NANDX1 U16228 (.A1(n15904), .A2(N4340), .ZN(n29100));
    NOR2X1 U16229 (.A1(N5703), .A2(n25208), .ZN(n29101));
    NOR2X1 U16230 (.A1(n24751), .A2(n16302), .ZN(n29102));
    NOR2X1 U16231 (.A1(N11352), .A2(n21656), .ZN(N29103));
    NOR2X1 U16232 (.A1(N4003), .A2(n25349), .ZN(n29104));
    NANDX1 U16233 (.A1(N1341), .A2(N2697), .ZN(n29105));
    NANDX1 U16234 (.A1(N8415), .A2(N11426), .ZN(n29106));
    NANDX1 U16235 (.A1(n19530), .A2(N8042), .ZN(n29107));
    NOR2X1 U16236 (.A1(n19454), .A2(N1114), .ZN(n29108));
    INVX1 U16237 (.I(N7766), .ZN(n29109));
    NOR2X1 U16238 (.A1(N6424), .A2(n21233), .ZN(n29110));
    NANDX1 U16239 (.A1(n25034), .A2(n25083), .ZN(N29111));
    INVX1 U16240 (.I(n13507), .ZN(N29112));
    INVX1 U16241 (.I(N8298), .ZN(n29113));
    INVX1 U16242 (.I(N9289), .ZN(n29114));
    INVX1 U16243 (.I(n14729), .ZN(N29115));
    INVX1 U16244 (.I(N1188), .ZN(n29116));
    NOR2X1 U16245 (.A1(n20665), .A2(N2528), .ZN(n29117));
    NOR2X1 U16246 (.A1(n21690), .A2(n25212), .ZN(n29118));
    NOR2X1 U16247 (.A1(N1754), .A2(N8007), .ZN(n29119));
    INVX1 U16248 (.I(n21807), .ZN(n29120));
    NOR2X1 U16249 (.A1(n15387), .A2(n12939), .ZN(N29121));
    NOR2X1 U16250 (.A1(n14062), .A2(n19362), .ZN(n29122));
    NOR2X1 U16251 (.A1(N3139), .A2(N7661), .ZN(N29123));
    INVX1 U16252 (.I(N12188), .ZN(N29124));
    NANDX1 U16253 (.A1(N5555), .A2(N9253), .ZN(n29125));
    NANDX1 U16254 (.A1(n14844), .A2(n17670), .ZN(N29126));
    NANDX1 U16255 (.A1(N1138), .A2(n18857), .ZN(N29127));
    INVX1 U16256 (.I(n21802), .ZN(N29128));
    NOR2X1 U16257 (.A1(n15886), .A2(N6757), .ZN(n29129));
    NANDX1 U16258 (.A1(N10886), .A2(N8510), .ZN(n29130));
    NOR2X1 U16259 (.A1(n13927), .A2(n19084), .ZN(n29131));
    NOR2X1 U16260 (.A1(N3812), .A2(n20790), .ZN(n29132));
    NANDX1 U16261 (.A1(N6641), .A2(n14650), .ZN(n29133));
    NANDX1 U16262 (.A1(n24049), .A2(N11078), .ZN(n29134));
    NOR2X1 U16263 (.A1(N10734), .A2(n21013), .ZN(n29135));
    NANDX1 U16264 (.A1(n19987), .A2(N9750), .ZN(n29136));
    NANDX1 U16265 (.A1(N922), .A2(n16254), .ZN(N29137));
    NANDX1 U16266 (.A1(n19779), .A2(N599), .ZN(N29138));
    NANDX1 U16267 (.A1(n18698), .A2(N5252), .ZN(n29139));
    NOR2X1 U16268 (.A1(n17327), .A2(n16137), .ZN(N29140));
    NOR2X1 U16269 (.A1(N12730), .A2(N4561), .ZN(N29141));
    NOR2X1 U16270 (.A1(N10090), .A2(n22642), .ZN(N29142));
    NOR2X1 U16271 (.A1(N5942), .A2(n18051), .ZN(N29143));
    NANDX1 U16272 (.A1(N10285), .A2(n16597), .ZN(n29144));
    NANDX1 U16273 (.A1(N8429), .A2(N1829), .ZN(N29145));
    NOR2X1 U16274 (.A1(N12128), .A2(N10583), .ZN(n29146));
    NOR2X1 U16275 (.A1(n19438), .A2(N11504), .ZN(n29147));
    NANDX1 U16276 (.A1(n16653), .A2(n20050), .ZN(n29148));
    NOR2X1 U16277 (.A1(n24437), .A2(n13246), .ZN(n29149));
    INVX1 U16278 (.I(n13475), .ZN(n29150));
    INVX1 U16279 (.I(n24984), .ZN(n29151));
    NOR2X1 U16280 (.A1(N6567), .A2(n18312), .ZN(N29152));
    NOR2X1 U16281 (.A1(n16656), .A2(N4220), .ZN(n29153));
    NOR2X1 U16282 (.A1(N11365), .A2(n22270), .ZN(n29154));
    NANDX1 U16283 (.A1(n21649), .A2(n13364), .ZN(N29155));
    INVX1 U16284 (.I(N4576), .ZN(n29156));
    INVX1 U16285 (.I(n19464), .ZN(n29157));
    NOR2X1 U16286 (.A1(n14542), .A2(n17440), .ZN(n29158));
    NOR2X1 U16287 (.A1(n14814), .A2(n20438), .ZN(n29159));
    INVX1 U16288 (.I(N9361), .ZN(n29160));
    NOR2X1 U16289 (.A1(n18032), .A2(N11374), .ZN(N29161));
    NOR2X1 U16290 (.A1(n20274), .A2(N5211), .ZN(n29162));
    NANDX1 U16291 (.A1(N8832), .A2(N545), .ZN(n29163));
    NANDX1 U16292 (.A1(n17059), .A2(n17201), .ZN(n29164));
    NOR2X1 U16293 (.A1(n14741), .A2(n17333), .ZN(n29165));
    NOR2X1 U16294 (.A1(N5294), .A2(n13480), .ZN(N29166));
    INVX1 U16295 (.I(n25298), .ZN(n29167));
    INVX1 U16296 (.I(n24055), .ZN(n29168));
    NANDX1 U16297 (.A1(N1061), .A2(N1862), .ZN(n29169));
    NOR2X1 U16298 (.A1(n14737), .A2(n16675), .ZN(n29170));
    NANDX1 U16299 (.A1(N8332), .A2(n14804), .ZN(N29171));
    INVX1 U16300 (.I(n15131), .ZN(n29172));
    NANDX1 U16301 (.A1(N810), .A2(N9902), .ZN(n29173));
    NOR2X1 U16302 (.A1(N10707), .A2(n18734), .ZN(n29174));
    NOR2X1 U16303 (.A1(n13414), .A2(n24560), .ZN(n29175));
    INVX1 U16304 (.I(N9108), .ZN(n29176));
    INVX1 U16305 (.I(n18499), .ZN(N29177));
    NOR2X1 U16306 (.A1(N7859), .A2(n20746), .ZN(N29178));
    NANDX1 U16307 (.A1(N7654), .A2(n16336), .ZN(n29179));
    INVX1 U16308 (.I(N1410), .ZN(n29180));
    INVX1 U16309 (.I(N10845), .ZN(n29181));
    NANDX1 U16310 (.A1(N6631), .A2(N2018), .ZN(n29182));
    INVX1 U16311 (.I(N3730), .ZN(n29183));
    NANDX1 U16312 (.A1(N3973), .A2(n18860), .ZN(N29184));
    INVX1 U16313 (.I(n19052), .ZN(n29185));
    INVX1 U16314 (.I(n15186), .ZN(n29186));
    NANDX1 U16315 (.A1(n25030), .A2(N10384), .ZN(N29187));
    NOR2X1 U16316 (.A1(n24088), .A2(N317), .ZN(n29188));
    INVX1 U16317 (.I(N1151), .ZN(N29189));
    NOR2X1 U16318 (.A1(n17114), .A2(N9010), .ZN(n29190));
    NOR2X1 U16319 (.A1(n13275), .A2(n16663), .ZN(n29191));
    NOR2X1 U16320 (.A1(n22258), .A2(N6841), .ZN(N29192));
    INVX1 U16321 (.I(N7601), .ZN(n29193));
    INVX1 U16322 (.I(N6453), .ZN(N29194));
    NANDX1 U16323 (.A1(N7524), .A2(n24452), .ZN(n29195));
    INVX1 U16324 (.I(N264), .ZN(n29196));
    NOR2X1 U16325 (.A1(N10236), .A2(n19316), .ZN(n29197));
    NOR2X1 U16326 (.A1(n25422), .A2(N12340), .ZN(n29198));
    INVX1 U16327 (.I(n24573), .ZN(N29199));
    NANDX1 U16328 (.A1(N10986), .A2(n13657), .ZN(N29200));
    NANDX1 U16329 (.A1(N12136), .A2(n21240), .ZN(n29201));
    NANDX1 U16330 (.A1(N9913), .A2(N1601), .ZN(N29202));
    NOR2X1 U16331 (.A1(n15344), .A2(N9530), .ZN(N29203));
    NANDX1 U16332 (.A1(N10952), .A2(N9352), .ZN(N29204));
    INVX1 U16333 (.I(n22203), .ZN(n29205));
    INVX1 U16334 (.I(N5215), .ZN(N29206));
    INVX1 U16335 (.I(N3521), .ZN(n29207));
    INVX1 U16336 (.I(n18757), .ZN(n29208));
    NOR2X1 U16337 (.A1(n19423), .A2(N12570), .ZN(N29209));
    NANDX1 U16338 (.A1(n19342), .A2(n24909), .ZN(n29210));
    NOR2X1 U16339 (.A1(N7180), .A2(N6952), .ZN(n29211));
    NANDX1 U16340 (.A1(n20837), .A2(n15771), .ZN(n29212));
    NANDX1 U16341 (.A1(N5342), .A2(N4970), .ZN(N29213));
    NANDX1 U16342 (.A1(N6942), .A2(N7444), .ZN(n29214));
    NANDX1 U16343 (.A1(n16471), .A2(N6673), .ZN(N29215));
    INVX1 U16344 (.I(n14590), .ZN(n29216));
    INVX1 U16345 (.I(n17928), .ZN(n29217));
    INVX1 U16346 (.I(n21754), .ZN(N29218));
    NANDX1 U16347 (.A1(N217), .A2(N5439), .ZN(n29219));
    NANDX1 U16348 (.A1(n24583), .A2(n24861), .ZN(N29220));
    NANDX1 U16349 (.A1(n22050), .A2(N7469), .ZN(n29221));
    NANDX1 U16350 (.A1(n20684), .A2(N3416), .ZN(n29222));
    NOR2X1 U16351 (.A1(n16034), .A2(n24252), .ZN(n29223));
    NOR2X1 U16352 (.A1(N1055), .A2(n18361), .ZN(N29224));
    NANDX1 U16353 (.A1(n21490), .A2(n25303), .ZN(n29225));
    INVX1 U16354 (.I(N6265), .ZN(n29226));
    INVX1 U16355 (.I(N1796), .ZN(n29227));
    INVX1 U16356 (.I(N8397), .ZN(n29228));
    INVX1 U16357 (.I(n22956), .ZN(N29229));
    NANDX1 U16358 (.A1(N316), .A2(N8372), .ZN(n29230));
    NOR2X1 U16359 (.A1(n20024), .A2(N1313), .ZN(n29231));
    NOR2X1 U16360 (.A1(n19382), .A2(N6824), .ZN(n29232));
    NANDX1 U16361 (.A1(n15618), .A2(n14779), .ZN(n29233));
    INVX1 U16362 (.I(n19034), .ZN(N29234));
    INVX1 U16363 (.I(n15190), .ZN(n29235));
    NANDX1 U16364 (.A1(N9357), .A2(n16244), .ZN(n29236));
    NANDX1 U16365 (.A1(N8269), .A2(N999), .ZN(N29237));
    NOR2X1 U16366 (.A1(n14624), .A2(n21533), .ZN(n29238));
    NOR2X1 U16367 (.A1(n16419), .A2(N1059), .ZN(n29239));
    NANDX1 U16368 (.A1(N9251), .A2(n24014), .ZN(n29240));
    INVX1 U16369 (.I(n23836), .ZN(n29241));
    NOR2X1 U16370 (.A1(N11814), .A2(n18357), .ZN(n29242));
    INVX1 U16371 (.I(n16203), .ZN(n29243));
    NOR2X1 U16372 (.A1(n18057), .A2(N5908), .ZN(n29244));
    INVX1 U16373 (.I(N7333), .ZN(n29245));
    NOR2X1 U16374 (.A1(n24423), .A2(N11515), .ZN(n29246));
    INVX1 U16375 (.I(n19742), .ZN(n29247));
    NOR2X1 U16376 (.A1(n25264), .A2(n19151), .ZN(n29248));
    NANDX1 U16377 (.A1(n15030), .A2(N7128), .ZN(n29249));
    NOR2X1 U16378 (.A1(N11061), .A2(n14413), .ZN(n29250));
    NOR2X1 U16379 (.A1(N887), .A2(N4593), .ZN(n29251));
    NOR2X1 U16380 (.A1(n24900), .A2(n25367), .ZN(N29252));
    INVX1 U16381 (.I(n20550), .ZN(n29253));
    NANDX1 U16382 (.A1(n15692), .A2(n17513), .ZN(n29254));
    INVX1 U16383 (.I(n16696), .ZN(n29255));
    NANDX1 U16384 (.A1(N11323), .A2(n22086), .ZN(N29256));
    INVX1 U16385 (.I(N5154), .ZN(n29257));
    INVX1 U16386 (.I(n17681), .ZN(N29258));
    NOR2X1 U16387 (.A1(N4013), .A2(n16088), .ZN(n29259));
    NANDX1 U16388 (.A1(N11931), .A2(N8493), .ZN(n29260));
    NOR2X1 U16389 (.A1(N7826), .A2(N4289), .ZN(N29261));
    NOR2X1 U16390 (.A1(n22239), .A2(N5272), .ZN(n29262));
    NOR2X1 U16391 (.A1(n15599), .A2(n15506), .ZN(n29263));
    NOR2X1 U16392 (.A1(N4231), .A2(n24073), .ZN(n29264));
    NANDX1 U16393 (.A1(N4676), .A2(N3030), .ZN(n29265));
    NANDX1 U16394 (.A1(N10091), .A2(n19726), .ZN(n29266));
    NOR2X1 U16395 (.A1(n21414), .A2(N5077), .ZN(N29267));
    NANDX1 U16396 (.A1(n15335), .A2(N3618), .ZN(N29268));
    NOR2X1 U16397 (.A1(n15239), .A2(n21901), .ZN(N29269));
    INVX1 U16398 (.I(n17941), .ZN(n29270));
    INVX1 U16399 (.I(n15428), .ZN(n29271));
    INVX1 U16400 (.I(N4923), .ZN(n29272));
    INVX1 U16401 (.I(N2229), .ZN(N29273));
    NANDX1 U16402 (.A1(n24988), .A2(N6405), .ZN(n29274));
    NOR2X1 U16403 (.A1(N3759), .A2(n24248), .ZN(n29275));
    NANDX1 U16404 (.A1(n16599), .A2(N405), .ZN(n29276));
    NOR2X1 U16405 (.A1(n19629), .A2(N5306), .ZN(N29277));
    INVX1 U16406 (.I(N2620), .ZN(n29278));
    NANDX1 U16407 (.A1(n23969), .A2(N7696), .ZN(n29279));
    INVX1 U16408 (.I(n13802), .ZN(n29280));
    NANDX1 U16409 (.A1(N6754), .A2(n17808), .ZN(n29281));
    INVX1 U16410 (.I(n13689), .ZN(n29282));
    INVX1 U16411 (.I(N4808), .ZN(N29283));
    NOR2X1 U16412 (.A1(n20417), .A2(N9730), .ZN(n29284));
    INVX1 U16413 (.I(n22645), .ZN(n29285));
    NANDX1 U16414 (.A1(N352), .A2(n17818), .ZN(n29286));
    NANDX1 U16415 (.A1(N4111), .A2(N5331), .ZN(n29287));
    INVX1 U16416 (.I(n20709), .ZN(N29288));
    NOR2X1 U16417 (.A1(n23169), .A2(n14835), .ZN(n29289));
    NOR2X1 U16418 (.A1(N11454), .A2(n17454), .ZN(N29290));
    NOR2X1 U16419 (.A1(N9921), .A2(n13917), .ZN(N29291));
    NOR2X1 U16420 (.A1(N12490), .A2(n13998), .ZN(n29292));
    INVX1 U16421 (.I(N4795), .ZN(n29293));
    NOR2X1 U16422 (.A1(n22731), .A2(n15040), .ZN(n29294));
    NANDX1 U16423 (.A1(n15113), .A2(n24224), .ZN(n29295));
    NOR2X1 U16424 (.A1(N1709), .A2(N10135), .ZN(n29296));
    INVX1 U16425 (.I(N2060), .ZN(N29297));
    INVX1 U16426 (.I(N11920), .ZN(n29298));
    INVX1 U16427 (.I(n22050), .ZN(n29299));
    INVX1 U16428 (.I(n15647), .ZN(n29300));
    NOR2X1 U16429 (.A1(n17825), .A2(n19249), .ZN(N29301));
    NOR2X1 U16430 (.A1(n18047), .A2(n25471), .ZN(N29302));
    NANDX1 U16431 (.A1(n16735), .A2(N2653), .ZN(N29303));
    NANDX1 U16432 (.A1(N3722), .A2(n16650), .ZN(n29304));
    NOR2X1 U16433 (.A1(N8516), .A2(n15894), .ZN(n29305));
    NANDX1 U16434 (.A1(N12323), .A2(n19944), .ZN(N29306));
    NANDX1 U16435 (.A1(N11045), .A2(n22492), .ZN(N29307));
    INVX1 U16436 (.I(n21179), .ZN(n29308));
    NOR2X1 U16437 (.A1(n18950), .A2(N12396), .ZN(n29309));
    INVX1 U16438 (.I(n13887), .ZN(n29310));
    NANDX1 U16439 (.A1(N9306), .A2(n18301), .ZN(n29311));
    NANDX1 U16440 (.A1(N1629), .A2(N816), .ZN(N29312));
    NANDX1 U16441 (.A1(N8443), .A2(n15054), .ZN(n29313));
    INVX1 U16442 (.I(n13945), .ZN(n29314));
    NANDX1 U16443 (.A1(n12896), .A2(n17666), .ZN(n29315));
    NOR2X1 U16444 (.A1(N12700), .A2(n14949), .ZN(n29316));
    NOR2X1 U16445 (.A1(n24001), .A2(N1769), .ZN(n29317));
    NANDX1 U16446 (.A1(n24913), .A2(N12813), .ZN(n29318));
    NOR2X1 U16447 (.A1(n16300), .A2(n22759), .ZN(n29319));
    INVX1 U16448 (.I(N9747), .ZN(n29320));
    INVX1 U16449 (.I(N11092), .ZN(n29321));
    NANDX1 U16450 (.A1(N10401), .A2(n20397), .ZN(n29322));
    INVX1 U16451 (.I(N2199), .ZN(n29323));
    NANDX1 U16452 (.A1(n20285), .A2(n24627), .ZN(n29324));
    INVX1 U16453 (.I(N9836), .ZN(n29325));
    NOR2X1 U16454 (.A1(n21947), .A2(n16310), .ZN(n29326));
    NANDX1 U16455 (.A1(n14110), .A2(n13931), .ZN(n29327));
    INVX1 U16456 (.I(n17826), .ZN(N29328));
    NANDX1 U16457 (.A1(N424), .A2(n19595), .ZN(n29329));
    NOR2X1 U16458 (.A1(n25336), .A2(n21175), .ZN(n29330));
    INVX1 U16459 (.I(N4901), .ZN(n29331));
    NOR2X1 U16460 (.A1(n17361), .A2(n14648), .ZN(n29332));
    NOR2X1 U16461 (.A1(n17220), .A2(n15817), .ZN(n29333));
    INVX1 U16462 (.I(N882), .ZN(N29334));
    INVX1 U16463 (.I(N6986), .ZN(n29335));
    NANDX1 U16464 (.A1(N4567), .A2(n20380), .ZN(N29336));
    NOR2X1 U16465 (.A1(n14402), .A2(N4904), .ZN(n29337));
    NOR2X1 U16466 (.A1(N5209), .A2(N5362), .ZN(N29338));
    NOR2X1 U16467 (.A1(N7907), .A2(n18518), .ZN(n29339));
    INVX1 U16468 (.I(n24119), .ZN(n29340));
    INVX1 U16469 (.I(n19685), .ZN(N29341));
    NOR2X1 U16470 (.A1(N7542), .A2(N4125), .ZN(N29342));
    NOR2X1 U16471 (.A1(N1211), .A2(N11324), .ZN(n29343));
    NOR2X1 U16472 (.A1(n15858), .A2(n16943), .ZN(n29344));
    INVX1 U16473 (.I(N6172), .ZN(N29345));
    INVX1 U16474 (.I(n19965), .ZN(n29346));
    NOR2X1 U16475 (.A1(N6250), .A2(N6137), .ZN(n29347));
    INVX1 U16476 (.I(N1128), .ZN(N29348));
    NOR2X1 U16477 (.A1(N12459), .A2(n20301), .ZN(N29349));
    NANDX1 U16478 (.A1(N6435), .A2(N160), .ZN(N29350));
    INVX1 U16479 (.I(n14342), .ZN(n29351));
    NANDX1 U16480 (.A1(N4863), .A2(N1726), .ZN(n29352));
    NOR2X1 U16481 (.A1(n13315), .A2(N2046), .ZN(n29353));
    INVX1 U16482 (.I(n17440), .ZN(n29354));
    NANDX1 U16483 (.A1(N12674), .A2(N3261), .ZN(n29355));
    NANDX1 U16484 (.A1(n17299), .A2(N8971), .ZN(N29356));
    NOR2X1 U16485 (.A1(N12238), .A2(n19468), .ZN(N29357));
    INVX1 U16486 (.I(n16960), .ZN(n29358));
    INVX1 U16487 (.I(N8096), .ZN(n29359));
    NOR2X1 U16488 (.A1(N1342), .A2(N11445), .ZN(N29360));
    INVX1 U16489 (.I(n21643), .ZN(N29361));
    NOR2X1 U16490 (.A1(n19639), .A2(N10570), .ZN(N29362));
    NANDX1 U16491 (.A1(n22748), .A2(N6783), .ZN(n29363));
    NOR2X1 U16492 (.A1(n24474), .A2(N10705), .ZN(n29364));
    NANDX1 U16493 (.A1(N1017), .A2(n22168), .ZN(n29365));
    INVX1 U16494 (.I(n13069), .ZN(n29366));
    NANDX1 U16495 (.A1(N1096), .A2(N12714), .ZN(n29367));
    NANDX1 U16496 (.A1(N10067), .A2(N5941), .ZN(N29368));
    NOR2X1 U16497 (.A1(N4032), .A2(n19132), .ZN(N29369));
    INVX1 U16498 (.I(N4246), .ZN(N29370));
    NOR2X1 U16499 (.A1(N8613), .A2(n19858), .ZN(n29371));
    NANDX1 U16500 (.A1(n21817), .A2(N4766), .ZN(n29372));
    NANDX1 U16501 (.A1(N4722), .A2(N4103), .ZN(N29373));
    NOR2X1 U16502 (.A1(N1967), .A2(N10886), .ZN(n29374));
    INVX1 U16503 (.I(N938), .ZN(n29375));
    NANDX1 U16504 (.A1(n19055), .A2(n16225), .ZN(n29376));
    NOR2X1 U16505 (.A1(n16890), .A2(N3791), .ZN(n29377));
    NANDX1 U16506 (.A1(n17985), .A2(n16504), .ZN(N29378));
    INVX1 U16507 (.I(N2549), .ZN(N29379));
    NOR2X1 U16508 (.A1(n22672), .A2(n20850), .ZN(N29380));
    NOR2X1 U16509 (.A1(N5036), .A2(n25096), .ZN(N29381));
    INVX1 U16510 (.I(n13649), .ZN(n29382));
    INVX1 U16511 (.I(n22773), .ZN(n29383));
    NOR2X1 U16512 (.A1(n12984), .A2(n18890), .ZN(n29384));
    NANDX1 U16513 (.A1(n17086), .A2(N2729), .ZN(n29385));
    INVX1 U16514 (.I(n16739), .ZN(n29386));
    NOR2X1 U16515 (.A1(n20626), .A2(N12826), .ZN(N29387));
    NANDX1 U16516 (.A1(N11348), .A2(n19848), .ZN(n29388));
    NANDX1 U16517 (.A1(N3906), .A2(n24976), .ZN(n29389));
    NANDX1 U16518 (.A1(N9178), .A2(n20006), .ZN(N29390));
    INVX1 U16519 (.I(n20389), .ZN(n29391));
    INVX1 U16520 (.I(N8510), .ZN(n29392));
    INVX1 U16521 (.I(N10979), .ZN(n29393));
    NANDX1 U16522 (.A1(N9331), .A2(n24627), .ZN(n29394));
    NOR2X1 U16523 (.A1(N6601), .A2(n23357), .ZN(N29395));
    NOR2X1 U16524 (.A1(n14258), .A2(n15577), .ZN(N29396));
    INVX1 U16525 (.I(n16986), .ZN(n29397));
    NANDX1 U16526 (.A1(N3930), .A2(n21638), .ZN(n29398));
    NANDX1 U16527 (.A1(n16756), .A2(n19842), .ZN(n29399));
    NANDX1 U16528 (.A1(n25371), .A2(n23703), .ZN(n29400));
    NANDX1 U16529 (.A1(n24845), .A2(N8815), .ZN(n29401));
    NANDX1 U16530 (.A1(N8116), .A2(n21977), .ZN(n29402));
    NOR2X1 U16531 (.A1(n14059), .A2(n19254), .ZN(n29403));
    NOR2X1 U16532 (.A1(n25037), .A2(N4893), .ZN(N29404));
    INVX1 U16533 (.I(n12929), .ZN(n29405));
    NANDX1 U16534 (.A1(n20434), .A2(n25053), .ZN(n29406));
    NANDX1 U16535 (.A1(N9189), .A2(n15127), .ZN(n29407));
    NOR2X1 U16536 (.A1(n14943), .A2(n24889), .ZN(n29408));
    NOR2X1 U16537 (.A1(N11078), .A2(N4273), .ZN(n29409));
    NOR2X1 U16538 (.A1(n19688), .A2(N9274), .ZN(n29410));
    NANDX1 U16539 (.A1(N6656), .A2(N6948), .ZN(N29411));
    NANDX1 U16540 (.A1(n15470), .A2(n13800), .ZN(n29412));
    NANDX1 U16541 (.A1(N712), .A2(n15538), .ZN(n29413));
    INVX1 U16542 (.I(N8734), .ZN(N29414));
    NOR2X1 U16543 (.A1(n14956), .A2(n13626), .ZN(N29415));
    NOR2X1 U16544 (.A1(n16652), .A2(N12374), .ZN(n29416));
    NOR2X1 U16545 (.A1(N4971), .A2(N6730), .ZN(N29417));
    NOR2X1 U16546 (.A1(n20097), .A2(N2547), .ZN(n29418));
    NANDX1 U16547 (.A1(N8252), .A2(n13526), .ZN(n29419));
    NOR2X1 U16548 (.A1(N12524), .A2(N4525), .ZN(n29420));
    NANDX1 U16549 (.A1(N10565), .A2(N9663), .ZN(N29421));
    NOR2X1 U16550 (.A1(N6280), .A2(n14143), .ZN(n29422));
    INVX1 U16551 (.I(n20079), .ZN(n29423));
    INVX1 U16552 (.I(n24874), .ZN(n29424));
    NANDX1 U16553 (.A1(N5426), .A2(N8105), .ZN(n29425));
    NANDX1 U16554 (.A1(N9150), .A2(N10498), .ZN(N29426));
    NANDX1 U16555 (.A1(N299), .A2(N11640), .ZN(N29427));
    INVX1 U16556 (.I(N5269), .ZN(n29428));
    NOR2X1 U16557 (.A1(N12428), .A2(n14134), .ZN(N29429));
    NANDX1 U16558 (.A1(N6164), .A2(n22385), .ZN(n29430));
    INVX1 U16559 (.I(N10978), .ZN(n29431));
    NOR2X1 U16560 (.A1(n16501), .A2(n24247), .ZN(n29432));
    NOR2X1 U16561 (.A1(N662), .A2(n18670), .ZN(n29433));
    NANDX1 U16562 (.A1(n14804), .A2(n17330), .ZN(n29434));
    INVX1 U16563 (.I(n19078), .ZN(n29435));
    INVX1 U16564 (.I(N11513), .ZN(n29436));
    INVX1 U16565 (.I(n13574), .ZN(n29437));
    NANDX1 U16566 (.A1(N8151), .A2(n24071), .ZN(n29438));
    NOR2X1 U16567 (.A1(n22719), .A2(N10208), .ZN(N29439));
    NANDX1 U16568 (.A1(N2486), .A2(n17345), .ZN(n29440));
    NOR2X1 U16569 (.A1(N5387), .A2(N1526), .ZN(n29441));
    NOR2X1 U16570 (.A1(N2269), .A2(n24734), .ZN(n29442));
    NANDX1 U16571 (.A1(n14712), .A2(n15732), .ZN(n29443));
    NOR2X1 U16572 (.A1(N12217), .A2(N5161), .ZN(n29444));
    NOR2X1 U16573 (.A1(n16001), .A2(N8733), .ZN(n29445));
    NANDX1 U16574 (.A1(N3130), .A2(N2308), .ZN(n29446));
    INVX1 U16575 (.I(n14643), .ZN(N29447));
    INVX1 U16576 (.I(n22620), .ZN(N29448));
    INVX1 U16577 (.I(N9459), .ZN(n29449));
    NANDX1 U16578 (.A1(N9909), .A2(N6676), .ZN(n29450));
    INVX1 U16579 (.I(n19606), .ZN(n29451));
    NANDX1 U16580 (.A1(N774), .A2(n19266), .ZN(N29452));
    NANDX1 U16581 (.A1(N2299), .A2(n25090), .ZN(n29453));
    INVX1 U16582 (.I(n15800), .ZN(n29454));
    INVX1 U16583 (.I(n23332), .ZN(n29455));
    INVX1 U16584 (.I(N9470), .ZN(n29456));
    NOR2X1 U16585 (.A1(n25460), .A2(n21221), .ZN(n29457));
    NOR2X1 U16586 (.A1(N8690), .A2(n24798), .ZN(n29458));
    NANDX1 U16587 (.A1(N10997), .A2(n22612), .ZN(n29459));
    INVX1 U16588 (.I(N1074), .ZN(n29460));
    NOR2X1 U16589 (.A1(N4194), .A2(n24802), .ZN(N29461));
    NOR2X1 U16590 (.A1(n14102), .A2(n20245), .ZN(N29462));
    INVX1 U16591 (.I(n22476), .ZN(n29463));
    NOR2X1 U16592 (.A1(N2655), .A2(N5007), .ZN(n29464));
    INVX1 U16593 (.I(n19223), .ZN(n29465));
    INVX1 U16594 (.I(n18875), .ZN(N29466));
    INVX1 U16595 (.I(N9750), .ZN(n29467));
    NANDX1 U16596 (.A1(n18586), .A2(N7988), .ZN(n29468));
    INVX1 U16597 (.I(n18543), .ZN(N29469));
    NANDX1 U16598 (.A1(n16061), .A2(n16000), .ZN(n29470));
    INVX1 U16599 (.I(N8502), .ZN(N29471));
    NOR2X1 U16600 (.A1(n14381), .A2(n15585), .ZN(n29472));
    NANDX1 U16601 (.A1(n22877), .A2(N8546), .ZN(N29473));
    INVX1 U16602 (.I(n15827), .ZN(n29474));
    NANDX1 U16603 (.A1(n25150), .A2(n17708), .ZN(n29475));
    NOR2X1 U16604 (.A1(N6588), .A2(N9130), .ZN(N29476));
    NOR2X1 U16605 (.A1(N5611), .A2(N2850), .ZN(n29477));
    NOR2X1 U16606 (.A1(n13253), .A2(N1137), .ZN(N29478));
    NANDX1 U16607 (.A1(n18725), .A2(N8491), .ZN(n29479));
    NOR2X1 U16608 (.A1(N8739), .A2(n15801), .ZN(n29480));
    INVX1 U16609 (.I(n13567), .ZN(n29481));
    NOR2X1 U16610 (.A1(n23004), .A2(N10836), .ZN(N29482));
    NOR2X1 U16611 (.A1(N11882), .A2(n15188), .ZN(n29483));
    NANDX1 U16612 (.A1(n23527), .A2(n23733), .ZN(n29484));
    NANDX1 U16613 (.A1(n13851), .A2(n23916), .ZN(n29485));
    NOR2X1 U16614 (.A1(n20327), .A2(n21071), .ZN(n29486));
    NANDX1 U16615 (.A1(n18224), .A2(n23233), .ZN(n29487));
    INVX1 U16616 (.I(N9842), .ZN(N29488));
    NANDX1 U16617 (.A1(n23973), .A2(N10978), .ZN(n29489));
    NOR2X1 U16618 (.A1(N5963), .A2(N8236), .ZN(n29490));
    NANDX1 U16619 (.A1(N3470), .A2(n24037), .ZN(n29491));
    NOR2X1 U16620 (.A1(n17036), .A2(n19103), .ZN(n29492));
    INVX1 U16621 (.I(n16640), .ZN(N29493));
    NOR2X1 U16622 (.A1(n15672), .A2(N6325), .ZN(n29494));
    INVX1 U16623 (.I(n13696), .ZN(n29495));
    INVX1 U16624 (.I(N5471), .ZN(n29496));
    INVX1 U16625 (.I(N2969), .ZN(N29497));
    NOR2X1 U16626 (.A1(n25408), .A2(N12807), .ZN(N29498));
    NANDX1 U16627 (.A1(n18130), .A2(n24808), .ZN(N29499));
    NANDX1 U16628 (.A1(N2469), .A2(n18062), .ZN(n29500));
    INVX1 U16629 (.I(N2214), .ZN(N29501));
    NANDX1 U16630 (.A1(n24257), .A2(N10450), .ZN(n29502));
    NOR2X1 U16631 (.A1(N2224), .A2(n23254), .ZN(n29503));
    NOR2X1 U16632 (.A1(N8027), .A2(N5622), .ZN(n29504));
    NOR2X1 U16633 (.A1(n24666), .A2(n24322), .ZN(n29505));
    INVX1 U16634 (.I(N5489), .ZN(n29506));
    NANDX1 U16635 (.A1(N5583), .A2(N10044), .ZN(N29507));
    INVX1 U16636 (.I(N10665), .ZN(n29508));
    NANDX1 U16637 (.A1(N6684), .A2(N10570), .ZN(n29509));
    INVX1 U16638 (.I(N1517), .ZN(n29510));
    INVX1 U16639 (.I(N2659), .ZN(n29511));
    NOR2X1 U16640 (.A1(N5665), .A2(N9488), .ZN(n29512));
    NANDX1 U16641 (.A1(N7879), .A2(n14844), .ZN(n29513));
    NANDX1 U16642 (.A1(N7096), .A2(N6485), .ZN(n29514));
    NOR2X1 U16643 (.A1(N4847), .A2(n18684), .ZN(n29515));
    NANDX1 U16644 (.A1(n24738), .A2(N6133), .ZN(n29516));
    NOR2X1 U16645 (.A1(n23557), .A2(N12290), .ZN(n29517));
    NANDX1 U16646 (.A1(n20777), .A2(n17873), .ZN(n29518));
    INVX1 U16647 (.I(n23467), .ZN(n29519));
    INVX1 U16648 (.I(N2875), .ZN(N29520));
    NOR2X1 U16649 (.A1(N2372), .A2(n20498), .ZN(n29521));
    INVX1 U16650 (.I(N5569), .ZN(n29522));
    INVX1 U16651 (.I(n16273), .ZN(n29523));
    NOR2X1 U16652 (.A1(N7142), .A2(n16134), .ZN(n29524));
    INVX1 U16653 (.I(N10754), .ZN(n29525));
    NANDX1 U16654 (.A1(N3742), .A2(n17238), .ZN(n29526));
    NANDX1 U16655 (.A1(n22858), .A2(n24690), .ZN(N29527));
    INVX1 U16656 (.I(n22093), .ZN(n29528));
    NANDX1 U16657 (.A1(n13053), .A2(n20147), .ZN(N29529));
    NANDX1 U16658 (.A1(n15337), .A2(n15421), .ZN(N29530));
    NOR2X1 U16659 (.A1(n16432), .A2(N2154), .ZN(n29531));
    INVX1 U16660 (.I(N8074), .ZN(n29532));
    NOR2X1 U16661 (.A1(n18423), .A2(N3070), .ZN(N29533));
    INVX1 U16662 (.I(N12759), .ZN(N29534));
    NANDX1 U16663 (.A1(N9812), .A2(N12759), .ZN(n29535));
    NANDX1 U16664 (.A1(N443), .A2(N9406), .ZN(n29536));
    NOR2X1 U16665 (.A1(n18229), .A2(n13147), .ZN(N29537));
    NANDX1 U16666 (.A1(N11351), .A2(N10503), .ZN(N29538));
    NOR2X1 U16667 (.A1(n16376), .A2(N7093), .ZN(N29539));
    INVX1 U16668 (.I(N3926), .ZN(n29540));
    INVX1 U16669 (.I(N1810), .ZN(n29541));
    NOR2X1 U16670 (.A1(n20196), .A2(n14827), .ZN(n29542));
    NANDX1 U16671 (.A1(n22349), .A2(n19645), .ZN(N29543));
    NOR2X1 U16672 (.A1(N6686), .A2(N12565), .ZN(n29544));
    INVX1 U16673 (.I(N226), .ZN(n29545));
    NOR2X1 U16674 (.A1(N2632), .A2(N10037), .ZN(n29546));
    NANDX1 U16675 (.A1(n13534), .A2(n24750), .ZN(n29547));
    NANDX1 U16676 (.A1(N9688), .A2(n17476), .ZN(n29548));
    NANDX1 U16677 (.A1(N11847), .A2(n17595), .ZN(N29549));
    NANDX1 U16678 (.A1(N1961), .A2(n22738), .ZN(N29550));
    INVX1 U16679 (.I(n22896), .ZN(n29551));
    NANDX1 U16680 (.A1(N9535), .A2(n13473), .ZN(N29552));
    NANDX1 U16681 (.A1(N4228), .A2(n17067), .ZN(n29553));
    INVX1 U16682 (.I(n15345), .ZN(N29554));
    NANDX1 U16683 (.A1(N3952), .A2(N10798), .ZN(n29555));
    NANDX1 U16684 (.A1(n17092), .A2(N11023), .ZN(n29556));
    NANDX1 U16685 (.A1(n19723), .A2(n21060), .ZN(n29557));
    NOR2X1 U16686 (.A1(N7754), .A2(N9075), .ZN(N29558));
    NANDX1 U16687 (.A1(N6209), .A2(n15318), .ZN(n29559));
    NOR2X1 U16688 (.A1(N6823), .A2(N7410), .ZN(n29560));
    NOR2X1 U16689 (.A1(N8783), .A2(N4645), .ZN(n29561));
    NOR2X1 U16690 (.A1(n20446), .A2(n20076), .ZN(N29562));
    INVX1 U16691 (.I(n22687), .ZN(N29563));
    INVX1 U16692 (.I(n22657), .ZN(n29564));
    NOR2X1 U16693 (.A1(N682), .A2(N1267), .ZN(n29565));
    INVX1 U16694 (.I(n18903), .ZN(n29566));
    NANDX1 U16695 (.A1(N1268), .A2(N10492), .ZN(n29567));
    NOR2X1 U16696 (.A1(N2398), .A2(N4712), .ZN(N29568));
    NOR2X1 U16697 (.A1(n19145), .A2(N1234), .ZN(n29569));
    NOR2X1 U16698 (.A1(n21142), .A2(N7442), .ZN(N29570));
    NANDX1 U16699 (.A1(n24573), .A2(n14265), .ZN(N29571));
    INVX1 U16700 (.I(N169), .ZN(N29572));
    INVX1 U16701 (.I(n21394), .ZN(N29573));
    INVX1 U16702 (.I(N6759), .ZN(n29574));
    INVX1 U16703 (.I(n13223), .ZN(n29575));
    NANDX1 U16704 (.A1(N8498), .A2(n24648), .ZN(N29576));
    INVX1 U16705 (.I(n23450), .ZN(n29577));
    NOR2X1 U16706 (.A1(n21189), .A2(n16850), .ZN(n29578));
    INVX1 U16707 (.I(n22456), .ZN(N29579));
    NANDX1 U16708 (.A1(n13099), .A2(n24853), .ZN(n29580));
    NOR2X1 U16709 (.A1(N9278), .A2(N7263), .ZN(N29581));
    NANDX1 U16710 (.A1(N262), .A2(N2902), .ZN(n29582));
    NOR2X1 U16711 (.A1(n20833), .A2(N1972), .ZN(n29583));
    NANDX1 U16712 (.A1(N12079), .A2(n16411), .ZN(N29584));
    NANDX1 U16713 (.A1(N7970), .A2(n25474), .ZN(N29585));
    INVX1 U16714 (.I(N12704), .ZN(n29586));
    INVX1 U16715 (.I(N7076), .ZN(n29587));
    INVX1 U16716 (.I(N1108), .ZN(N29588));
    INVX1 U16717 (.I(N7917), .ZN(n29589));
    NANDX1 U16718 (.A1(n23993), .A2(n24766), .ZN(N29590));
    NOR2X1 U16719 (.A1(N9714), .A2(n15373), .ZN(n29591));
    NANDX1 U16720 (.A1(n23334), .A2(N10692), .ZN(n29592));
    NOR2X1 U16721 (.A1(N5094), .A2(N7243), .ZN(n29593));
    NANDX1 U16722 (.A1(n22265), .A2(N4), .ZN(N29594));
    NANDX1 U16723 (.A1(n13004), .A2(N7029), .ZN(n29595));
    INVX1 U16724 (.I(N3912), .ZN(n29596));
    NOR2X1 U16725 (.A1(N10119), .A2(N3884), .ZN(n29597));
    NOR2X1 U16726 (.A1(N11591), .A2(N5846), .ZN(n29598));
    NOR2X1 U16727 (.A1(n21560), .A2(n21223), .ZN(n29599));
    INVX1 U16728 (.I(n18244), .ZN(n29600));
    NANDX1 U16729 (.A1(N3676), .A2(N6275), .ZN(N29601));
    NANDX1 U16730 (.A1(n13389), .A2(n21648), .ZN(n29602));
    NOR2X1 U16731 (.A1(N11220), .A2(N6837), .ZN(n29603));
    NOR2X1 U16732 (.A1(n16313), .A2(N2847), .ZN(n29604));
    INVX1 U16733 (.I(N1843), .ZN(N29605));
    NOR2X1 U16734 (.A1(n15498), .A2(n14846), .ZN(N29606));
    NANDX1 U16735 (.A1(n17647), .A2(n18758), .ZN(n29607));
    INVX1 U16736 (.I(N2263), .ZN(n29608));
    NANDX1 U16737 (.A1(n16783), .A2(N2621), .ZN(n29609));
    NOR2X1 U16738 (.A1(n16126), .A2(n12948), .ZN(N29610));
    INVX1 U16739 (.I(n21311), .ZN(n29611));
    NOR2X1 U16740 (.A1(N2018), .A2(n24986), .ZN(n29612));
    NANDX1 U16741 (.A1(N11133), .A2(N12872), .ZN(n29613));
    NOR2X1 U16742 (.A1(n13643), .A2(N12859), .ZN(N29614));
    NANDX1 U16743 (.A1(n21865), .A2(n17939), .ZN(n29615));
    NANDX1 U16744 (.A1(n21790), .A2(n19781), .ZN(n29616));
    NANDX1 U16745 (.A1(N11785), .A2(N9124), .ZN(n29617));
    INVX1 U16746 (.I(N3929), .ZN(n29618));
    INVX1 U16747 (.I(N10106), .ZN(n29619));
    NANDX1 U16748 (.A1(n13787), .A2(N1386), .ZN(N29620));
    NANDX1 U16749 (.A1(n19808), .A2(N6279), .ZN(n29621));
    NOR2X1 U16750 (.A1(n21549), .A2(N2087), .ZN(n29622));
    INVX1 U16751 (.I(N12335), .ZN(n29623));
    NOR2X1 U16752 (.A1(N8753), .A2(n23467), .ZN(N29624));
    NOR2X1 U16753 (.A1(N5629), .A2(N11607), .ZN(n29625));
    INVX1 U16754 (.I(N12379), .ZN(n29626));
    INVX1 U16755 (.I(N8503), .ZN(N29627));
    NOR2X1 U16756 (.A1(n18527), .A2(N2781), .ZN(N29628));
    NANDX1 U16757 (.A1(n19079), .A2(N11905), .ZN(n29629));
    NANDX1 U16758 (.A1(N11775), .A2(N3051), .ZN(n29630));
    INVX1 U16759 (.I(n21003), .ZN(N29631));
    NANDX1 U16760 (.A1(N6002), .A2(N7350), .ZN(N29632));
    NOR2X1 U16761 (.A1(N1048), .A2(n20915), .ZN(N29633));
    NOR2X1 U16762 (.A1(N3135), .A2(N3434), .ZN(n29634));
    INVX1 U16763 (.I(N4704), .ZN(n29635));
    NOR2X1 U16764 (.A1(N9294), .A2(N7913), .ZN(n29636));
    NANDX1 U16765 (.A1(N9668), .A2(n23979), .ZN(n29637));
    NANDX1 U16766 (.A1(N6405), .A2(N6980), .ZN(n29638));
    INVX1 U16767 (.I(n24931), .ZN(n29639));
    NOR2X1 U16768 (.A1(n24351), .A2(n18507), .ZN(N29640));
    NOR2X1 U16769 (.A1(n18861), .A2(n19049), .ZN(N29641));
    NANDX1 U16770 (.A1(N12245), .A2(n14550), .ZN(n29642));
    INVX1 U16771 (.I(n18246), .ZN(N29643));
    NOR2X1 U16772 (.A1(n22036), .A2(n19293), .ZN(n29644));
    NOR2X1 U16773 (.A1(N6761), .A2(N11195), .ZN(N29645));
    NOR2X1 U16774 (.A1(n18090), .A2(N4667), .ZN(N29646));
    NANDX1 U16775 (.A1(n16151), .A2(N12579), .ZN(n29647));
    NOR2X1 U16776 (.A1(N317), .A2(n25325), .ZN(N29648));
    NANDX1 U16777 (.A1(N6721), .A2(n21072), .ZN(N29649));
    INVX1 U16778 (.I(n20420), .ZN(n29650));
    NANDX1 U16779 (.A1(N2319), .A2(n13424), .ZN(N29651));
    NANDX1 U16780 (.A1(n21180), .A2(N6971), .ZN(N29652));
    INVX1 U16781 (.I(N7922), .ZN(n29653));
    INVX1 U16782 (.I(N3402), .ZN(N29654));
    NOR2X1 U16783 (.A1(n20954), .A2(n25438), .ZN(N29655));
    INVX1 U16784 (.I(N1531), .ZN(n29656));
    NANDX1 U16785 (.A1(N8688), .A2(N11042), .ZN(N29657));
    NOR2X1 U16786 (.A1(n13354), .A2(n21507), .ZN(N29658));
    INVX1 U16787 (.I(n14700), .ZN(N29659));
    NOR2X1 U16788 (.A1(n18788), .A2(N3290), .ZN(n29660));
    NOR2X1 U16789 (.A1(N7), .A2(n13130), .ZN(n29661));
    NOR2X1 U16790 (.A1(n20426), .A2(n21497), .ZN(N29662));
    NANDX1 U16791 (.A1(n22617), .A2(n14793), .ZN(N29663));
    NOR2X1 U16792 (.A1(n18355), .A2(n24610), .ZN(n29664));
    NOR2X1 U16793 (.A1(N3140), .A2(N2509), .ZN(n29665));
    NANDX1 U16794 (.A1(n24094), .A2(n16714), .ZN(N29666));
    INVX1 U16795 (.I(n14392), .ZN(n29667));
    NOR2X1 U16796 (.A1(N9125), .A2(n14201), .ZN(N29668));
    NOR2X1 U16797 (.A1(n22478), .A2(n24475), .ZN(N29669));
    INVX1 U16798 (.I(N443), .ZN(N29670));
    NOR2X1 U16799 (.A1(N754), .A2(n18002), .ZN(n29671));
    NANDX1 U16800 (.A1(N760), .A2(n19899), .ZN(n29672));
    INVX1 U16801 (.I(N9953), .ZN(n29673));
    NANDX1 U16802 (.A1(n18469), .A2(n21337), .ZN(n29674));
    NOR2X1 U16803 (.A1(N6753), .A2(n14190), .ZN(n29675));
    INVX1 U16804 (.I(n17227), .ZN(N29676));
    NANDX1 U16805 (.A1(n21069), .A2(n17134), .ZN(n29677));
    INVX1 U16806 (.I(N1049), .ZN(n29678));
    NANDX1 U16807 (.A1(N7847), .A2(n13226), .ZN(N29679));
    NANDX1 U16808 (.A1(n22048), .A2(N2222), .ZN(n29680));
    INVX1 U16809 (.I(n21020), .ZN(n29681));
    NANDX1 U16810 (.A1(N1648), .A2(n21810), .ZN(N29682));
    NOR2X1 U16811 (.A1(n19649), .A2(N9418), .ZN(n29683));
    NOR2X1 U16812 (.A1(N2814), .A2(n24048), .ZN(n29684));
    INVX1 U16813 (.I(n18706), .ZN(n29685));
    NANDX1 U16814 (.A1(n20026), .A2(N1425), .ZN(N29686));
    INVX1 U16815 (.I(n22983), .ZN(n29687));
    NANDX1 U16816 (.A1(n15491), .A2(N3577), .ZN(n29688));
    NANDX1 U16817 (.A1(n21392), .A2(n22535), .ZN(n29689));
    NANDX1 U16818 (.A1(n13460), .A2(N4879), .ZN(N29690));
    INVX1 U16819 (.I(N3420), .ZN(N29691));
    NOR2X1 U16820 (.A1(N9582), .A2(n15857), .ZN(n29692));
    NANDX1 U16821 (.A1(n19270), .A2(n17504), .ZN(N29693));
    INVX1 U16822 (.I(n18480), .ZN(n29694));
    INVX1 U16823 (.I(N5705), .ZN(n29695));
    NANDX1 U16824 (.A1(N3232), .A2(N4250), .ZN(n29696));
    NOR2X1 U16825 (.A1(N10705), .A2(N10032), .ZN(n29697));
    INVX1 U16826 (.I(N12130), .ZN(n29698));
    NANDX1 U16827 (.A1(N12178), .A2(n20882), .ZN(N29699));
    NANDX1 U16828 (.A1(n15754), .A2(n25201), .ZN(N29700));
    NANDX1 U16829 (.A1(N1554), .A2(n19336), .ZN(n29701));
    NOR2X1 U16830 (.A1(N6433), .A2(N12426), .ZN(n29702));
    NOR2X1 U16831 (.A1(N10894), .A2(N10775), .ZN(N29703));
    NOR2X1 U16832 (.A1(N10873), .A2(N4543), .ZN(n29704));
    INVX1 U16833 (.I(N7160), .ZN(n29705));
    INVX1 U16834 (.I(n25405), .ZN(n29706));
    INVX1 U16835 (.I(n19005), .ZN(n29707));
    NANDX1 U16836 (.A1(n20151), .A2(n13677), .ZN(n29708));
    NANDX1 U16837 (.A1(N4681), .A2(N2872), .ZN(n29709));
    INVX1 U16838 (.I(N1744), .ZN(n29710));
    INVX1 U16839 (.I(n24385), .ZN(N29711));
    NOR2X1 U16840 (.A1(n19571), .A2(N12852), .ZN(N29712));
    NANDX1 U16841 (.A1(n21124), .A2(N6685), .ZN(N29713));
    NANDX1 U16842 (.A1(n16324), .A2(N7879), .ZN(n29714));
    INVX1 U16843 (.I(N1716), .ZN(n29715));
    NOR2X1 U16844 (.A1(n21290), .A2(N12588), .ZN(n29716));
    NANDX1 U16845 (.A1(n20775), .A2(N8515), .ZN(n29717));
    NANDX1 U16846 (.A1(N9445), .A2(N10146), .ZN(n29718));
    NANDX1 U16847 (.A1(N1347), .A2(N4795), .ZN(n29719));
    INVX1 U16848 (.I(n18223), .ZN(n29720));
    INVX1 U16849 (.I(N107), .ZN(n29721));
    INVX1 U16850 (.I(n25488), .ZN(n29722));
    INVX1 U16851 (.I(N9376), .ZN(n29723));
    NOR2X1 U16852 (.A1(N12261), .A2(n22227), .ZN(N29724));
    INVX1 U16853 (.I(n22153), .ZN(n29725));
    NOR2X1 U16854 (.A1(n14277), .A2(n12974), .ZN(N29726));
    NANDX1 U16855 (.A1(n16851), .A2(N3457), .ZN(N29727));
    INVX1 U16856 (.I(N12639), .ZN(n29728));
    NANDX1 U16857 (.A1(N5169), .A2(N7911), .ZN(N29729));
    INVX1 U16858 (.I(N3418), .ZN(n29730));
    NANDX1 U16859 (.A1(N12241), .A2(n23710), .ZN(N29731));
    INVX1 U16860 (.I(N5803), .ZN(n29732));
    NANDX1 U16861 (.A1(N189), .A2(N4045), .ZN(n29733));
    NANDX1 U16862 (.A1(N10682), .A2(n18300), .ZN(N29734));
    NOR2X1 U16863 (.A1(N8826), .A2(n21351), .ZN(n29735));
    NOR2X1 U16864 (.A1(N5550), .A2(n24679), .ZN(n29736));
    NOR2X1 U16865 (.A1(n23229), .A2(n13453), .ZN(n29737));
    NANDX1 U16866 (.A1(n23284), .A2(N4802), .ZN(n29738));
    NOR2X1 U16867 (.A1(n16490), .A2(n17440), .ZN(n29739));
    INVX1 U16868 (.I(n21658), .ZN(n29740));
    NOR2X1 U16869 (.A1(N9254), .A2(n13843), .ZN(n29741));
    NANDX1 U16870 (.A1(N10262), .A2(N12051), .ZN(N29742));
    NOR2X1 U16871 (.A1(n16064), .A2(n18725), .ZN(n29743));
    INVX1 U16872 (.I(N8876), .ZN(n29744));
    INVX1 U16873 (.I(n16115), .ZN(n29745));
    NANDX1 U16874 (.A1(N2511), .A2(n24940), .ZN(N29746));
    NANDX1 U16875 (.A1(n14242), .A2(n19257), .ZN(N29747));
    INVX1 U16876 (.I(N11391), .ZN(N29748));
    NOR2X1 U16877 (.A1(N10151), .A2(N10282), .ZN(n29749));
    INVX1 U16878 (.I(N3720), .ZN(N29750));
    NANDX1 U16879 (.A1(n20022), .A2(N9927), .ZN(N29751));
    NOR2X1 U16880 (.A1(N4945), .A2(n24044), .ZN(n29752));
    NANDX1 U16881 (.A1(n18788), .A2(N7550), .ZN(n29753));
    INVX1 U16882 (.I(N5336), .ZN(n29754));
    INVX1 U16883 (.I(n21670), .ZN(n29755));
    INVX1 U16884 (.I(n15188), .ZN(n29756));
    INVX1 U16885 (.I(n15868), .ZN(n29757));
    NANDX1 U16886 (.A1(n20987), .A2(n18378), .ZN(n29758));
    INVX1 U16887 (.I(N7276), .ZN(n29759));
    NOR2X1 U16888 (.A1(n13262), .A2(N3974), .ZN(N29760));
    NOR2X1 U16889 (.A1(n19013), .A2(N2893), .ZN(n29761));
    NANDX1 U16890 (.A1(N11313), .A2(n20882), .ZN(n29762));
    INVX1 U16891 (.I(n20103), .ZN(n29763));
    NOR2X1 U16892 (.A1(N5044), .A2(n25047), .ZN(N29764));
    NANDX1 U16893 (.A1(N389), .A2(n18332), .ZN(N29765));
    INVX1 U16894 (.I(N5995), .ZN(n29766));
    NOR2X1 U16895 (.A1(n24190), .A2(n16432), .ZN(N29767));
    NOR2X1 U16896 (.A1(N2644), .A2(N10243), .ZN(N29768));
    INVX1 U16897 (.I(N8443), .ZN(n29769));
    NOR2X1 U16898 (.A1(n22773), .A2(N2448), .ZN(n29770));
    INVX1 U16899 (.I(n18658), .ZN(n29771));
    NOR2X1 U16900 (.A1(n20014), .A2(n14701), .ZN(n29772));
    INVX1 U16901 (.I(N11674), .ZN(n29773));
    NANDX1 U16902 (.A1(n23569), .A2(N7054), .ZN(n29774));
    NOR2X1 U16903 (.A1(n18169), .A2(N1128), .ZN(n29775));
    INVX1 U16904 (.I(n17714), .ZN(n29776));
    INVX1 U16905 (.I(N482), .ZN(n29777));
    NANDX1 U16906 (.A1(n22448), .A2(N6476), .ZN(n29778));
    NOR2X1 U16907 (.A1(N9903), .A2(N11675), .ZN(N29779));
    NANDX1 U16908 (.A1(N12546), .A2(N10686), .ZN(n29780));
    INVX1 U16909 (.I(N9757), .ZN(n29781));
    INVX1 U16910 (.I(N1938), .ZN(n29782));
    NANDX1 U16911 (.A1(n21220), .A2(n20595), .ZN(n29783));
    NANDX1 U16912 (.A1(N4500), .A2(n24063), .ZN(n29784));
    NOR2X1 U16913 (.A1(n16173), .A2(n22624), .ZN(N29785));
    NOR2X1 U16914 (.A1(N11994), .A2(N3404), .ZN(N29786));
    NANDX1 U16915 (.A1(n13121), .A2(N3497), .ZN(N29787));
    NOR2X1 U16916 (.A1(N9902), .A2(n18248), .ZN(n29788));
    NANDX1 U16917 (.A1(N6847), .A2(n13491), .ZN(N29789));
    INVX1 U16918 (.I(n16749), .ZN(n29790));
    NOR2X1 U16919 (.A1(N11976), .A2(n18063), .ZN(n29791));
    INVX1 U16920 (.I(n16643), .ZN(n29792));
    NANDX1 U16921 (.A1(N4296), .A2(n18580), .ZN(n29793));
    INVX1 U16922 (.I(n14283), .ZN(N29794));
    INVX1 U16923 (.I(N8735), .ZN(N29795));
    NOR2X1 U16924 (.A1(n15270), .A2(N936), .ZN(N29796));
    INVX1 U16925 (.I(N12392), .ZN(n29797));
    INVX1 U16926 (.I(N10214), .ZN(N29798));
    NANDX1 U16927 (.A1(n13909), .A2(N12103), .ZN(n29799));
    NANDX1 U16928 (.A1(N3324), .A2(n22004), .ZN(n29800));
    NOR2X1 U16929 (.A1(N3282), .A2(n17618), .ZN(n29801));
    NOR2X1 U16930 (.A1(N3752), .A2(n23134), .ZN(N29802));
    NANDX1 U16931 (.A1(N4495), .A2(n15694), .ZN(n29803));
    INVX1 U16932 (.I(n21137), .ZN(N29804));
    NOR2X1 U16933 (.A1(n20405), .A2(N2982), .ZN(n29805));
    INVX1 U16934 (.I(N9185), .ZN(n29806));
    INVX1 U16935 (.I(N7567), .ZN(n29807));
    NOR2X1 U16936 (.A1(N9459), .A2(N8502), .ZN(N29808));
    NOR2X1 U16937 (.A1(n21850), .A2(N2743), .ZN(n29809));
    NANDX1 U16938 (.A1(n15180), .A2(n16651), .ZN(n29810));
    INVX1 U16939 (.I(N12006), .ZN(N29811));
    NANDX1 U16940 (.A1(N11307), .A2(N1577), .ZN(N29812));
    NOR2X1 U16941 (.A1(N3422), .A2(n18908), .ZN(N29813));
    NANDX1 U16942 (.A1(N1054), .A2(N10399), .ZN(n29814));
    NANDX1 U16943 (.A1(N5515), .A2(N12238), .ZN(n29815));
    NOR2X1 U16944 (.A1(N12293), .A2(n21410), .ZN(N29816));
    NANDX1 U16945 (.A1(n22357), .A2(n19363), .ZN(N29817));
    NOR2X1 U16946 (.A1(N4422), .A2(N10595), .ZN(n29818));
    NANDX1 U16947 (.A1(N1691), .A2(n14317), .ZN(n29819));
    INVX1 U16948 (.I(N4433), .ZN(N29820));
    INVX1 U16949 (.I(n14632), .ZN(n29821));
    INVX1 U16950 (.I(n17556), .ZN(N29822));
    NANDX1 U16951 (.A1(N4324), .A2(n17630), .ZN(n29823));
    NOR2X1 U16952 (.A1(N5115), .A2(n21052), .ZN(n29824));
    NOR2X1 U16953 (.A1(N9657), .A2(N10873), .ZN(N29825));
    NOR2X1 U16954 (.A1(N7462), .A2(N5155), .ZN(n29826));
    NOR2X1 U16955 (.A1(N902), .A2(n17447), .ZN(n29827));
    INVX1 U16956 (.I(N11593), .ZN(n29828));
    NANDX1 U16957 (.A1(N326), .A2(N5240), .ZN(N29829));
    NOR2X1 U16958 (.A1(N10920), .A2(n19578), .ZN(n29830));
    NANDX1 U16959 (.A1(n25236), .A2(n19030), .ZN(n29831));
    NANDX1 U16960 (.A1(n16753), .A2(N8160), .ZN(n29832));
    NOR2X1 U16961 (.A1(N8806), .A2(n23564), .ZN(N29833));
    NANDX1 U16962 (.A1(N934), .A2(N3811), .ZN(n29834));
    NOR2X1 U16963 (.A1(N10753), .A2(N2964), .ZN(n29835));
    NOR2X1 U16964 (.A1(N10393), .A2(N12516), .ZN(N29836));
    NANDX1 U16965 (.A1(n15547), .A2(N8804), .ZN(N29837));
    INVX1 U16966 (.I(n21762), .ZN(n29838));
    INVX1 U16967 (.I(n20623), .ZN(n29839));
    INVX1 U16968 (.I(n15594), .ZN(N29840));
    NOR2X1 U16969 (.A1(n21089), .A2(n15281), .ZN(n29841));
    INVX1 U16970 (.I(n19037), .ZN(n29842));
    NANDX1 U16971 (.A1(N2233), .A2(N10186), .ZN(N29843));
    NOR2X1 U16972 (.A1(n24662), .A2(N11186), .ZN(n29844));
    NOR2X1 U16973 (.A1(n22723), .A2(N5277), .ZN(N29845));
    NANDX1 U16974 (.A1(n15301), .A2(n18752), .ZN(N29846));
    NANDX1 U16975 (.A1(n18265), .A2(n16382), .ZN(n29847));
    INVX1 U16976 (.I(N5278), .ZN(n29848));
    NANDX1 U16977 (.A1(N7765), .A2(N2849), .ZN(N29849));
    NOR2X1 U16978 (.A1(n18294), .A2(n18117), .ZN(N29850));
    NOR2X1 U16979 (.A1(n17622), .A2(n22478), .ZN(n29851));
    NANDX1 U16980 (.A1(n13208), .A2(N12256), .ZN(N29852));
    INVX1 U16981 (.I(n21013), .ZN(N29853));
    INVX1 U16982 (.I(N11417), .ZN(n29854));
    INVX1 U16983 (.I(N11069), .ZN(N29855));
    NANDX1 U16984 (.A1(N5650), .A2(N3674), .ZN(n29856));
    NOR2X1 U16985 (.A1(n25196), .A2(N11482), .ZN(N29857));
    NOR2X1 U16986 (.A1(n18446), .A2(N4540), .ZN(n29858));
    INVX1 U16987 (.I(N9325), .ZN(n29859));
    INVX1 U16988 (.I(n24174), .ZN(n29860));
    NOR2X1 U16989 (.A1(N4522), .A2(N1521), .ZN(n29861));
    NOR2X1 U16990 (.A1(n22816), .A2(N8405), .ZN(n29862));
    NANDX1 U16991 (.A1(N3703), .A2(n19651), .ZN(N29863));
    INVX1 U16992 (.I(N5679), .ZN(n29864));
    NOR2X1 U16993 (.A1(N652), .A2(N1189), .ZN(n29865));
    INVX1 U16994 (.I(N836), .ZN(N29866));
    INVX1 U16995 (.I(N11045), .ZN(n29867));
    INVX1 U16996 (.I(n15571), .ZN(n29868));
    NOR2X1 U16997 (.A1(N11013), .A2(n15265), .ZN(n29869));
    NANDX1 U16998 (.A1(N11645), .A2(N8208), .ZN(n29870));
    NANDX1 U16999 (.A1(N5039), .A2(N6300), .ZN(n29871));
    NOR2X1 U17000 (.A1(n17980), .A2(n14632), .ZN(n29872));
    NANDX1 U17001 (.A1(n19500), .A2(N2462), .ZN(N29873));
    INVX1 U17002 (.I(n16673), .ZN(N29874));
    NANDX1 U17003 (.A1(n24838), .A2(N10821), .ZN(N29875));
    NOR2X1 U17004 (.A1(N5014), .A2(N5992), .ZN(N29876));
    NANDX1 U17005 (.A1(N6202), .A2(N5968), .ZN(n29877));
    INVX1 U17006 (.I(N1853), .ZN(N29878));
    NOR2X1 U17007 (.A1(N12085), .A2(n17424), .ZN(N29879));
    NANDX1 U17008 (.A1(n23097), .A2(n21456), .ZN(n29880));
    INVX1 U17009 (.I(n23509), .ZN(n29881));
    INVX1 U17010 (.I(n21272), .ZN(n29882));
    NANDX1 U17011 (.A1(n13498), .A2(N800), .ZN(n29883));
    NOR2X1 U17012 (.A1(n16897), .A2(N10352), .ZN(n29884));
    INVX1 U17013 (.I(n19358), .ZN(N29885));
    NOR2X1 U17014 (.A1(N9230), .A2(N12807), .ZN(N29886));
    NANDX1 U17015 (.A1(N8818), .A2(N8955), .ZN(n29887));
    NOR2X1 U17016 (.A1(n14809), .A2(n20025), .ZN(n29888));
    INVX1 U17017 (.I(N9545), .ZN(n29889));
    INVX1 U17018 (.I(N7154), .ZN(n29890));
    INVX1 U17019 (.I(n18513), .ZN(n29891));
    NOR2X1 U17020 (.A1(n13357), .A2(N4875), .ZN(n29892));
    INVX1 U17021 (.I(n15123), .ZN(n29893));
    NANDX1 U17022 (.A1(n16496), .A2(N10893), .ZN(N29894));
    NOR2X1 U17023 (.A1(N4491), .A2(N11692), .ZN(n29895));
    NOR2X1 U17024 (.A1(n21387), .A2(N10811), .ZN(n29896));
    INVX1 U17025 (.I(N4010), .ZN(n29897));
    NANDX1 U17026 (.A1(N6270), .A2(N5584), .ZN(n29898));
    INVX1 U17027 (.I(n15087), .ZN(N29899));
    NOR2X1 U17028 (.A1(N9981), .A2(n18664), .ZN(n29900));
    NOR2X1 U17029 (.A1(n15281), .A2(n16976), .ZN(N29901));
    NOR2X1 U17030 (.A1(N11202), .A2(n21067), .ZN(n29902));
    NANDX1 U17031 (.A1(n13314), .A2(n23191), .ZN(n29903));
    NANDX1 U17032 (.A1(N11379), .A2(N12812), .ZN(n29904));
    INVX1 U17033 (.I(N2372), .ZN(n29905));
    NANDX1 U17034 (.A1(n25215), .A2(n21132), .ZN(n29906));
    NANDX1 U17035 (.A1(N4196), .A2(N5784), .ZN(N29907));
    INVX1 U17036 (.I(N1237), .ZN(n29908));
    NOR2X1 U17037 (.A1(N3802), .A2(N7506), .ZN(n29909));
    NOR2X1 U17038 (.A1(N3450), .A2(N11361), .ZN(n29910));
    INVX1 U17039 (.I(n13430), .ZN(n29911));
    NANDX1 U17040 (.A1(n16510), .A2(N3209), .ZN(n29912));
    INVX1 U17041 (.I(N9534), .ZN(N29913));
    INVX1 U17042 (.I(n17061), .ZN(n29914));
    NANDX1 U17043 (.A1(N2222), .A2(n14750), .ZN(n29915));
    INVX1 U17044 (.I(N2368), .ZN(n29916));
    INVX1 U17045 (.I(N5766), .ZN(n29917));
    INVX1 U17046 (.I(N3298), .ZN(N29918));
    INVX1 U17047 (.I(n14639), .ZN(n29919));
    NOR2X1 U17048 (.A1(N12711), .A2(n20423), .ZN(n29920));
    INVX1 U17049 (.I(n13947), .ZN(n29921));
    NANDX1 U17050 (.A1(N7036), .A2(N10221), .ZN(n29922));
    NOR2X1 U17051 (.A1(N10486), .A2(n21581), .ZN(N29923));
    INVX1 U17052 (.I(n23915), .ZN(n29924));
    NOR2X1 U17053 (.A1(N10351), .A2(n15891), .ZN(N29925));
    INVX1 U17054 (.I(n19884), .ZN(N29926));
    INVX1 U17055 (.I(N5460), .ZN(N29927));
    INVX1 U17056 (.I(n21290), .ZN(N29928));
    INVX1 U17057 (.I(N1926), .ZN(n29929));
    NANDX1 U17058 (.A1(n25305), .A2(n21961), .ZN(n29930));
    NOR2X1 U17059 (.A1(n17370), .A2(n16206), .ZN(N29931));
    INVX1 U17060 (.I(N8096), .ZN(n29932));
    NANDX1 U17061 (.A1(n15491), .A2(N11330), .ZN(n29933));
    INVX1 U17062 (.I(N8971), .ZN(N29934));
    INVX1 U17063 (.I(n16349), .ZN(N29935));
    NOR2X1 U17064 (.A1(N6387), .A2(N1195), .ZN(n29936));
    INVX1 U17065 (.I(N4799), .ZN(n29937));
    NANDX1 U17066 (.A1(N10786), .A2(N9458), .ZN(n29938));
    NOR2X1 U17067 (.A1(N5167), .A2(n14256), .ZN(n29939));
    NOR2X1 U17068 (.A1(N9385), .A2(n24313), .ZN(n29940));
    INVX1 U17069 (.I(N78), .ZN(n29941));
    NANDX1 U17070 (.A1(N7469), .A2(n22038), .ZN(N29942));
    NANDX1 U17071 (.A1(n24839), .A2(N12741), .ZN(n29943));
    NOR2X1 U17072 (.A1(n21702), .A2(n16155), .ZN(N29944));
    NANDX1 U17073 (.A1(n21799), .A2(n22283), .ZN(n29945));
    NANDX1 U17074 (.A1(n17700), .A2(n13129), .ZN(N29946));
    NOR2X1 U17075 (.A1(n24086), .A2(n14323), .ZN(N29947));
    NOR2X1 U17076 (.A1(n17653), .A2(n19154), .ZN(N29948));
    NANDX1 U17077 (.A1(N1608), .A2(n23616), .ZN(n29949));
    INVX1 U17078 (.I(n15863), .ZN(n29950));
    NANDX1 U17079 (.A1(N6826), .A2(n14673), .ZN(n29951));
    NOR2X1 U17080 (.A1(N6903), .A2(N405), .ZN(N29952));
    NANDX1 U17081 (.A1(N3439), .A2(n14533), .ZN(N29953));
    INVX1 U17082 (.I(n16179), .ZN(n29954));
    NANDX1 U17083 (.A1(N10511), .A2(n21101), .ZN(N29955));
    NOR2X1 U17084 (.A1(N6807), .A2(n17881), .ZN(N29956));
    NOR2X1 U17085 (.A1(n24507), .A2(n19777), .ZN(N29957));
    NOR2X1 U17086 (.A1(N11858), .A2(n22867), .ZN(n29958));
    NOR2X1 U17087 (.A1(N4008), .A2(N5286), .ZN(N29959));
    INVX1 U17088 (.I(N5615), .ZN(N29960));
    NOR2X1 U17089 (.A1(n20058), .A2(N10245), .ZN(n29961));
    NANDX1 U17090 (.A1(N1381), .A2(n13685), .ZN(n29962));
    NANDX1 U17091 (.A1(n22553), .A2(n14090), .ZN(n29963));
    NOR2X1 U17092 (.A1(N489), .A2(n17390), .ZN(n29964));
    INVX1 U17093 (.I(N5436), .ZN(N29965));
    INVX1 U17094 (.I(n18964), .ZN(N29966));
    NOR2X1 U17095 (.A1(N4833), .A2(n14539), .ZN(n29967));
    NANDX1 U17096 (.A1(n13436), .A2(N2311), .ZN(n29968));
    NANDX1 U17097 (.A1(n14324), .A2(n14168), .ZN(N29969));
    NOR2X1 U17098 (.A1(n22203), .A2(n18176), .ZN(n29970));
    INVX1 U17099 (.I(n19317), .ZN(n29971));
    NANDX1 U17100 (.A1(n14082), .A2(N2640), .ZN(N29972));
    NANDX1 U17101 (.A1(n17321), .A2(N4020), .ZN(n29973));
    NOR2X1 U17102 (.A1(n25028), .A2(n15341), .ZN(n29974));
    NANDX1 U17103 (.A1(N7939), .A2(n15829), .ZN(N29975));
    NANDX1 U17104 (.A1(n16392), .A2(N10032), .ZN(N29976));
    NANDX1 U17105 (.A1(n24124), .A2(n25336), .ZN(n29977));
    NANDX1 U17106 (.A1(N1928), .A2(N10554), .ZN(n29978));
    NOR2X1 U17107 (.A1(n18508), .A2(n15548), .ZN(n29979));
    NANDX1 U17108 (.A1(N7173), .A2(n17907), .ZN(N29980));
    INVX1 U17109 (.I(n14116), .ZN(N29981));
    INVX1 U17110 (.I(n25026), .ZN(n29982));
    NOR2X1 U17111 (.A1(N5937), .A2(N2163), .ZN(n29983));
    INVX1 U17112 (.I(n23257), .ZN(N29984));
    NOR2X1 U17113 (.A1(n23726), .A2(N11550), .ZN(n29985));
    INVX1 U17114 (.I(N12066), .ZN(n29986));
    NOR2X1 U17115 (.A1(n14887), .A2(N6563), .ZN(N29987));
    NOR2X1 U17116 (.A1(n13687), .A2(n16676), .ZN(N29988));
    NOR2X1 U17117 (.A1(N2288), .A2(n20389), .ZN(n29989));
    INVX1 U17118 (.I(N12841), .ZN(n29990));
    NANDX1 U17119 (.A1(N6969), .A2(N2886), .ZN(n29991));
    INVX1 U17120 (.I(N2909), .ZN(n29992));
    NOR2X1 U17121 (.A1(N1251), .A2(N5793), .ZN(n29993));
    NOR2X1 U17122 (.A1(N774), .A2(n21234), .ZN(n29994));
    INVX1 U17123 (.I(n17207), .ZN(n29995));
    INVX1 U17124 (.I(N5106), .ZN(n29996));
    INVX1 U17125 (.I(n20966), .ZN(n29997));
    NOR2X1 U17126 (.A1(N11215), .A2(n21799), .ZN(n29998));
    INVX1 U17127 (.I(N599), .ZN(n29999));
    NANDX1 U17128 (.A1(n24056), .A2(n14285), .ZN(n30000));
    NANDX1 U17129 (.A1(N10590), .A2(N5340), .ZN(n30001));
    NANDX1 U17130 (.A1(n13321), .A2(n18180), .ZN(n30002));
    NOR2X1 U17131 (.A1(N9057), .A2(N9834), .ZN(n30003));
    NOR2X1 U17132 (.A1(N11965), .A2(n19394), .ZN(n30004));
    NANDX1 U17133 (.A1(n17757), .A2(n20809), .ZN(n30005));
    NANDX1 U17134 (.A1(N2256), .A2(N2658), .ZN(n30006));
    NOR2X1 U17135 (.A1(N10728), .A2(N7763), .ZN(N30007));
    INVX1 U17136 (.I(n20462), .ZN(N30008));
    INVX1 U17137 (.I(N8438), .ZN(N30009));
    INVX1 U17138 (.I(N12593), .ZN(n30010));
    NOR2X1 U17139 (.A1(n22655), .A2(n25416), .ZN(n30011));
    NANDX1 U17140 (.A1(N5454), .A2(N10503), .ZN(N30012));
    INVX1 U17141 (.I(n22912), .ZN(n30013));
    NANDX1 U17142 (.A1(n24376), .A2(n15672), .ZN(n30014));
    NOR2X1 U17143 (.A1(N8707), .A2(n18243), .ZN(N30015));
    NOR2X1 U17144 (.A1(n16868), .A2(n22065), .ZN(n30016));
    NOR2X1 U17145 (.A1(N12174), .A2(N1159), .ZN(n30017));
    INVX1 U17146 (.I(N3599), .ZN(n30018));
    INVX1 U17147 (.I(N5153), .ZN(n30019));
    INVX1 U17148 (.I(N8952), .ZN(n30020));
    NANDX1 U17149 (.A1(n13314), .A2(n17389), .ZN(n30021));
    NOR2X1 U17150 (.A1(N404), .A2(N3961), .ZN(n30022));
    NOR2X1 U17151 (.A1(N318), .A2(N4818), .ZN(n30023));
    NANDX1 U17152 (.A1(n25090), .A2(N11014), .ZN(n30024));
    NANDX1 U17153 (.A1(N947), .A2(N9887), .ZN(n30025));
    NANDX1 U17154 (.A1(n22593), .A2(N7362), .ZN(n30026));
    NANDX1 U17155 (.A1(N8238), .A2(n24229), .ZN(N30027));
    INVX1 U17156 (.I(N11640), .ZN(n30028));
    NOR2X1 U17157 (.A1(N6629), .A2(n17297), .ZN(n30029));
    NOR2X1 U17158 (.A1(n18356), .A2(N11217), .ZN(n30030));
    NANDX1 U17159 (.A1(n16075), .A2(N97), .ZN(N30031));
    INVX1 U17160 (.I(n22232), .ZN(n30032));
    NANDX1 U17161 (.A1(N5880), .A2(N690), .ZN(n30033));
    NANDX1 U17162 (.A1(n20467), .A2(N5507), .ZN(N30034));
    INVX1 U17163 (.I(N8823), .ZN(N30035));
    NOR2X1 U17164 (.A1(N9067), .A2(N9769), .ZN(N30036));
    INVX1 U17165 (.I(N10964), .ZN(n30037));
    NOR2X1 U17166 (.A1(n22536), .A2(N5602), .ZN(n30038));
    NOR2X1 U17167 (.A1(N10030), .A2(n22304), .ZN(n30039));
    INVX1 U17168 (.I(N9698), .ZN(n30040));
    INVX1 U17169 (.I(n21568), .ZN(n30041));
    NOR2X1 U17170 (.A1(N10553), .A2(N7282), .ZN(N30042));
    NANDX1 U17171 (.A1(N1126), .A2(N7378), .ZN(n30043));
    NOR2X1 U17172 (.A1(n23357), .A2(n16149), .ZN(N30044));
    NOR2X1 U17173 (.A1(n24046), .A2(N5245), .ZN(N30045));
    NOR2X1 U17174 (.A1(N4051), .A2(N5622), .ZN(N30046));
    NANDX1 U17175 (.A1(n20570), .A2(N3456), .ZN(n30047));
    NOR2X1 U17176 (.A1(N10242), .A2(n14420), .ZN(n30048));
    NOR2X1 U17177 (.A1(n21545), .A2(N8789), .ZN(n30049));
    NANDX1 U17178 (.A1(N6073), .A2(n19860), .ZN(N30050));
    NOR2X1 U17179 (.A1(N4538), .A2(N12057), .ZN(n30051));
    NANDX1 U17180 (.A1(n20540), .A2(n22609), .ZN(n30052));
    NANDX1 U17181 (.A1(n14435), .A2(N12502), .ZN(n30053));
    INVX1 U17182 (.I(N2574), .ZN(n30054));
    NOR2X1 U17183 (.A1(n15744), .A2(n22095), .ZN(n30055));
    NOR2X1 U17184 (.A1(n20988), .A2(N11078), .ZN(n30056));
    NOR2X1 U17185 (.A1(n15377), .A2(N8883), .ZN(N30057));
    NOR2X1 U17186 (.A1(n18833), .A2(n16456), .ZN(n30058));
    INVX1 U17187 (.I(n22020), .ZN(N30059));
    NANDX1 U17188 (.A1(N6107), .A2(n19576), .ZN(N30060));
    INVX1 U17189 (.I(N947), .ZN(n30061));
    NANDX1 U17190 (.A1(N1319), .A2(n19755), .ZN(n30062));
    NOR2X1 U17191 (.A1(n22989), .A2(n14792), .ZN(n30063));
    NOR2X1 U17192 (.A1(N936), .A2(n17995), .ZN(N30064));
    NANDX1 U17193 (.A1(N11762), .A2(N9336), .ZN(n30065));
    NANDX1 U17194 (.A1(n16273), .A2(N5928), .ZN(N30066));
    INVX1 U17195 (.I(N11759), .ZN(n30067));
    NANDX1 U17196 (.A1(n22872), .A2(n15903), .ZN(n30068));
    NANDX1 U17197 (.A1(N8425), .A2(n23503), .ZN(n30069));
    INVX1 U17198 (.I(N7257), .ZN(N30070));
    INVX1 U17199 (.I(N2799), .ZN(n30071));
    INVX1 U17200 (.I(n14093), .ZN(n30072));
    INVX1 U17201 (.I(N3078), .ZN(n30073));
    INVX1 U17202 (.I(n22641), .ZN(n30074));
    NANDX1 U17203 (.A1(n17279), .A2(n20127), .ZN(n30075));
    NANDX1 U17204 (.A1(N3640), .A2(n21062), .ZN(n30076));
    INVX1 U17205 (.I(N2502), .ZN(N30077));
    INVX1 U17206 (.I(n16987), .ZN(n30078));
    INVX1 U17207 (.I(N12362), .ZN(N30079));
    INVX1 U17208 (.I(N7372), .ZN(N30080));
    NOR2X1 U17209 (.A1(N3185), .A2(N4741), .ZN(n30081));
    INVX1 U17210 (.I(n17839), .ZN(n30082));
    INVX1 U17211 (.I(N1289), .ZN(n30083));
    NANDX1 U17212 (.A1(N9189), .A2(N10077), .ZN(N30084));
    NANDX1 U17213 (.A1(N11320), .A2(n12937), .ZN(N30085));
    NANDX1 U17214 (.A1(N3165), .A2(N4228), .ZN(n30086));
    NANDX1 U17215 (.A1(N3532), .A2(n21506), .ZN(n30087));
    NOR2X1 U17216 (.A1(n18690), .A2(n25145), .ZN(n30088));
    INVX1 U17217 (.I(n15109), .ZN(n30089));
    NANDX1 U17218 (.A1(n22784), .A2(N6593), .ZN(n30090));
    INVX1 U17219 (.I(n23914), .ZN(N30091));
    INVX1 U17220 (.I(n24272), .ZN(n30092));
    NOR2X1 U17221 (.A1(N10226), .A2(n17780), .ZN(N30093));
    NOR2X1 U17222 (.A1(n16833), .A2(n19713), .ZN(n30094));
    NANDX1 U17223 (.A1(n17815), .A2(n17669), .ZN(n30095));
    INVX1 U17224 (.I(n21595), .ZN(N30096));
    NOR2X1 U17225 (.A1(n16424), .A2(n21195), .ZN(N30097));
    NANDX1 U17226 (.A1(n20651), .A2(N3663), .ZN(N30098));
    NANDX1 U17227 (.A1(n16655), .A2(N9296), .ZN(n30099));
    INVX1 U17228 (.I(N5065), .ZN(n30100));
    NOR2X1 U17229 (.A1(n21515), .A2(n21479), .ZN(n30101));
    INVX1 U17230 (.I(n16875), .ZN(N30102));
    NANDX1 U17231 (.A1(n20451), .A2(n23916), .ZN(n30103));
    NANDX1 U17232 (.A1(N6248), .A2(n22910), .ZN(N30104));
    INVX1 U17233 (.I(N9602), .ZN(N30105));
    NOR2X1 U17234 (.A1(N1171), .A2(N3013), .ZN(n30106));
    INVX1 U17235 (.I(N7608), .ZN(n30107));
    INVX1 U17236 (.I(n16914), .ZN(N30108));
    NANDX1 U17237 (.A1(n22924), .A2(N12606), .ZN(N30109));
    NANDX1 U17238 (.A1(n18072), .A2(N5036), .ZN(N30110));
    INVX1 U17239 (.I(N9224), .ZN(N30111));
    INVX1 U17240 (.I(N6709), .ZN(n30112));
    NOR2X1 U17241 (.A1(n13588), .A2(n16991), .ZN(n30113));
    INVX1 U17242 (.I(N10125), .ZN(n30114));
    NOR2X1 U17243 (.A1(N677), .A2(n19344), .ZN(n30115));
    INVX1 U17244 (.I(N1090), .ZN(N30116));
    NANDX1 U17245 (.A1(N7222), .A2(N8050), .ZN(n30117));
    NOR2X1 U17246 (.A1(N10229), .A2(N9221), .ZN(N30118));
    NOR2X1 U17247 (.A1(N5548), .A2(N5596), .ZN(N30119));
    INVX1 U17248 (.I(n22461), .ZN(n30120));
    NOR2X1 U17249 (.A1(n19661), .A2(n23834), .ZN(n30121));
    INVX1 U17250 (.I(N12231), .ZN(n30122));
    INVX1 U17251 (.I(n18345), .ZN(N30123));
    NANDX1 U17252 (.A1(n20736), .A2(n13821), .ZN(N30124));
    INVX1 U17253 (.I(N8821), .ZN(n30125));
    NANDX1 U17254 (.A1(N1078), .A2(N7714), .ZN(n30126));
    INVX1 U17255 (.I(n16024), .ZN(N30127));
    NOR2X1 U17256 (.A1(N12254), .A2(N5881), .ZN(n30128));
    NANDX1 U17257 (.A1(n19475), .A2(n13931), .ZN(n30129));
    INVX1 U17258 (.I(n18471), .ZN(n30130));
    NOR2X1 U17259 (.A1(n18878), .A2(n24018), .ZN(n30131));
    INVX1 U17260 (.I(n15616), .ZN(n30132));
    INVX1 U17261 (.I(N505), .ZN(n30133));
    NANDX1 U17262 (.A1(N8075), .A2(n18547), .ZN(n30134));
    NANDX1 U17263 (.A1(N210), .A2(N157), .ZN(N30135));
    NANDX1 U17264 (.A1(N9713), .A2(n13977), .ZN(n30136));
    NOR2X1 U17265 (.A1(n18534), .A2(N8054), .ZN(N30137));
    NOR2X1 U17266 (.A1(n25676), .A2(N9614), .ZN(N30138));
    NOR2X1 U17267 (.A1(n14238), .A2(N4989), .ZN(N30139));
    INVX1 U17268 (.I(n21442), .ZN(N30140));
    INVX1 U17269 (.I(n15314), .ZN(N30141));
    NOR2X1 U17270 (.A1(n19387), .A2(n27086), .ZN(N30142));
    INVX1 U17271 (.I(N3636), .ZN(N30143));
    INVX1 U17272 (.I(n16711), .ZN(N30144));
    NOR2X1 U17273 (.A1(n29372), .A2(N6377), .ZN(n30145));
    INVX1 U17274 (.I(n21628), .ZN(N30146));
    NANDX1 U17275 (.A1(N3583), .A2(N2819), .ZN(n30147));
    NOR2X1 U17276 (.A1(N2107), .A2(n16885), .ZN(N30148));
    NANDX1 U17277 (.A1(n23393), .A2(n21190), .ZN(N30149));
    NANDX1 U17278 (.A1(n18931), .A2(N667), .ZN(N30150));
    INVX1 U17279 (.I(n21730), .ZN(n30151));
    NOR2X1 U17280 (.A1(n13193), .A2(N1595), .ZN(n30152));
    NOR2X1 U17281 (.A1(n17068), .A2(n28063), .ZN(n30153));
    NOR2X1 U17282 (.A1(n14016), .A2(N6495), .ZN(n30154));
    NOR2X1 U17283 (.A1(n27093), .A2(n23206), .ZN(N30155));
    NOR2X1 U17284 (.A1(n26327), .A2(n18143), .ZN(n30156));
    INVX1 U17285 (.I(N6378), .ZN(N30157));
    NOR2X1 U17286 (.A1(N11418), .A2(N9196), .ZN(N30158));
    NANDX1 U17287 (.A1(N2085), .A2(n14642), .ZN(n30159));
    NANDX1 U17288 (.A1(n25478), .A2(N5694), .ZN(n30160));
    NOR2X1 U17289 (.A1(N2832), .A2(n25058), .ZN(N30161));
    NANDX1 U17290 (.A1(n24561), .A2(N7834), .ZN(N30162));
    NOR2X1 U17291 (.A1(n14716), .A2(n23249), .ZN(N30163));
    NANDX1 U17292 (.A1(N12642), .A2(n27913), .ZN(N30164));
    INVX1 U17293 (.I(n19136), .ZN(N30165));
    INVX1 U17294 (.I(n26694), .ZN(n30166));
    NANDX1 U17295 (.A1(N7430), .A2(N11445), .ZN(n30167));
    NANDX1 U17296 (.A1(n15265), .A2(n17822), .ZN(n30168));
    INVX1 U17297 (.I(n26682), .ZN(N30169));
    NOR2X1 U17298 (.A1(N996), .A2(n28767), .ZN(N30170));
    NOR2X1 U17299 (.A1(N8056), .A2(N12668), .ZN(N30171));
    NANDX1 U17300 (.A1(n20678), .A2(n15499), .ZN(n30172));
    NOR2X1 U17301 (.A1(n17581), .A2(N9923), .ZN(n30173));
    NANDX1 U17302 (.A1(n27677), .A2(n13199), .ZN(N30174));
    INVX1 U17303 (.I(n24702), .ZN(n30175));
    NANDX1 U17304 (.A1(n25374), .A2(N12865), .ZN(N30176));
    NANDX1 U17305 (.A1(N8571), .A2(N9421), .ZN(N30177));
    NOR2X1 U17306 (.A1(N4561), .A2(n20865), .ZN(N30178));
    NOR2X1 U17307 (.A1(n19825), .A2(N8550), .ZN(N30179));
    INVX1 U17308 (.I(n16369), .ZN(N30180));
    NOR2X1 U17309 (.A1(n24183), .A2(N3559), .ZN(N30181));
    NOR2X1 U17310 (.A1(N2101), .A2(n16226), .ZN(n30182));
    INVX1 U17311 (.I(N11340), .ZN(N30183));
    NANDX1 U17312 (.A1(n15062), .A2(n28920), .ZN(N30184));
    NANDX1 U17313 (.A1(n19412), .A2(n26459), .ZN(n30185));
    NOR2X1 U17314 (.A1(n16873), .A2(N9585), .ZN(N30186));
    NOR2X1 U17315 (.A1(N12109), .A2(N11010), .ZN(N30187));
    INVX1 U17316 (.I(N9240), .ZN(N30188));
    INVX1 U17317 (.I(n23793), .ZN(N30189));
    INVX1 U17318 (.I(n29856), .ZN(N30190));
    INVX1 U17319 (.I(N3487), .ZN(N30191));
    NOR2X1 U17320 (.A1(n17036), .A2(N8417), .ZN(N30192));
    NOR2X1 U17321 (.A1(N11081), .A2(N11975), .ZN(N30193));
    NANDX1 U17322 (.A1(N1743), .A2(n16762), .ZN(N30194));
    NOR2X1 U17323 (.A1(n13082), .A2(N6910), .ZN(N30195));
    INVX1 U17324 (.I(N11864), .ZN(N30196));
    NANDX1 U17325 (.A1(n22290), .A2(n26884), .ZN(N30197));
    NANDX1 U17326 (.A1(N9025), .A2(n25029), .ZN(N30198));
    NANDX1 U17327 (.A1(N9694), .A2(N5901), .ZN(N30199));
    NOR2X1 U17328 (.A1(n18934), .A2(n14891), .ZN(n30200));
    NANDX1 U17329 (.A1(N2596), .A2(n14609), .ZN(N30201));
    NANDX1 U17330 (.A1(n24781), .A2(N11437), .ZN(n30202));
    NANDX1 U17331 (.A1(N3060), .A2(N2255), .ZN(N30203));
    NOR2X1 U17332 (.A1(N3595), .A2(n24541), .ZN(n30204));
    NANDX1 U17333 (.A1(n20356), .A2(n23797), .ZN(N30205));
    NANDX1 U17334 (.A1(n27265), .A2(n26675), .ZN(N30206));
    INVX1 U17335 (.I(n22805), .ZN(n30207));
    NOR2X1 U17336 (.A1(N7826), .A2(n20175), .ZN(N30208));
    NOR2X1 U17337 (.A1(n21415), .A2(N3637), .ZN(n30209));
    INVX1 U17338 (.I(n15876), .ZN(N30210));
    NANDX1 U17339 (.A1(n22160), .A2(N630), .ZN(n30211));
    NOR2X1 U17340 (.A1(n13317), .A2(N3799), .ZN(N30212));
    NANDX1 U17341 (.A1(n26658), .A2(n15236), .ZN(N30213));
    INVX1 U17342 (.I(n29717), .ZN(N30214));
    INVX1 U17343 (.I(n16230), .ZN(N30215));
    NANDX1 U17344 (.A1(N455), .A2(n13804), .ZN(N30216));
    INVX1 U17345 (.I(n24251), .ZN(N30217));
    INVX1 U17346 (.I(n27916), .ZN(N30218));
    INVX1 U17347 (.I(N5401), .ZN(N30219));
    NANDX1 U17348 (.A1(N5297), .A2(N1788), .ZN(n30220));
    NANDX1 U17349 (.A1(N10269), .A2(N11763), .ZN(N30221));
    NOR2X1 U17350 (.A1(n13495), .A2(n27639), .ZN(N30222));
    NANDX1 U17351 (.A1(n24216), .A2(n16829), .ZN(N30223));
    INVX1 U17352 (.I(n26093), .ZN(N30224));
    NANDX1 U17353 (.A1(N7091), .A2(n22613), .ZN(N30225));
    NANDX1 U17354 (.A1(n16049), .A2(n22192), .ZN(N30226));
    INVX1 U17355 (.I(n20839), .ZN(N30227));
    NANDX1 U17356 (.A1(N12230), .A2(n23203), .ZN(N30228));
    NOR2X1 U17357 (.A1(n25041), .A2(n17524), .ZN(n30229));
    NANDX1 U17358 (.A1(n22950), .A2(N11485), .ZN(N30230));
    INVX1 U17359 (.I(n28246), .ZN(n30231));
    NANDX1 U17360 (.A1(N9242), .A2(N8377), .ZN(n30232));
    NANDX1 U17361 (.A1(N12059), .A2(N10432), .ZN(N30233));
    NANDX1 U17362 (.A1(n21605), .A2(N4510), .ZN(n30234));
    NANDX1 U17363 (.A1(N4488), .A2(N465), .ZN(n30235));
    INVX1 U17364 (.I(N139), .ZN(N30236));
    NOR2X1 U17365 (.A1(N1261), .A2(N4748), .ZN(N30237));
    NOR2X1 U17366 (.A1(n13036), .A2(n25586), .ZN(n30238));
    NOR2X1 U17367 (.A1(n13826), .A2(n18651), .ZN(N30239));
    NANDX1 U17368 (.A1(n27427), .A2(n24735), .ZN(n30240));
    NOR2X1 U17369 (.A1(n20239), .A2(n24781), .ZN(N30241));
    INVX1 U17370 (.I(n18347), .ZN(N30242));
    INVX1 U17371 (.I(n22274), .ZN(N30243));
    NOR2X1 U17372 (.A1(N10071), .A2(N4196), .ZN(n30244));
    INVX1 U17373 (.I(N9728), .ZN(N30245));
    NOR2X1 U17374 (.A1(n18786), .A2(n26213), .ZN(n30246));
    NANDX1 U17375 (.A1(N7811), .A2(N3051), .ZN(N30247));
    NOR2X1 U17376 (.A1(n19449), .A2(N4311), .ZN(N30248));
    INVX1 U17377 (.I(N11701), .ZN(N30249));
    NANDX1 U17378 (.A1(n15003), .A2(n17879), .ZN(n30250));
    INVX1 U17379 (.I(N3516), .ZN(n30251));
    NANDX1 U17380 (.A1(n17021), .A2(n16812), .ZN(N30252));
    NANDX1 U17381 (.A1(n25820), .A2(N11455), .ZN(N30253));
    NOR2X1 U17382 (.A1(N2590), .A2(N7930), .ZN(n30254));
    NANDX1 U17383 (.A1(N6434), .A2(n18001), .ZN(N30255));
    INVX1 U17384 (.I(n20709), .ZN(N30256));
    NANDX1 U17385 (.A1(N876), .A2(n28055), .ZN(n30257));
    NANDX1 U17386 (.A1(n26983), .A2(n24427), .ZN(N30258));
    NANDX1 U17387 (.A1(n23091), .A2(n13738), .ZN(N30259));
    NANDX1 U17388 (.A1(N12507), .A2(n25438), .ZN(N30260));
    NOR2X1 U17389 (.A1(n27509), .A2(N1741), .ZN(n30261));
    INVX1 U17390 (.I(n19586), .ZN(N30262));
    NOR2X1 U17391 (.A1(N9367), .A2(N6260), .ZN(N30263));
    NANDX1 U17392 (.A1(N5049), .A2(n17714), .ZN(N30264));
    NANDX1 U17393 (.A1(N7638), .A2(n14204), .ZN(N30265));
    NANDX1 U17394 (.A1(n14071), .A2(n20765), .ZN(N30266));
    NANDX1 U17395 (.A1(n23340), .A2(N6917), .ZN(N30267));
    INVX1 U17396 (.I(n21258), .ZN(N30268));
    NOR2X1 U17397 (.A1(N8583), .A2(n15547), .ZN(n30269));
    NANDX1 U17398 (.A1(n20234), .A2(n17845), .ZN(N30270));
    NOR2X1 U17399 (.A1(n21301), .A2(n13145), .ZN(n30271));
    NOR2X1 U17400 (.A1(N7234), .A2(n14885), .ZN(N30272));
    INVX1 U17401 (.I(n15380), .ZN(N30273));
    NOR2X1 U17402 (.A1(n28746), .A2(n21639), .ZN(n30274));
    NOR2X1 U17403 (.A1(n22355), .A2(n27913), .ZN(N30275));
    INVX1 U17404 (.I(n18553), .ZN(n30276));
    NOR2X1 U17405 (.A1(n25865), .A2(N2486), .ZN(n30277));
    NOR2X1 U17406 (.A1(N6590), .A2(n14386), .ZN(N30278));
    NANDX1 U17407 (.A1(n18327), .A2(n24204), .ZN(N30279));
    INVX1 U17408 (.I(n15470), .ZN(N30280));
    NANDX1 U17409 (.A1(n29180), .A2(n24264), .ZN(N30281));
    NOR2X1 U17410 (.A1(N446), .A2(N3988), .ZN(n30282));
    NOR2X1 U17411 (.A1(n16040), .A2(n29919), .ZN(N30283));
    NOR2X1 U17412 (.A1(N5282), .A2(n15161), .ZN(N30284));
    INVX1 U17413 (.I(n22588), .ZN(n30285));
    NOR2X1 U17414 (.A1(n24481), .A2(n14805), .ZN(N30286));
    INVX1 U17415 (.I(n25999), .ZN(n30287));
    NANDX1 U17416 (.A1(N12236), .A2(N10288), .ZN(N30288));
    NANDX1 U17417 (.A1(n22101), .A2(n16877), .ZN(n30289));
    NANDX1 U17418 (.A1(N8745), .A2(n23764), .ZN(n30290));
    INVX1 U17419 (.I(n14669), .ZN(n30291));
    INVX1 U17420 (.I(N891), .ZN(N30292));
    INVX1 U17421 (.I(N10481), .ZN(N30293));
    INVX1 U17422 (.I(N2717), .ZN(n30294));
    NANDX1 U17423 (.A1(N4495), .A2(N7317), .ZN(N30295));
    NANDX1 U17424 (.A1(n25663), .A2(N12598), .ZN(N30296));
    NOR2X1 U17425 (.A1(N239), .A2(N5048), .ZN(N30297));
    NOR2X1 U17426 (.A1(n24719), .A2(N8413), .ZN(N30298));
    INVX1 U17427 (.I(N9142), .ZN(n30299));
    NANDX1 U17428 (.A1(n25685), .A2(n19429), .ZN(n30300));
    NOR2X1 U17429 (.A1(n17648), .A2(n24866), .ZN(N30301));
    NANDX1 U17430 (.A1(n26392), .A2(N7053), .ZN(n30302));
    NOR2X1 U17431 (.A1(n29621), .A2(n23407), .ZN(N30303));
    NOR2X1 U17432 (.A1(n20453), .A2(N3750), .ZN(n30304));
    NOR2X1 U17433 (.A1(N11730), .A2(n25476), .ZN(N30305));
    INVX1 U17434 (.I(n19046), .ZN(n30306));
    NANDX1 U17435 (.A1(N765), .A2(n20204), .ZN(N30307));
    NOR2X1 U17436 (.A1(n19702), .A2(n25251), .ZN(n30308));
    NOR2X1 U17437 (.A1(N2844), .A2(n22224), .ZN(N30309));
    NOR2X1 U17438 (.A1(N11985), .A2(N3718), .ZN(n30310));
    INVX1 U17439 (.I(n19974), .ZN(n30311));
    NANDX1 U17440 (.A1(n21640), .A2(N3263), .ZN(n30312));
    INVX1 U17441 (.I(N6456), .ZN(N30313));
    INVX1 U17442 (.I(n14366), .ZN(N30314));
    NANDX1 U17443 (.A1(N3584), .A2(N9642), .ZN(n30315));
    NANDX1 U17444 (.A1(n26031), .A2(N10387), .ZN(N30316));
    NANDX1 U17445 (.A1(n21370), .A2(n15626), .ZN(N30317));
    NOR2X1 U17446 (.A1(N8079), .A2(N4952), .ZN(n30318));
    NANDX1 U17447 (.A1(N12759), .A2(n24653), .ZN(N30319));
    NOR2X1 U17448 (.A1(n19193), .A2(n27496), .ZN(n30320));
    NOR2X1 U17449 (.A1(n27638), .A2(n28042), .ZN(N30321));
    NOR2X1 U17450 (.A1(n12932), .A2(n17878), .ZN(N30322));
    INVX1 U17451 (.I(n23132), .ZN(N30323));
    INVX1 U17452 (.I(n21988), .ZN(n30324));
    NANDX1 U17453 (.A1(n20016), .A2(N6217), .ZN(N30325));
    NANDX1 U17454 (.A1(N12161), .A2(N4419), .ZN(N30326));
    NOR2X1 U17455 (.A1(n26752), .A2(N3367), .ZN(n30327));
    INVX1 U17456 (.I(N6545), .ZN(n30328));
    INVX1 U17457 (.I(N9597), .ZN(n30329));
    INVX1 U17458 (.I(N12504), .ZN(N30330));
    INVX1 U17459 (.I(n15943), .ZN(N30331));
    NANDX1 U17460 (.A1(N11844), .A2(n23697), .ZN(n30332));
    NOR2X1 U17461 (.A1(N11959), .A2(n21197), .ZN(N30333));
    NANDX1 U17462 (.A1(n15792), .A2(n22689), .ZN(N30334));
    NOR2X1 U17463 (.A1(N6361), .A2(n15683), .ZN(n30335));
    NOR2X1 U17464 (.A1(n16909), .A2(n15133), .ZN(N30336));
    NANDX1 U17465 (.A1(N11686), .A2(N9082), .ZN(N30337));
    NANDX1 U17466 (.A1(n16105), .A2(N6544), .ZN(N30338));
    INVX1 U17467 (.I(N8032), .ZN(N30339));
    NOR2X1 U17468 (.A1(N8000), .A2(n15584), .ZN(n30340));
    INVX1 U17469 (.I(N11184), .ZN(N30341));
    INVX1 U17470 (.I(N2522), .ZN(n30342));
    NOR2X1 U17471 (.A1(N4969), .A2(n14365), .ZN(N30343));
    NANDX1 U17472 (.A1(n28044), .A2(n26323), .ZN(N30344));
    INVX1 U17473 (.I(n18886), .ZN(N30345));
    NOR2X1 U17474 (.A1(N11554), .A2(N4728), .ZN(n30346));
    NANDX1 U17475 (.A1(n27237), .A2(N11709), .ZN(N30347));
    NANDX1 U17476 (.A1(N793), .A2(n27267), .ZN(N30348));
    NOR2X1 U17477 (.A1(n28572), .A2(n13409), .ZN(n30349));
    INVX1 U17478 (.I(N4978), .ZN(N30350));
    INVX1 U17479 (.I(n25311), .ZN(n30351));
    NANDX1 U17480 (.A1(n22863), .A2(N10757), .ZN(N30352));
    NOR2X1 U17481 (.A1(N3909), .A2(N8707), .ZN(n30353));
    INVX1 U17482 (.I(n19595), .ZN(N30354));
    INVX1 U17483 (.I(N9680), .ZN(n30355));
    NANDX1 U17484 (.A1(N143), .A2(n24564), .ZN(n30356));
    NOR2X1 U17485 (.A1(N7590), .A2(n25102), .ZN(N30357));
    INVX1 U17486 (.I(N878), .ZN(N30358));
    INVX1 U17487 (.I(N3481), .ZN(N30359));
    NOR2X1 U17488 (.A1(n21489), .A2(N4273), .ZN(n30360));
    NANDX1 U17489 (.A1(N3966), .A2(N2707), .ZN(N30361));
    INVX1 U17490 (.I(n21245), .ZN(n30362));
    NOR2X1 U17491 (.A1(N3670), .A2(n16418), .ZN(N30363));
    NANDX1 U17492 (.A1(n26532), .A2(n27175), .ZN(N30364));
    NOR2X1 U17493 (.A1(n19001), .A2(n24442), .ZN(N30365));
    INVX1 U17494 (.I(n27157), .ZN(N30366));
    INVX1 U17495 (.I(n18259), .ZN(N30367));
    INVX1 U17496 (.I(n15382), .ZN(n30368));
    INVX1 U17497 (.I(n20687), .ZN(N30369));
    INVX1 U17498 (.I(n14908), .ZN(N30370));
    INVX1 U17499 (.I(N12409), .ZN(n30371));
    NOR2X1 U17500 (.A1(N11850), .A2(n13555), .ZN(N30372));
    INVX1 U17501 (.I(n16122), .ZN(N30373));
    NANDX1 U17502 (.A1(N7907), .A2(N7389), .ZN(N30374));
    NOR2X1 U17503 (.A1(n17712), .A2(n22331), .ZN(N30375));
    INVX1 U17504 (.I(N3993), .ZN(N30376));
    INVX1 U17505 (.I(N702), .ZN(N30377));
    NOR2X1 U17506 (.A1(n14487), .A2(N8263), .ZN(N30378));
    NOR2X1 U17507 (.A1(n23065), .A2(N5282), .ZN(n30379));
    NANDX1 U17508 (.A1(n29884), .A2(n19702), .ZN(n30380));
    NANDX1 U17509 (.A1(N992), .A2(n28950), .ZN(N30381));
    NANDX1 U17510 (.A1(n15899), .A2(N7182), .ZN(N30382));
    NOR2X1 U17511 (.A1(N9790), .A2(n19032), .ZN(N30383));
    NOR2X1 U17512 (.A1(n13731), .A2(n23714), .ZN(n30384));
    NANDX1 U17513 (.A1(N10198), .A2(n19664), .ZN(n30385));
    NANDX1 U17514 (.A1(n27909), .A2(N418), .ZN(N30386));
    NOR2X1 U17515 (.A1(n20462), .A2(N1641), .ZN(n30387));
    NOR2X1 U17516 (.A1(N10052), .A2(n16127), .ZN(n30388));
    NANDX1 U17517 (.A1(N12645), .A2(n27753), .ZN(N30389));
    NOR2X1 U17518 (.A1(N11778), .A2(n27499), .ZN(n30390));
    NOR2X1 U17519 (.A1(n14853), .A2(n28491), .ZN(N30391));
    NOR2X1 U17520 (.A1(n29459), .A2(N2813), .ZN(n30392));
    INVX1 U17521 (.I(n26336), .ZN(N30393));
    NANDX1 U17522 (.A1(N10284), .A2(n25328), .ZN(n30394));
    NOR2X1 U17523 (.A1(n22559), .A2(N6014), .ZN(N30395));
    INVX1 U17524 (.I(N646), .ZN(N30396));
    INVX1 U17525 (.I(n22862), .ZN(n30397));
    NOR2X1 U17526 (.A1(N3104), .A2(n13187), .ZN(N30398));
    NOR2X1 U17527 (.A1(n19571), .A2(N11799), .ZN(n30399));
    INVX1 U17528 (.I(N2725), .ZN(n30400));
    NOR2X1 U17529 (.A1(n23704), .A2(N9859), .ZN(N30401));
    NOR2X1 U17530 (.A1(N9627), .A2(n25255), .ZN(n30402));
    NANDX1 U17531 (.A1(n26678), .A2(N9326), .ZN(n30403));
    NANDX1 U17532 (.A1(n29490), .A2(N578), .ZN(N30404));
    NANDX1 U17533 (.A1(N516), .A2(n29560), .ZN(N30405));
    NANDX1 U17534 (.A1(n15409), .A2(n21981), .ZN(N30406));
    NOR2X1 U17535 (.A1(N10362), .A2(N11187), .ZN(N30407));
    INVX1 U17536 (.I(n21785), .ZN(n30408));
    INVX1 U17537 (.I(N3918), .ZN(n30409));
    NANDX1 U17538 (.A1(n22211), .A2(N12049), .ZN(n30410));
    NOR2X1 U17539 (.A1(N6724), .A2(N3335), .ZN(N30411));
    INVX1 U17540 (.I(N290), .ZN(N30412));
    NOR2X1 U17541 (.A1(N12840), .A2(n28614), .ZN(N30413));
    NANDX1 U17542 (.A1(N10897), .A2(n13715), .ZN(N30414));
    INVX1 U17543 (.I(n26972), .ZN(N30415));
    NANDX1 U17544 (.A1(N6773), .A2(N9109), .ZN(N30416));
    NANDX1 U17545 (.A1(n24893), .A2(N5134), .ZN(n30417));
    INVX1 U17546 (.I(n16736), .ZN(N30418));
    NOR2X1 U17547 (.A1(n16475), .A2(n16483), .ZN(N30419));
    NOR2X1 U17548 (.A1(N8122), .A2(n17293), .ZN(N30420));
    NANDX1 U17549 (.A1(n12955), .A2(n28064), .ZN(N30421));
    NOR2X1 U17550 (.A1(n18148), .A2(N4650), .ZN(n30422));
    NANDX1 U17551 (.A1(N6207), .A2(n23638), .ZN(n30423));
    INVX1 U17552 (.I(N7607), .ZN(N30424));
    NANDX1 U17553 (.A1(n21729), .A2(n18503), .ZN(n30425));
    NOR2X1 U17554 (.A1(n27924), .A2(N3899), .ZN(N30426));
    NANDX1 U17555 (.A1(n23257), .A2(N1568), .ZN(N30427));
    NOR2X1 U17556 (.A1(n18013), .A2(N6701), .ZN(N30428));
    INVX1 U17557 (.I(n23309), .ZN(n30429));
    NOR2X1 U17558 (.A1(N1914), .A2(n28353), .ZN(n30430));
    INVX1 U17559 (.I(N10035), .ZN(n30431));
    NANDX1 U17560 (.A1(n29580), .A2(N11551), .ZN(N30432));
    NOR2X1 U17561 (.A1(N516), .A2(n18259), .ZN(n30433));
    INVX1 U17562 (.I(n23621), .ZN(N30434));
    INVX1 U17563 (.I(N145), .ZN(N30435));
    INVX1 U17564 (.I(n20632), .ZN(n30436));
    NOR2X1 U17565 (.A1(N9933), .A2(n27696), .ZN(N30437));
    NOR2X1 U17566 (.A1(n26417), .A2(N1457), .ZN(N30438));
    NANDX1 U17567 (.A1(N8098), .A2(N3024), .ZN(n30439));
    NANDX1 U17568 (.A1(n26110), .A2(N9724), .ZN(N30440));
    NOR2X1 U17569 (.A1(N7842), .A2(N12156), .ZN(n30441));
    NOR2X1 U17570 (.A1(N6057), .A2(n22574), .ZN(N30442));
    NANDX1 U17571 (.A1(N10125), .A2(n22017), .ZN(N30443));
    NOR2X1 U17572 (.A1(N12120), .A2(N11093), .ZN(N30444));
    NOR2X1 U17573 (.A1(n18764), .A2(N4577), .ZN(n30445));
    INVX1 U17574 (.I(N7469), .ZN(N30446));
    INVX1 U17575 (.I(N6810), .ZN(N30447));
    NANDX1 U17576 (.A1(N2714), .A2(N4368), .ZN(N30448));
    NOR2X1 U17577 (.A1(n29130), .A2(N5824), .ZN(N30449));
    INVX1 U17578 (.I(N7090), .ZN(n30450));
    NANDX1 U17579 (.A1(N11843), .A2(n21760), .ZN(n30451));
    NANDX1 U17580 (.A1(n26393), .A2(n18163), .ZN(N30452));
    NANDX1 U17581 (.A1(N1279), .A2(n24219), .ZN(N30453));
    NANDX1 U17582 (.A1(n16337), .A2(N4207), .ZN(N30454));
    INVX1 U17583 (.I(N1369), .ZN(N30455));
    INVX1 U17584 (.I(N10515), .ZN(N30456));
    NANDX1 U17585 (.A1(n23650), .A2(n15091), .ZN(N30457));
    NOR2X1 U17586 (.A1(n19679), .A2(N7871), .ZN(N30458));
    NOR2X1 U17587 (.A1(N7828), .A2(n29282), .ZN(N30459));
    INVX1 U17588 (.I(N8307), .ZN(N30460));
    NANDX1 U17589 (.A1(n15097), .A2(n21176), .ZN(N30461));
    INVX1 U17590 (.I(N1065), .ZN(N30462));
    NOR2X1 U17591 (.A1(N4109), .A2(n26894), .ZN(N30463));
    NOR2X1 U17592 (.A1(n22271), .A2(N4604), .ZN(n30464));
    NOR2X1 U17593 (.A1(N4913), .A2(n23585), .ZN(n30465));
    INVX1 U17594 (.I(n27817), .ZN(N30466));
    NANDX1 U17595 (.A1(n25379), .A2(N2566), .ZN(N30467));
    NANDX1 U17596 (.A1(n18598), .A2(n14776), .ZN(N30468));
    NANDX1 U17597 (.A1(n16694), .A2(N4317), .ZN(N30469));
    INVX1 U17598 (.I(N2901), .ZN(N30470));
    NANDX1 U17599 (.A1(N2611), .A2(N12173), .ZN(N30471));
    INVX1 U17600 (.I(n19446), .ZN(n30472));
    NOR2X1 U17601 (.A1(n18748), .A2(N1794), .ZN(n30473));
    NANDX1 U17602 (.A1(N10190), .A2(N5902), .ZN(N30474));
    NOR2X1 U17603 (.A1(n28023), .A2(n16733), .ZN(n30475));
    INVX1 U17604 (.I(N5559), .ZN(N30476));
    INVX1 U17605 (.I(n18960), .ZN(N30477));
    NOR2X1 U17606 (.A1(n19325), .A2(N390), .ZN(n30478));
    INVX1 U17607 (.I(N10452), .ZN(N30479));
    NANDX1 U17608 (.A1(n20529), .A2(n25227), .ZN(N30480));
    NOR2X1 U17609 (.A1(N7085), .A2(n29544), .ZN(N30481));
    NANDX1 U17610 (.A1(N9985), .A2(N112), .ZN(n30482));
    NANDX1 U17611 (.A1(N10719), .A2(N9123), .ZN(n30483));
    NOR2X1 U17612 (.A1(n15109), .A2(n16432), .ZN(N30484));
    NOR2X1 U17613 (.A1(n20564), .A2(n26621), .ZN(N30485));
    INVX1 U17614 (.I(n22775), .ZN(n30486));
    INVX1 U17615 (.I(n26438), .ZN(N30487));
    NOR2X1 U17616 (.A1(n30065), .A2(n17946), .ZN(N30488));
    INVX1 U17617 (.I(n18057), .ZN(n30489));
    NANDX1 U17618 (.A1(n26060), .A2(N1290), .ZN(n30490));
    INVX1 U17619 (.I(n18394), .ZN(N30491));
    NOR2X1 U17620 (.A1(n19933), .A2(n17761), .ZN(n30492));
    INVX1 U17621 (.I(n19339), .ZN(N30493));
    INVX1 U17622 (.I(n27448), .ZN(n30494));
    NANDX1 U17623 (.A1(n14598), .A2(n26727), .ZN(N30495));
    INVX1 U17624 (.I(n28047), .ZN(N30496));
    NOR2X1 U17625 (.A1(N3428), .A2(n13153), .ZN(N30497));
    NOR2X1 U17626 (.A1(n18609), .A2(n22858), .ZN(N30498));
    NANDX1 U17627 (.A1(n12977), .A2(N7719), .ZN(N30499));
    INVX1 U17628 (.I(N1465), .ZN(N30500));
    INVX1 U17629 (.I(n27143), .ZN(n30501));
    INVX1 U17630 (.I(N9920), .ZN(N30502));
    NOR2X1 U17631 (.A1(N9371), .A2(N4626), .ZN(N30503));
    NOR2X1 U17632 (.A1(n19750), .A2(n24558), .ZN(N30504));
    NANDX1 U17633 (.A1(n18515), .A2(N2321), .ZN(N30505));
    NOR2X1 U17634 (.A1(N4386), .A2(N10331), .ZN(N30506));
    NANDX1 U17635 (.A1(n19674), .A2(n27464), .ZN(N30507));
    NANDX1 U17636 (.A1(n19933), .A2(n19452), .ZN(N30508));
    INVX1 U17637 (.I(N10618), .ZN(N30509));
    NOR2X1 U17638 (.A1(n18119), .A2(n24078), .ZN(N30510));
    INVX1 U17639 (.I(n25837), .ZN(n30511));
    INVX1 U17640 (.I(n29623), .ZN(n30512));
    NOR2X1 U17641 (.A1(n29815), .A2(N7568), .ZN(n30513));
    NANDX1 U17642 (.A1(N11304), .A2(N5499), .ZN(N30514));
    INVX1 U17643 (.I(N11186), .ZN(N30515));
    NOR2X1 U17644 (.A1(n26149), .A2(n17390), .ZN(n30516));
    INVX1 U17645 (.I(n28469), .ZN(N30517));
    INVX1 U17646 (.I(n25270), .ZN(n30518));
    NANDX1 U17647 (.A1(N9688), .A2(n14806), .ZN(N30519));
    INVX1 U17648 (.I(N3236), .ZN(N30520));
    NOR2X1 U17649 (.A1(N2562), .A2(N9936), .ZN(N30521));
    INVX1 U17650 (.I(n29183), .ZN(N30522));
    INVX1 U17651 (.I(n27857), .ZN(N30523));
    INVX1 U17652 (.I(n23754), .ZN(N30524));
    INVX1 U17653 (.I(n15250), .ZN(n30525));
    INVX1 U17654 (.I(n18767), .ZN(n30526));
    NOR2X1 U17655 (.A1(N507), .A2(n30071), .ZN(N30527));
    NOR2X1 U17656 (.A1(N2097), .A2(N11119), .ZN(N30528));
    NOR2X1 U17657 (.A1(n28245), .A2(n17069), .ZN(N30529));
    NANDX1 U17658 (.A1(n15137), .A2(n26938), .ZN(N30530));
    NANDX1 U17659 (.A1(n23799), .A2(n25187), .ZN(N30531));
    INVX1 U17660 (.I(N6909), .ZN(N30532));
    INVX1 U17661 (.I(n13091), .ZN(N30533));
    NANDX1 U17662 (.A1(N8221), .A2(n16869), .ZN(N30534));
    NANDX1 U17663 (.A1(n24835), .A2(N3149), .ZN(n30535));
    NANDX1 U17664 (.A1(N7012), .A2(n22238), .ZN(N30536));
    NOR2X1 U17665 (.A1(n29251), .A2(N10868), .ZN(N30537));
    NANDX1 U17666 (.A1(n29757), .A2(N10801), .ZN(n30538));
    NANDX1 U17667 (.A1(N1716), .A2(N10480), .ZN(N30539));
    NOR2X1 U17668 (.A1(n18522), .A2(n27549), .ZN(N30540));
    INVX1 U17669 (.I(N3521), .ZN(n30541));
    NOR2X1 U17670 (.A1(N294), .A2(n27319), .ZN(n30542));
    NOR2X1 U17671 (.A1(N8784), .A2(n22788), .ZN(n30543));
    INVX1 U17672 (.I(n21874), .ZN(N30544));
    NOR2X1 U17673 (.A1(N3025), .A2(n27303), .ZN(N30545));
    INVX1 U17674 (.I(n27859), .ZN(N30546));
    NOR2X1 U17675 (.A1(N597), .A2(n23432), .ZN(n30547));
    NANDX1 U17676 (.A1(n28686), .A2(n22545), .ZN(n30548));
    INVX1 U17677 (.I(n26576), .ZN(n30549));
    NANDX1 U17678 (.A1(N2643), .A2(n29904), .ZN(n30550));
    NOR2X1 U17679 (.A1(N1684), .A2(N3642), .ZN(N30551));
    NANDX1 U17680 (.A1(n29232), .A2(n17509), .ZN(n30552));
    INVX1 U17681 (.I(N565), .ZN(N30553));
    NANDX1 U17682 (.A1(n20224), .A2(N8524), .ZN(N30554));
    NANDX1 U17683 (.A1(N1436), .A2(N3328), .ZN(n30555));
    NOR2X1 U17684 (.A1(n22254), .A2(N6352), .ZN(n30556));
    NANDX1 U17685 (.A1(n28708), .A2(n22771), .ZN(N30557));
    NANDX1 U17686 (.A1(n29304), .A2(n16065), .ZN(n30558));
    INVX1 U17687 (.I(n16413), .ZN(N30559));
    NANDX1 U17688 (.A1(N3136), .A2(N1413), .ZN(N30560));
    NOR2X1 U17689 (.A1(n24477), .A2(N1179), .ZN(N30561));
    INVX1 U17690 (.I(n26160), .ZN(n30562));
    NOR2X1 U17691 (.A1(N9581), .A2(n13815), .ZN(n30563));
    NANDX1 U17692 (.A1(n13925), .A2(n14379), .ZN(N30564));
    NOR2X1 U17693 (.A1(n22710), .A2(N11463), .ZN(n30565));
    NANDX1 U17694 (.A1(n24145), .A2(n14790), .ZN(n30566));
    INVX1 U17695 (.I(N4822), .ZN(n30567));
    INVX1 U17696 (.I(n16265), .ZN(n30568));
    NANDX1 U17697 (.A1(N2336), .A2(n16446), .ZN(n30569));
    NANDX1 U17698 (.A1(N6961), .A2(n27739), .ZN(n30570));
    NOR2X1 U17699 (.A1(N3994), .A2(n19435), .ZN(n30571));
    NANDX1 U17700 (.A1(N11750), .A2(n13774), .ZN(N30572));
    INVX1 U17701 (.I(N1809), .ZN(n30573));
    NANDX1 U17702 (.A1(n22200), .A2(N11390), .ZN(n30574));
    NOR2X1 U17703 (.A1(N2951), .A2(n13875), .ZN(N30575));
    NOR2X1 U17704 (.A1(n20201), .A2(n25145), .ZN(n30576));
    NANDX1 U17705 (.A1(N11020), .A2(n19152), .ZN(N30577));
    NOR2X1 U17706 (.A1(n15979), .A2(N12534), .ZN(N30578));
    INVX1 U17707 (.I(N2107), .ZN(N30579));
    NANDX1 U17708 (.A1(N11823), .A2(N7113), .ZN(N30580));
    NOR2X1 U17709 (.A1(n18784), .A2(n23412), .ZN(n30581));
    NOR2X1 U17710 (.A1(n22777), .A2(N12709), .ZN(N30582));
    NANDX1 U17711 (.A1(N4389), .A2(n15044), .ZN(n30583));
    NANDX1 U17712 (.A1(N6198), .A2(n13400), .ZN(N30584));
    NOR2X1 U17713 (.A1(N6148), .A2(n14132), .ZN(N30585));
    NANDX1 U17714 (.A1(n20022), .A2(n29242), .ZN(N30586));
    NOR2X1 U17715 (.A1(n15030), .A2(n14238), .ZN(n30587));
    NANDX1 U17716 (.A1(n22742), .A2(n14024), .ZN(N30588));
    NOR2X1 U17717 (.A1(N5139), .A2(N4814), .ZN(N30589));
    NOR2X1 U17718 (.A1(N9625), .A2(n16636), .ZN(N30590));
    INVX1 U17719 (.I(n16669), .ZN(N30591));
    NOR2X1 U17720 (.A1(n28409), .A2(N8366), .ZN(N30592));
    INVX1 U17721 (.I(n29678), .ZN(N30593));
    NANDX1 U17722 (.A1(n21008), .A2(n14584), .ZN(n30594));
    NANDX1 U17723 (.A1(n27205), .A2(n16545), .ZN(N30595));
    NANDX1 U17724 (.A1(n21913), .A2(N539), .ZN(N30596));
    NOR2X1 U17725 (.A1(N358), .A2(n18341), .ZN(N30597));
    NOR2X1 U17726 (.A1(n15387), .A2(N2441), .ZN(N30598));
    NANDX1 U17727 (.A1(n26690), .A2(N5026), .ZN(n30599));
    NANDX1 U17728 (.A1(n20389), .A2(N9839), .ZN(n30600));
    INVX1 U17729 (.I(n30013), .ZN(N30601));
    NANDX1 U17730 (.A1(N1570), .A2(n16544), .ZN(N30602));
    NOR2X1 U17731 (.A1(n18539), .A2(n24909), .ZN(N30603));
    INVX1 U17732 (.I(n18079), .ZN(n30604));
    INVX1 U17733 (.I(n16366), .ZN(N30605));
    NANDX1 U17734 (.A1(n19368), .A2(N1994), .ZN(n30606));
    NANDX1 U17735 (.A1(n14904), .A2(n23906), .ZN(n30607));
    INVX1 U17736 (.I(N4776), .ZN(N30608));
    NOR2X1 U17737 (.A1(n15070), .A2(n16445), .ZN(N30609));
    NANDX1 U17738 (.A1(N6071), .A2(n19353), .ZN(n30610));
    NANDX1 U17739 (.A1(N11096), .A2(n29479), .ZN(N30611));
    INVX1 U17740 (.I(N9495), .ZN(N30612));
    NOR2X1 U17741 (.A1(N3450), .A2(n13091), .ZN(N30613));
    INVX1 U17742 (.I(N8554), .ZN(n30614));
    INVX1 U17743 (.I(n16021), .ZN(N30615));
    INVX1 U17744 (.I(n17326), .ZN(N30616));
    NOR2X1 U17745 (.A1(n14363), .A2(n22253), .ZN(N30617));
    NANDX1 U17746 (.A1(n22291), .A2(N12807), .ZN(N30618));
    NOR2X1 U17747 (.A1(N7057), .A2(N6576), .ZN(n30619));
    INVX1 U17748 (.I(N393), .ZN(N30620));
    NANDX1 U17749 (.A1(N3037), .A2(n16837), .ZN(N30621));
    INVX1 U17750 (.I(N9108), .ZN(N30622));
    INVX1 U17751 (.I(n19358), .ZN(N30623));
    NOR2X1 U17752 (.A1(n24091), .A2(n22932), .ZN(n30624));
    NANDX1 U17753 (.A1(n20004), .A2(n14943), .ZN(N30625));
    NOR2X1 U17754 (.A1(n17486), .A2(n23496), .ZN(n30626));
    INVX1 U17755 (.I(N3369), .ZN(N30627));
    NOR2X1 U17756 (.A1(n17626), .A2(N7331), .ZN(N30628));
    INVX1 U17757 (.I(N9741), .ZN(n30629));
    NANDX1 U17758 (.A1(n29156), .A2(N11109), .ZN(n30630));
    NOR2X1 U17759 (.A1(n24773), .A2(n17684), .ZN(N30631));
    NOR2X1 U17760 (.A1(n25166), .A2(n25644), .ZN(n30632));
    NANDX1 U17761 (.A1(N426), .A2(n20238), .ZN(N30633));
    NOR2X1 U17762 (.A1(n25176), .A2(N9458), .ZN(N30634));
    NANDX1 U17763 (.A1(N7690), .A2(n20951), .ZN(N30635));
    INVX1 U17764 (.I(n27694), .ZN(N30636));
    NANDX1 U17765 (.A1(n29219), .A2(n15042), .ZN(n30637));
    NANDX1 U17766 (.A1(N10821), .A2(n18411), .ZN(N30638));
    NANDX1 U17767 (.A1(n17008), .A2(n14302), .ZN(N30639));
    NOR2X1 U17768 (.A1(n15309), .A2(N5240), .ZN(n30640));
    INVX1 U17769 (.I(n26417), .ZN(N30641));
    INVX1 U17770 (.I(n22274), .ZN(N30642));
    NANDX1 U17771 (.A1(N10577), .A2(n17302), .ZN(N30643));
    INVX1 U17772 (.I(n25334), .ZN(N30644));
    NOR2X1 U17773 (.A1(n18268), .A2(n19061), .ZN(n30645));
    INVX1 U17774 (.I(n16286), .ZN(n30646));
    NANDX1 U17775 (.A1(n27714), .A2(N7099), .ZN(n30647));
    INVX1 U17776 (.I(n25270), .ZN(n30648));
    INVX1 U17777 (.I(N7064), .ZN(N30649));
    NOR2X1 U17778 (.A1(n19227), .A2(N6446), .ZN(N30650));
    NANDX1 U17779 (.A1(N10844), .A2(n23453), .ZN(N30651));
    INVX1 U17780 (.I(n20765), .ZN(N30652));
    NANDX1 U17781 (.A1(n13808), .A2(n18266), .ZN(n30653));
    NOR2X1 U17782 (.A1(N12664), .A2(n29101), .ZN(N30654));
    INVX1 U17783 (.I(N11801), .ZN(N30655));
    INVX1 U17784 (.I(N12716), .ZN(N30656));
    NOR2X1 U17785 (.A1(N11114), .A2(n19544), .ZN(n30657));
    NOR2X1 U17786 (.A1(N1001), .A2(N5692), .ZN(N30658));
    INVX1 U17787 (.I(n17276), .ZN(N30659));
    NOR2X1 U17788 (.A1(N2574), .A2(N969), .ZN(N30660));
    NOR2X1 U17789 (.A1(n28336), .A2(n29841), .ZN(n30661));
    NANDX1 U17790 (.A1(N4644), .A2(n24108), .ZN(N30662));
    INVX1 U17791 (.I(n16657), .ZN(N30663));
    NANDX1 U17792 (.A1(N585), .A2(N2402), .ZN(N30664));
    NANDX1 U17793 (.A1(N7411), .A2(n26003), .ZN(N30665));
    NOR2X1 U17794 (.A1(N6374), .A2(N10552), .ZN(N30666));
    NANDX1 U17795 (.A1(N11200), .A2(n23267), .ZN(N30667));
    INVX1 U17796 (.I(n22313), .ZN(N30668));
    NANDX1 U17797 (.A1(n20847), .A2(N11875), .ZN(N30669));
    NANDX1 U17798 (.A1(N3999), .A2(n29150), .ZN(N30670));
    INVX1 U17799 (.I(N6573), .ZN(N30671));
    NANDX1 U17800 (.A1(n29740), .A2(n23469), .ZN(N30672));
    INVX1 U17801 (.I(N10155), .ZN(N30673));
    INVX1 U17802 (.I(N914), .ZN(N30674));
    NANDX1 U17803 (.A1(N3192), .A2(N3453), .ZN(N30675));
    INVX1 U17804 (.I(N5593), .ZN(N30676));
    NANDX1 U17805 (.A1(N9408), .A2(n20157), .ZN(N30677));
    INVX1 U17806 (.I(n15782), .ZN(N30678));
    INVX1 U17807 (.I(n25163), .ZN(N30679));
    NANDX1 U17808 (.A1(N12398), .A2(N1255), .ZN(n30680));
    NANDX1 U17809 (.A1(n13631), .A2(N10662), .ZN(N30681));
    NOR2X1 U17810 (.A1(n20555), .A2(n14660), .ZN(N30682));
    NANDX1 U17811 (.A1(n17392), .A2(N9793), .ZN(N30683));
    INVX1 U17812 (.I(n16994), .ZN(n30684));
    INVX1 U17813 (.I(n21347), .ZN(N30685));
    NANDX1 U17814 (.A1(N8357), .A2(n22260), .ZN(n30686));
    INVX1 U17815 (.I(N109), .ZN(N30687));
    NOR2X1 U17816 (.A1(n19119), .A2(n24400), .ZN(N30688));
    NANDX1 U17817 (.A1(n17088), .A2(n14419), .ZN(N30689));
    NOR2X1 U17818 (.A1(N2732), .A2(N3550), .ZN(n30690));
    NANDX1 U17819 (.A1(n18273), .A2(n15947), .ZN(N30691));
    NANDX1 U17820 (.A1(n14550), .A2(n29577), .ZN(N30692));
    INVX1 U17821 (.I(N11263), .ZN(N30693));
    NANDX1 U17822 (.A1(n28585), .A2(N6987), .ZN(N30694));
    NOR2X1 U17823 (.A1(n26938), .A2(n21390), .ZN(n30695));
    INVX1 U17824 (.I(n18623), .ZN(N30696));
    NOR2X1 U17825 (.A1(n28511), .A2(n26979), .ZN(n30697));
    INVX1 U17826 (.I(n15495), .ZN(n30698));
    NANDX1 U17827 (.A1(n18994), .A2(n23175), .ZN(N30699));
    INVX1 U17828 (.I(N11489), .ZN(n30700));
    NOR2X1 U17829 (.A1(n24329), .A2(N11214), .ZN(n30701));
    NANDX1 U17830 (.A1(n27878), .A2(N5965), .ZN(n30702));
    NOR2X1 U17831 (.A1(n13687), .A2(n20667), .ZN(N30703));
    NOR2X1 U17832 (.A1(n13126), .A2(N4455), .ZN(N30704));
    NOR2X1 U17833 (.A1(n21680), .A2(n21600), .ZN(N30705));
    NANDX1 U17834 (.A1(N6050), .A2(N6961), .ZN(N30706));
    INVX1 U17835 (.I(n18851), .ZN(n30707));
    NANDX1 U17836 (.A1(n22021), .A2(N5785), .ZN(n30708));
    NANDX1 U17837 (.A1(N3864), .A2(n21280), .ZN(n30709));
    INVX1 U17838 (.I(n22857), .ZN(N30710));
    INVX1 U17839 (.I(n17846), .ZN(n30711));
    INVX1 U17840 (.I(n13002), .ZN(N30712));
    INVX1 U17841 (.I(N3983), .ZN(N30713));
    NANDX1 U17842 (.A1(n28475), .A2(N9947), .ZN(N30714));
    INVX1 U17843 (.I(N585), .ZN(n30715));
    NANDX1 U17844 (.A1(n22587), .A2(n13710), .ZN(N30716));
    NOR2X1 U17845 (.A1(n15072), .A2(n23950), .ZN(N30717));
    NOR2X1 U17846 (.A1(N3104), .A2(n29999), .ZN(N30718));
    INVX1 U17847 (.I(N12525), .ZN(N30719));
    INVX1 U17848 (.I(n13316), .ZN(n30720));
    NOR2X1 U17849 (.A1(N1619), .A2(n24301), .ZN(N30721));
    INVX1 U17850 (.I(n22898), .ZN(n30722));
    NANDX1 U17851 (.A1(N8250), .A2(n14336), .ZN(n30723));
    NOR2X1 U17852 (.A1(N1018), .A2(n27337), .ZN(N30724));
    NOR2X1 U17853 (.A1(N5000), .A2(N178), .ZN(N30725));
    INVX1 U17854 (.I(N3507), .ZN(N30726));
    NOR2X1 U17855 (.A1(n15282), .A2(N11242), .ZN(N30727));
    NOR2X1 U17856 (.A1(n17552), .A2(N11991), .ZN(n30728));
    NOR2X1 U17857 (.A1(n30063), .A2(N4203), .ZN(n30729));
    INVX1 U17858 (.I(n18485), .ZN(N30730));
    NANDX1 U17859 (.A1(N11675), .A2(n14319), .ZN(N30731));
    NANDX1 U17860 (.A1(n23342), .A2(n15938), .ZN(N30732));
    NOR2X1 U17861 (.A1(n20173), .A2(n27396), .ZN(n30733));
    INVX1 U17862 (.I(n28422), .ZN(n30734));
    INVX1 U17863 (.I(n24536), .ZN(N30735));
    NOR2X1 U17864 (.A1(n27492), .A2(n29457), .ZN(n30736));
    INVX1 U17865 (.I(n27670), .ZN(N30737));
    NANDX1 U17866 (.A1(n15068), .A2(n16196), .ZN(n30738));
    NOR2X1 U17867 (.A1(n14870), .A2(n27309), .ZN(N30739));
    INVX1 U17868 (.I(n26860), .ZN(n30740));
    NOR2X1 U17869 (.A1(n23898), .A2(N925), .ZN(N30741));
    INVX1 U17870 (.I(N12245), .ZN(N30742));
    INVX1 U17871 (.I(n22742), .ZN(N30743));
    NOR2X1 U17872 (.A1(n28248), .A2(n15946), .ZN(N30744));
    NOR2X1 U17873 (.A1(n16223), .A2(n24679), .ZN(n30745));
    INVX1 U17874 (.I(n13555), .ZN(n30746));
    NANDX1 U17875 (.A1(N9777), .A2(N7953), .ZN(N30747));
    INVX1 U17876 (.I(n25830), .ZN(n30748));
    NANDX1 U17877 (.A1(N10948), .A2(N11923), .ZN(N30749));
    INVX1 U17878 (.I(n26015), .ZN(N30750));
    NANDX1 U17879 (.A1(n27710), .A2(N10747), .ZN(N30751));
    NOR2X1 U17880 (.A1(n21545), .A2(n26168), .ZN(n30752));
    NOR2X1 U17881 (.A1(N3866), .A2(n27092), .ZN(N30753));
    INVX1 U17882 (.I(N4672), .ZN(n30754));
    NANDX1 U17883 (.A1(n29438), .A2(n19796), .ZN(N30755));
    NANDX1 U17884 (.A1(N3807), .A2(n20720), .ZN(N30756));
    INVX1 U17885 (.I(n28485), .ZN(n30757));
    NOR2X1 U17886 (.A1(N6262), .A2(N9872), .ZN(N30758));
    NANDX1 U17887 (.A1(N2776), .A2(n27957), .ZN(N30759));
    NANDX1 U17888 (.A1(n28746), .A2(N8768), .ZN(n30760));
    NOR2X1 U17889 (.A1(N8459), .A2(n23343), .ZN(N30761));
    INVX1 U17890 (.I(n24729), .ZN(n30762));
    NOR2X1 U17891 (.A1(n25245), .A2(N4698), .ZN(N30763));
    NANDX1 U17892 (.A1(N2177), .A2(n27261), .ZN(n30764));
    NANDX1 U17893 (.A1(n20312), .A2(N1795), .ZN(n30765));
    INVX1 U17894 (.I(n19612), .ZN(N30766));
    INVX1 U17895 (.I(N632), .ZN(N30767));
    NOR2X1 U17896 (.A1(N733), .A2(N12037), .ZN(N30768));
    INVX1 U17897 (.I(n26894), .ZN(N30769));
    NANDX1 U17898 (.A1(N8759), .A2(N2557), .ZN(n30770));
    INVX1 U17899 (.I(N6578), .ZN(n30771));
    NOR2X1 U17900 (.A1(N8243), .A2(n15345), .ZN(N30772));
    NANDX1 U17901 (.A1(N5262), .A2(N8551), .ZN(N30773));
    NOR2X1 U17902 (.A1(n18551), .A2(N1064), .ZN(N30774));
    INVX1 U17903 (.I(N11809), .ZN(n30775));
    NANDX1 U17904 (.A1(n21961), .A2(n27631), .ZN(n30776));
    INVX1 U17905 (.I(N696), .ZN(N30777));
    NANDX1 U17906 (.A1(n17949), .A2(n20307), .ZN(n30778));
    NOR2X1 U17907 (.A1(N7141), .A2(N2148), .ZN(N30779));
    NANDX1 U17908 (.A1(N7739), .A2(N1034), .ZN(N30780));
    NANDX1 U17909 (.A1(n14598), .A2(N9792), .ZN(N30781));
    NANDX1 U17910 (.A1(n24232), .A2(n16370), .ZN(N30782));
    INVX1 U17911 (.I(n21035), .ZN(n30783));
    NANDX1 U17912 (.A1(N3935), .A2(n14857), .ZN(N30784));
    NOR2X1 U17913 (.A1(N9914), .A2(n21968), .ZN(N30785));
    INVX1 U17914 (.I(n29698), .ZN(N30786));
    INVX1 U17915 (.I(N8055), .ZN(N30787));
    NOR2X1 U17916 (.A1(n19831), .A2(n20555), .ZN(n30788));
    NANDX1 U17917 (.A1(N7679), .A2(n27064), .ZN(N30789));
    NANDX1 U17918 (.A1(N5678), .A2(n22765), .ZN(N30790));
    NANDX1 U17919 (.A1(n23108), .A2(N366), .ZN(N30791));
    NANDX1 U17920 (.A1(N7156), .A2(N3524), .ZN(N30792));
    NOR2X1 U17921 (.A1(N12459), .A2(n16316), .ZN(N30793));
    INVX1 U17922 (.I(n21809), .ZN(N30794));
    NOR2X1 U17923 (.A1(n16244), .A2(n14305), .ZN(N30795));
    NOR2X1 U17924 (.A1(N3493), .A2(N12779), .ZN(N30796));
    INVX1 U17925 (.I(n21941), .ZN(n30797));
    INVX1 U17926 (.I(n13359), .ZN(n30798));
    NOR2X1 U17927 (.A1(N10981), .A2(n21750), .ZN(n30799));
    NOR2X1 U17928 (.A1(n21757), .A2(n29428), .ZN(n30800));
    NOR2X1 U17929 (.A1(N11263), .A2(N4969), .ZN(N30801));
    NOR2X1 U17930 (.A1(n21614), .A2(n28076), .ZN(n30802));
    NOR2X1 U17931 (.A1(n21559), .A2(N5094), .ZN(N30803));
    INVX1 U17932 (.I(N1159), .ZN(N30804));
    NOR2X1 U17933 (.A1(n25991), .A2(n27265), .ZN(n30805));
    NOR2X1 U17934 (.A1(n21764), .A2(N1933), .ZN(N30806));
    NOR2X1 U17935 (.A1(n20955), .A2(N5425), .ZN(n30807));
    NANDX1 U17936 (.A1(N11976), .A2(n15926), .ZN(N30808));
    NOR2X1 U17937 (.A1(n13895), .A2(N4345), .ZN(N30809));
    NANDX1 U17938 (.A1(N5507), .A2(N1879), .ZN(N30810));
    NOR2X1 U17939 (.A1(N4797), .A2(n15037), .ZN(n30811));
    NANDX1 U17940 (.A1(n28463), .A2(N2125), .ZN(n30812));
    NANDX1 U17941 (.A1(n26401), .A2(n26974), .ZN(N30813));
    NOR2X1 U17942 (.A1(n20056), .A2(N6511), .ZN(n30814));
    NANDX1 U17943 (.A1(n26168), .A2(n21062), .ZN(N30815));
    INVX1 U17944 (.I(N12513), .ZN(N30816));
    NOR2X1 U17945 (.A1(N2943), .A2(N1723), .ZN(N30817));
    NOR2X1 U17946 (.A1(N8367), .A2(n15150), .ZN(N30818));
    INVX1 U17947 (.I(n24293), .ZN(N30819));
    INVX1 U17948 (.I(n17936), .ZN(n30820));
    INVX1 U17949 (.I(n20465), .ZN(n30821));
    NOR2X1 U17950 (.A1(N7638), .A2(n14512), .ZN(N30822));
    NANDX1 U17951 (.A1(n22674), .A2(n27080), .ZN(N30823));
    NOR2X1 U17952 (.A1(n13359), .A2(N987), .ZN(N30824));
    INVX1 U17953 (.I(N10195), .ZN(n30825));
    NOR2X1 U17954 (.A1(N8565), .A2(n16706), .ZN(N30826));
    NANDX1 U17955 (.A1(n23294), .A2(n26328), .ZN(N30827));
    NANDX1 U17956 (.A1(N5669), .A2(N8879), .ZN(N30828));
    NANDX1 U17957 (.A1(N7392), .A2(N945), .ZN(N30829));
    NANDX1 U17958 (.A1(N11102), .A2(N4986), .ZN(n30830));
    NOR2X1 U17959 (.A1(n17700), .A2(N11482), .ZN(n30831));
    NANDX1 U17960 (.A1(N8027), .A2(n23484), .ZN(N30832));
    NOR2X1 U17961 (.A1(N11100), .A2(n28844), .ZN(N30833));
    INVX1 U17962 (.I(n26740), .ZN(N30834));
    NOR2X1 U17963 (.A1(N3223), .A2(n27727), .ZN(n30835));
    INVX1 U17964 (.I(N1978), .ZN(N30836));
    INVX1 U17965 (.I(n29603), .ZN(N30837));
    NANDX1 U17966 (.A1(n13075), .A2(n22759), .ZN(N30838));
    NANDX1 U17967 (.A1(n14420), .A2(n16988), .ZN(N30839));
    NOR2X1 U17968 (.A1(n18708), .A2(n24379), .ZN(N30840));
    NOR2X1 U17969 (.A1(N1226), .A2(n24042), .ZN(n30841));
    NANDX1 U17970 (.A1(n26733), .A2(N11604), .ZN(N30842));
    NOR2X1 U17971 (.A1(n27862), .A2(N8191), .ZN(N30843));
    NOR2X1 U17972 (.A1(n25189), .A2(N7851), .ZN(n30844));
    NOR2X1 U17973 (.A1(N3614), .A2(N4454), .ZN(N30845));
    NANDX1 U17974 (.A1(N6836), .A2(n20741), .ZN(N30846));
    NOR2X1 U17975 (.A1(n27511), .A2(N3343), .ZN(N30847));
    NOR2X1 U17976 (.A1(N4618), .A2(N4978), .ZN(n30848));
    NOR2X1 U17977 (.A1(N8052), .A2(n19397), .ZN(N30849));
    NOR2X1 U17978 (.A1(N8925), .A2(n26666), .ZN(N30850));
    NOR2X1 U17979 (.A1(N10743), .A2(n27891), .ZN(N30851));
    NOR2X1 U17980 (.A1(n24806), .A2(n13047), .ZN(N30852));
    NOR2X1 U17981 (.A1(N1515), .A2(n29470), .ZN(N30853));
    NANDX1 U17982 (.A1(N8966), .A2(n13082), .ZN(n30854));
    INVX1 U17983 (.I(n15124), .ZN(N30855));
    INVX1 U17984 (.I(n20406), .ZN(N30856));
    INVX1 U17985 (.I(N12091), .ZN(n30857));
    INVX1 U17986 (.I(N11682), .ZN(N30858));
    INVX1 U17987 (.I(N2912), .ZN(n30859));
    NOR2X1 U17988 (.A1(n14082), .A2(n26587), .ZN(n30860));
    NANDX1 U17989 (.A1(N10694), .A2(N4407), .ZN(N30861));
    NANDX1 U17990 (.A1(n19618), .A2(N935), .ZN(N30862));
    NANDX1 U17991 (.A1(n18922), .A2(n17386), .ZN(N30863));
    INVX1 U17992 (.I(n13590), .ZN(N30864));
    NOR2X1 U17993 (.A1(n23414), .A2(N3665), .ZN(N30865));
    NANDX1 U17994 (.A1(N12817), .A2(N1191), .ZN(N30866));
    NANDX1 U17995 (.A1(n17330), .A2(n16314), .ZN(n30867));
    NOR2X1 U17996 (.A1(N7598), .A2(n28547), .ZN(n30868));
    NANDX1 U17997 (.A1(n25865), .A2(n28789), .ZN(N30869));
    NANDX1 U17998 (.A1(n28776), .A2(N5068), .ZN(n30870));
    NANDX1 U17999 (.A1(n13786), .A2(n21716), .ZN(N30871));
    NANDX1 U18000 (.A1(n18193), .A2(N12570), .ZN(N30872));
    INVX1 U18001 (.I(N7688), .ZN(N30873));
    NOR2X1 U18002 (.A1(N8241), .A2(n25074), .ZN(n30874));
    INVX1 U18003 (.I(N10391), .ZN(N30875));
    INVX1 U18004 (.I(n26045), .ZN(N30876));
    INVX1 U18005 (.I(N2118), .ZN(N30877));
    INVX1 U18006 (.I(N3806), .ZN(n30878));
    INVX1 U18007 (.I(n14615), .ZN(N30879));
    NOR2X1 U18008 (.A1(N9912), .A2(N10774), .ZN(N30880));
    INVX1 U18009 (.I(n28528), .ZN(N30881));
    INVX1 U18010 (.I(n13000), .ZN(N30882));
    NANDX1 U18011 (.A1(n23838), .A2(n18067), .ZN(N30883));
    NANDX1 U18012 (.A1(n26184), .A2(n28344), .ZN(n30884));
    INVX1 U18013 (.I(n14239), .ZN(N30885));
    NANDX1 U18014 (.A1(n27651), .A2(N10488), .ZN(N30886));
    NOR2X1 U18015 (.A1(N5754), .A2(n24122), .ZN(N30887));
    NOR2X1 U18016 (.A1(N4705), .A2(N7914), .ZN(N30888));
    NANDX1 U18017 (.A1(N7320), .A2(n28729), .ZN(n30889));
    NOR2X1 U18018 (.A1(n29824), .A2(n20676), .ZN(N30890));
    NANDX1 U18019 (.A1(N8367), .A2(n19149), .ZN(n30891));
    NOR2X1 U18020 (.A1(N4017), .A2(N6100), .ZN(n30892));
    INVX1 U18021 (.I(N5577), .ZN(N30893));
    NOR2X1 U18022 (.A1(N7138), .A2(n23644), .ZN(n30894));
    NANDX1 U18023 (.A1(N3184), .A2(N10411), .ZN(N30895));
    NOR2X1 U18024 (.A1(N5984), .A2(N9747), .ZN(N30896));
    INVX1 U18025 (.I(n16471), .ZN(n30897));
    NANDX1 U18026 (.A1(n29509), .A2(n29153), .ZN(N30898));
    NOR2X1 U18027 (.A1(n22774), .A2(N6929), .ZN(n30899));
    INVX1 U18028 (.I(n30094), .ZN(N30900));
    NANDX1 U18029 (.A1(n26636), .A2(n29780), .ZN(N30901));
    NANDX1 U18030 (.A1(N4101), .A2(n26707), .ZN(N30902));
    INVX1 U18031 (.I(n22477), .ZN(N30903));
    NOR2X1 U18032 (.A1(n28564), .A2(N5777), .ZN(N30904));
    NANDX1 U18033 (.A1(n19557), .A2(N1475), .ZN(N30905));
    INVX1 U18034 (.I(n26164), .ZN(n30906));
    NANDX1 U18035 (.A1(n28776), .A2(n22268), .ZN(N30907));
    NOR2X1 U18036 (.A1(N8386), .A2(n15886), .ZN(N30908));
    INVX1 U18037 (.I(N8037), .ZN(n30909));
    INVX1 U18038 (.I(N3248), .ZN(n30910));
    NANDX1 U18039 (.A1(n26591), .A2(n28874), .ZN(n30911));
    NOR2X1 U18040 (.A1(n15108), .A2(n22954), .ZN(N30912));
    NOR2X1 U18041 (.A1(N3311), .A2(n26271), .ZN(N30913));
    NANDX1 U18042 (.A1(n30017), .A2(n18598), .ZN(N30914));
    INVX1 U18043 (.I(N7724), .ZN(N30915));
    NANDX1 U18044 (.A1(n16967), .A2(N2447), .ZN(N30916));
    NANDX1 U18045 (.A1(n18441), .A2(N9373), .ZN(N30917));
    NOR2X1 U18046 (.A1(N11659), .A2(N8012), .ZN(N30918));
    NANDX1 U18047 (.A1(n29559), .A2(N4958), .ZN(N30919));
    NOR2X1 U18048 (.A1(N3654), .A2(N1555), .ZN(n30920));
    INVX1 U18049 (.I(n25600), .ZN(N30921));
    NANDX1 U18050 (.A1(n25274), .A2(n24336), .ZN(N30922));
    INVX1 U18051 (.I(n28943), .ZN(N30923));
    NOR2X1 U18052 (.A1(n20265), .A2(n20814), .ZN(n30924));
    INVX1 U18053 (.I(n20418), .ZN(N30925));
    NANDX1 U18054 (.A1(n20444), .A2(n12910), .ZN(N30926));
    NANDX1 U18055 (.A1(n14590), .A2(n18437), .ZN(n30927));
    NOR2X1 U18056 (.A1(n16853), .A2(n25438), .ZN(n30928));
    NOR2X1 U18057 (.A1(n15143), .A2(n25657), .ZN(n30929));
    INVX1 U18058 (.I(N5563), .ZN(N30930));
    NOR2X1 U18059 (.A1(N189), .A2(N429), .ZN(n30931));
    INVX1 U18060 (.I(n20441), .ZN(n30932));
    NOR2X1 U18061 (.A1(N12755), .A2(n22220), .ZN(N30933));
    INVX1 U18062 (.I(N6953), .ZN(N30934));
    NOR2X1 U18063 (.A1(N11751), .A2(n24105), .ZN(N30935));
    NANDX1 U18064 (.A1(N2428), .A2(n25951), .ZN(N30936));
    NANDX1 U18065 (.A1(N11682), .A2(N4819), .ZN(N30937));
    NOR2X1 U18066 (.A1(n28659), .A2(N7969), .ZN(n30938));
    INVX1 U18067 (.I(N6507), .ZN(N30939));
    NANDX1 U18068 (.A1(n19167), .A2(N5166), .ZN(n30940));
    NOR2X1 U18069 (.A1(n14686), .A2(N397), .ZN(n30941));
    NOR2X1 U18070 (.A1(n28325), .A2(n19283), .ZN(N30942));
    NANDX1 U18071 (.A1(n15480), .A2(N9586), .ZN(n30943));
    INVX1 U18072 (.I(n28234), .ZN(N30944));
    INVX1 U18073 (.I(N4995), .ZN(N30945));
    NANDX1 U18074 (.A1(n25222), .A2(n16746), .ZN(N30946));
    NOR2X1 U18075 (.A1(n20204), .A2(N7734), .ZN(N30947));
    INVX1 U18076 (.I(N5466), .ZN(N30948));
    NANDX1 U18077 (.A1(n25605), .A2(n22335), .ZN(N30949));
    INVX1 U18078 (.I(N3437), .ZN(N30950));
    NOR2X1 U18079 (.A1(N1564), .A2(n16819), .ZN(n30951));
    NOR2X1 U18080 (.A1(n25427), .A2(n15206), .ZN(N30952));
    NANDX1 U18081 (.A1(n25823), .A2(n19155), .ZN(N30953));
    NOR2X1 U18082 (.A1(N3529), .A2(N12093), .ZN(n30954));
    INVX1 U18083 (.I(N1676), .ZN(n30955));
    NOR2X1 U18084 (.A1(n27360), .A2(n22042), .ZN(n30956));
    INVX1 U18085 (.I(N9531), .ZN(N30957));
    NOR2X1 U18086 (.A1(n25881), .A2(n15806), .ZN(n30958));
    INVX1 U18087 (.I(n22175), .ZN(N30959));
    NOR2X1 U18088 (.A1(N12657), .A2(N13), .ZN(N30960));
    NOR2X1 U18089 (.A1(n23552), .A2(n13769), .ZN(n30961));
    NOR2X1 U18090 (.A1(n28176), .A2(N3893), .ZN(N30962));
    INVX1 U18091 (.I(n21829), .ZN(N30963));
    NOR2X1 U18092 (.A1(n14504), .A2(n18728), .ZN(N30964));
    NANDX1 U18093 (.A1(n22219), .A2(n13815), .ZN(N30965));
    INVX1 U18094 (.I(N4174), .ZN(N30966));
    NOR2X1 U18095 (.A1(n18770), .A2(N8315), .ZN(n30967));
    NANDX1 U18096 (.A1(N10674), .A2(n17450), .ZN(N30968));
    NANDX1 U18097 (.A1(n27799), .A2(n13194), .ZN(n30969));
    NANDX1 U18098 (.A1(N4853), .A2(n23929), .ZN(N30970));
    NANDX1 U18099 (.A1(N6070), .A2(N12503), .ZN(N30971));
    INVX1 U18100 (.I(n29621), .ZN(N30972));
    INVX1 U18101 (.I(N10736), .ZN(n30973));
    INVX1 U18102 (.I(N26), .ZN(N30974));
    INVX1 U18103 (.I(N7911), .ZN(N30975));
    NOR2X1 U18104 (.A1(n13098), .A2(n26638), .ZN(N30976));
    NOR2X1 U18105 (.A1(n23877), .A2(n29013), .ZN(N30977));
    NOR2X1 U18106 (.A1(n28050), .A2(N11817), .ZN(n30978));
    NANDX1 U18107 (.A1(N6227), .A2(n29239), .ZN(N30979));
    NOR2X1 U18108 (.A1(N12238), .A2(n26054), .ZN(n30980));
    INVX1 U18109 (.I(n13992), .ZN(N30981));
    NANDX1 U18110 (.A1(n20247), .A2(N7783), .ZN(N30982));
    NOR2X1 U18111 (.A1(n26316), .A2(n20285), .ZN(N30983));
    NANDX1 U18112 (.A1(n14360), .A2(N4979), .ZN(n30984));
    NANDX1 U18113 (.A1(N442), .A2(N5005), .ZN(n30985));
    NOR2X1 U18114 (.A1(n27050), .A2(n22910), .ZN(N30986));
    INVX1 U18115 (.I(n23550), .ZN(N30987));
    INVX1 U18116 (.I(n26278), .ZN(N30988));
    NOR2X1 U18117 (.A1(n23974), .A2(n24190), .ZN(n30989));
    NOR2X1 U18118 (.A1(N897), .A2(n18978), .ZN(n30990));
    INVX1 U18119 (.I(n18630), .ZN(N30991));
    INVX1 U18120 (.I(n17820), .ZN(N30992));
    NANDX1 U18121 (.A1(N3630), .A2(n14917), .ZN(N30993));
    NANDX1 U18122 (.A1(N11412), .A2(n19649), .ZN(N30994));
    NOR2X1 U18123 (.A1(n20258), .A2(n22500), .ZN(n30995));
    NOR2X1 U18124 (.A1(n25236), .A2(n24648), .ZN(n30996));
    NOR2X1 U18125 (.A1(n18801), .A2(n13951), .ZN(n30997));
    NOR2X1 U18126 (.A1(N135), .A2(n16351), .ZN(N30998));
    NOR2X1 U18127 (.A1(n24378), .A2(N12491), .ZN(N30999));
    NOR2X1 U18128 (.A1(n18215), .A2(n25242), .ZN(N31000));
    NOR2X1 U18129 (.A1(N7672), .A2(n14082), .ZN(n31001));
    NOR2X1 U18130 (.A1(n26302), .A2(n22418), .ZN(n31002));
    INVX1 U18131 (.I(n18749), .ZN(N31003));
    NANDX1 U18132 (.A1(n26530), .A2(N1306), .ZN(N31004));
    INVX1 U18133 (.I(n16041), .ZN(N31005));
    INVX1 U18134 (.I(n16139), .ZN(N31006));
    INVX1 U18135 (.I(N10530), .ZN(N31007));
    NOR2X1 U18136 (.A1(N10173), .A2(N11323), .ZN(n31008));
    NOR2X1 U18137 (.A1(n24123), .A2(n27727), .ZN(N31009));
    INVX1 U18138 (.I(N10336), .ZN(N31010));
    NANDX1 U18139 (.A1(n12974), .A2(N11388), .ZN(n31011));
    INVX1 U18140 (.I(n19749), .ZN(n31012));
    NOR2X1 U18141 (.A1(n22977), .A2(n15981), .ZN(n31013));
    NOR2X1 U18142 (.A1(n16771), .A2(N12145), .ZN(n31014));
    NOR2X1 U18143 (.A1(n28384), .A2(N757), .ZN(n31015));
    INVX1 U18144 (.I(n13337), .ZN(N31016));
    NANDX1 U18145 (.A1(n23341), .A2(n17938), .ZN(N31017));
    NOR2X1 U18146 (.A1(N9343), .A2(n14902), .ZN(N31018));
    NANDX1 U18147 (.A1(N9141), .A2(n13635), .ZN(N31019));
    NOR2X1 U18148 (.A1(n27739), .A2(n26318), .ZN(N31020));
    INVX1 U18149 (.I(N4896), .ZN(N31021));
    NOR2X1 U18150 (.A1(n16206), .A2(n17869), .ZN(N31022));
    NANDX1 U18151 (.A1(n14276), .A2(n26178), .ZN(N31023));
    INVX1 U18152 (.I(n25813), .ZN(n31024));
    INVX1 U18153 (.I(n22089), .ZN(n31025));
    NANDX1 U18154 (.A1(N12727), .A2(n23502), .ZN(n31026));
    NANDX1 U18155 (.A1(N2044), .A2(N9385), .ZN(n31027));
    INVX1 U18156 (.I(n22803), .ZN(N31028));
    INVX1 U18157 (.I(N389), .ZN(N31029));
    INVX1 U18158 (.I(N491), .ZN(n31030));
    NANDX1 U18159 (.A1(N12051), .A2(n28329), .ZN(n31031));
    INVX1 U18160 (.I(N11823), .ZN(N31032));
    NOR2X1 U18161 (.A1(n13667), .A2(N9184), .ZN(N31033));
    INVX1 U18162 (.I(N8744), .ZN(n31034));
    NOR2X1 U18163 (.A1(N7118), .A2(n15208), .ZN(N31035));
    NANDX1 U18164 (.A1(n21856), .A2(n16724), .ZN(N31036));
    NANDX1 U18165 (.A1(N3739), .A2(N8675), .ZN(N31037));
    NOR2X1 U18166 (.A1(N5026), .A2(n20737), .ZN(N31038));
    NANDX1 U18167 (.A1(N7069), .A2(n18682), .ZN(N31039));
    NANDX1 U18168 (.A1(n29871), .A2(N9830), .ZN(n31040));
    NOR2X1 U18169 (.A1(N11896), .A2(N10321), .ZN(N31041));
    INVX1 U18170 (.I(n23946), .ZN(n31042));
    NOR2X1 U18171 (.A1(N5456), .A2(N5631), .ZN(N31043));
    NOR2X1 U18172 (.A1(N7683), .A2(n14814), .ZN(n31044));
    NOR2X1 U18173 (.A1(n16426), .A2(n17324), .ZN(N31045));
    NOR2X1 U18174 (.A1(n20194), .A2(n15411), .ZN(n31046));
    INVX1 U18175 (.I(N6780), .ZN(N31047));
    NOR2X1 U18176 (.A1(n22085), .A2(n15454), .ZN(N31048));
    NOR2X1 U18177 (.A1(n27110), .A2(n24751), .ZN(n31049));
    INVX1 U18178 (.I(N4042), .ZN(N31050));
    INVX1 U18179 (.I(N7648), .ZN(N31051));
    NANDX1 U18180 (.A1(n23124), .A2(n21903), .ZN(N31052));
    INVX1 U18181 (.I(n22005), .ZN(N31053));
    INVX1 U18182 (.I(n16737), .ZN(N31054));
    NANDX1 U18183 (.A1(n15328), .A2(N10928), .ZN(n31055));
    NANDX1 U18184 (.A1(n23010), .A2(n14302), .ZN(N31056));
    NOR2X1 U18185 (.A1(n27996), .A2(N1488), .ZN(N31057));
    NANDX1 U18186 (.A1(n18052), .A2(N5459), .ZN(N31058));
    INVX1 U18187 (.I(n13392), .ZN(N31059));
    NOR2X1 U18188 (.A1(N841), .A2(n17406), .ZN(n31060));
    NANDX1 U18189 (.A1(n16511), .A2(N12019), .ZN(N31061));
    NANDX1 U18190 (.A1(N9113), .A2(n13874), .ZN(N31062));
    INVX1 U18191 (.I(n20147), .ZN(n31063));
    INVX1 U18192 (.I(N10663), .ZN(N31064));
    NANDX1 U18193 (.A1(n17426), .A2(n20535), .ZN(N31065));
    NOR2X1 U18194 (.A1(N6366), .A2(n24423), .ZN(n31066));
    INVX1 U18195 (.I(n18308), .ZN(n31067));
    INVX1 U18196 (.I(N1889), .ZN(N31068));
    NOR2X1 U18197 (.A1(n22412), .A2(N3376), .ZN(N31069));
    NOR2X1 U18198 (.A1(N10326), .A2(n27533), .ZN(n31070));
    NOR2X1 U18199 (.A1(N12278), .A2(n19285), .ZN(N31071));
    INVX1 U18200 (.I(n29683), .ZN(N31072));
    NOR2X1 U18201 (.A1(n13537), .A2(N11564), .ZN(n31073));
    NANDX1 U18202 (.A1(N11211), .A2(n13998), .ZN(n31074));
    NOR2X1 U18203 (.A1(N1220), .A2(n20857), .ZN(n31075));
    NOR2X1 U18204 (.A1(n14157), .A2(n26843), .ZN(n31076));
    INVX1 U18205 (.I(n13694), .ZN(N31077));
    NANDX1 U18206 (.A1(n24849), .A2(N1281), .ZN(N31078));
    INVX1 U18207 (.I(N567), .ZN(n31079));
    INVX1 U18208 (.I(N10865), .ZN(N31080));
    NOR2X1 U18209 (.A1(n25242), .A2(N9597), .ZN(N31081));
    INVX1 U18210 (.I(n22637), .ZN(N31082));
    NOR2X1 U18211 (.A1(N4004), .A2(N346), .ZN(N31083));
    INVX1 U18212 (.I(N3549), .ZN(n31084));
    NOR2X1 U18213 (.A1(n27785), .A2(N3673), .ZN(N31085));
    INVX1 U18214 (.I(N8858), .ZN(n31086));
    NOR2X1 U18215 (.A1(N2419), .A2(N10077), .ZN(n31087));
    NANDX1 U18216 (.A1(n23887), .A2(N12794), .ZN(N31088));
    NANDX1 U18217 (.A1(N5615), .A2(n26488), .ZN(N31089));
    INVX1 U18218 (.I(N326), .ZN(n31090));
    NOR2X1 U18219 (.A1(n25363), .A2(n19590), .ZN(n31091));
    NOR2X1 U18220 (.A1(n24789), .A2(N991), .ZN(n31092));
    NANDX1 U18221 (.A1(N4248), .A2(N11415), .ZN(N31093));
    NANDX1 U18222 (.A1(N10031), .A2(n15418), .ZN(N31094));
    NANDX1 U18223 (.A1(n24278), .A2(N7527), .ZN(n31095));
    NANDX1 U18224 (.A1(N10486), .A2(n29897), .ZN(N31096));
    NOR2X1 U18225 (.A1(N7904), .A2(N5990), .ZN(N31097));
    INVX1 U18226 (.I(N6541), .ZN(N31098));
    NANDX1 U18227 (.A1(N2188), .A2(n19335), .ZN(n31099));
    INVX1 U18228 (.I(n26501), .ZN(n31100));
    NANDX1 U18229 (.A1(N579), .A2(n15387), .ZN(N31101));
    INVX1 U18230 (.I(n25942), .ZN(n31102));
    NOR2X1 U18231 (.A1(N9933), .A2(n20593), .ZN(N31103));
    INVX1 U18232 (.I(n13094), .ZN(n31104));
    INVX1 U18233 (.I(N5806), .ZN(N31105));
    INVX1 U18234 (.I(n23431), .ZN(n31106));
    INVX1 U18235 (.I(N4761), .ZN(N31107));
    NANDX1 U18236 (.A1(n17311), .A2(N470), .ZN(N31108));
    NOR2X1 U18237 (.A1(N5631), .A2(N6490), .ZN(n31109));
    NOR2X1 U18238 (.A1(N11621), .A2(N3489), .ZN(N31110));
    NANDX1 U18239 (.A1(N3121), .A2(N5676), .ZN(N31111));
    NOR2X1 U18240 (.A1(N6974), .A2(n20737), .ZN(N31112));
    INVX1 U18241 (.I(n26250), .ZN(N31113));
    INVX1 U18242 (.I(N3501), .ZN(n31114));
    NANDX1 U18243 (.A1(n29524), .A2(N1994), .ZN(N31115));
    INVX1 U18244 (.I(n23914), .ZN(N31116));
    NOR2X1 U18245 (.A1(N3032), .A2(n29719), .ZN(N31117));
    INVX1 U18246 (.I(n26462), .ZN(N31118));
    INVX1 U18247 (.I(n17164), .ZN(n31119));
    NOR2X1 U18248 (.A1(n15237), .A2(N6194), .ZN(n31120));
    NOR2X1 U18249 (.A1(N9428), .A2(N1244), .ZN(n31121));
    NOR2X1 U18250 (.A1(N9609), .A2(N4732), .ZN(n31122));
    NANDX1 U18251 (.A1(N12729), .A2(n29106), .ZN(N31123));
    NANDX1 U18252 (.A1(N8263), .A2(n19705), .ZN(n31124));
    NANDX1 U18253 (.A1(N4376), .A2(n14252), .ZN(N31125));
    INVX1 U18254 (.I(n14990), .ZN(n31126));
    NOR2X1 U18255 (.A1(n26142), .A2(N4621), .ZN(N31127));
    INVX1 U18256 (.I(n29790), .ZN(N31128));
    NANDX1 U18257 (.A1(n25694), .A2(N617), .ZN(N31129));
    NOR2X1 U18258 (.A1(n23620), .A2(n17780), .ZN(n31130));
    NOR2X1 U18259 (.A1(n27417), .A2(N12534), .ZN(N31131));
    NOR2X1 U18260 (.A1(N6708), .A2(n13778), .ZN(n31132));
    NANDX1 U18261 (.A1(n16316), .A2(n18509), .ZN(N31133));
    NOR2X1 U18262 (.A1(n17606), .A2(N6038), .ZN(N31134));
    NANDX1 U18263 (.A1(n25868), .A2(n25743), .ZN(n31135));
    INVX1 U18264 (.I(n18804), .ZN(n31136));
    NANDX1 U18265 (.A1(N2775), .A2(N3657), .ZN(N31137));
    NANDX1 U18266 (.A1(n28916), .A2(n26975), .ZN(N31138));
    NOR2X1 U18267 (.A1(n17130), .A2(n23187), .ZN(n31139));
    INVX1 U18268 (.I(n17746), .ZN(n31140));
    INVX1 U18269 (.I(n15768), .ZN(N31141));
    NOR2X1 U18270 (.A1(n17975), .A2(n13047), .ZN(n31142));
    INVX1 U18271 (.I(n27862), .ZN(n31143));
    NANDX1 U18272 (.A1(n20259), .A2(n16890), .ZN(n31144));
    INVX1 U18273 (.I(n27329), .ZN(N31145));
    NANDX1 U18274 (.A1(n19358), .A2(N3229), .ZN(n31146));
    INVX1 U18275 (.I(n15088), .ZN(n31147));
    NOR2X1 U18276 (.A1(n24438), .A2(n22453), .ZN(N31148));
    NANDX1 U18277 (.A1(n15773), .A2(n14670), .ZN(N31149));
    INVX1 U18278 (.I(N3113), .ZN(n31150));
    INVX1 U18279 (.I(n24596), .ZN(n31151));
    NOR2X1 U18280 (.A1(N4556), .A2(n16743), .ZN(N31152));
    NOR2X1 U18281 (.A1(N8839), .A2(n21071), .ZN(N31153));
    NANDX1 U18282 (.A1(n26814), .A2(n22679), .ZN(n31154));
    NOR2X1 U18283 (.A1(n13099), .A2(n19554), .ZN(N31155));
    NOR2X1 U18284 (.A1(n29989), .A2(N2608), .ZN(n31156));
    NANDX1 U18285 (.A1(n15972), .A2(n21965), .ZN(N31157));
    NOR2X1 U18286 (.A1(n20207), .A2(n25614), .ZN(N31158));
    NOR2X1 U18287 (.A1(N3069), .A2(n17929), .ZN(N31159));
    NANDX1 U18288 (.A1(n18841), .A2(N2461), .ZN(N31160));
    NANDX1 U18289 (.A1(n21953), .A2(N2528), .ZN(n31161));
    NANDX1 U18290 (.A1(N618), .A2(N7083), .ZN(n31162));
    NANDX1 U18291 (.A1(n27165), .A2(n15921), .ZN(N31163));
    NANDX1 U18292 (.A1(N6084), .A2(N1158), .ZN(N31164));
    INVX1 U18293 (.I(N10183), .ZN(N31165));
    NOR2X1 U18294 (.A1(n20417), .A2(N4403), .ZN(N31166));
    NOR2X1 U18295 (.A1(n23025), .A2(n14512), .ZN(N31167));
    INVX1 U18296 (.I(N3413), .ZN(n31168));
    NOR2X1 U18297 (.A1(n27407), .A2(n29026), .ZN(N31169));
    NOR2X1 U18298 (.A1(N338), .A2(N5378), .ZN(n31170));
    INVX1 U18299 (.I(N7740), .ZN(N31171));
    INVX1 U18300 (.I(n17133), .ZN(N31172));
    NOR2X1 U18301 (.A1(n29063), .A2(N10520), .ZN(n31173));
    NANDX1 U18302 (.A1(N6008), .A2(n27909), .ZN(N31174));
    NOR2X1 U18303 (.A1(N10490), .A2(n17533), .ZN(n31175));
    INVX1 U18304 (.I(N11647), .ZN(N31176));
    NOR2X1 U18305 (.A1(N9286), .A2(n14464), .ZN(n31177));
    NOR2X1 U18306 (.A1(N2249), .A2(n17132), .ZN(N31178));
    NANDX1 U18307 (.A1(N5321), .A2(n24332), .ZN(n31179));
    NANDX1 U18308 (.A1(N10291), .A2(n21602), .ZN(N31180));
    INVX1 U18309 (.I(N4555), .ZN(n31181));
    NOR2X1 U18310 (.A1(n16500), .A2(N11319), .ZN(N31182));
    NOR2X1 U18311 (.A1(n12898), .A2(n17013), .ZN(n31183));
    INVX1 U18312 (.I(N11824), .ZN(N31184));
    INVX1 U18313 (.I(N2347), .ZN(N31185));
    NOR2X1 U18314 (.A1(n25303), .A2(N6805), .ZN(N31186));
    NANDX1 U18315 (.A1(N1259), .A2(n24606), .ZN(n31187));
    NANDX1 U18316 (.A1(N8215), .A2(n22452), .ZN(N31188));
    NANDX1 U18317 (.A1(n24149), .A2(n24700), .ZN(N31189));
    INVX1 U18318 (.I(N2832), .ZN(n31190));
    NOR2X1 U18319 (.A1(n20000), .A2(n15065), .ZN(n31191));
    NANDX1 U18320 (.A1(N11464), .A2(n14748), .ZN(N31192));
    NOR2X1 U18321 (.A1(N10525), .A2(n19808), .ZN(N31193));
    NOR2X1 U18322 (.A1(n17324), .A2(n21266), .ZN(N31194));
    NOR2X1 U18323 (.A1(N12239), .A2(n21650), .ZN(n31195));
    NANDX1 U18324 (.A1(n14585), .A2(n28042), .ZN(N31196));
    NOR2X1 U18325 (.A1(N9951), .A2(N3346), .ZN(N31197));
    NOR2X1 U18326 (.A1(N4419), .A2(N8995), .ZN(n31198));
    NANDX1 U18327 (.A1(n26871), .A2(n17669), .ZN(N31199));
    NANDX1 U18328 (.A1(N9994), .A2(n13337), .ZN(N31200));
    NOR2X1 U18329 (.A1(n28575), .A2(N3199), .ZN(n31201));
    NANDX1 U18330 (.A1(n27309), .A2(N3224), .ZN(N31202));
    NOR2X1 U18331 (.A1(n19158), .A2(n13748), .ZN(N31203));
    NOR2X1 U18332 (.A1(n22325), .A2(N934), .ZN(N31204));
    NOR2X1 U18333 (.A1(N12368), .A2(n13173), .ZN(N31205));
    INVX1 U18334 (.I(N7064), .ZN(N31206));
    INVX1 U18335 (.I(n17981), .ZN(N31207));
    NANDX1 U18336 (.A1(n26268), .A2(N9888), .ZN(n31208));
    NANDX1 U18337 (.A1(N550), .A2(N7443), .ZN(n31209));
    NANDX1 U18338 (.A1(n15981), .A2(n25111), .ZN(N31210));
    NOR2X1 U18339 (.A1(n14535), .A2(N8310), .ZN(N31211));
    NOR2X1 U18340 (.A1(n12972), .A2(N70), .ZN(N31212));
    NOR2X1 U18341 (.A1(n28841), .A2(N3293), .ZN(N31213));
    NANDX1 U18342 (.A1(n17861), .A2(n17040), .ZN(n31214));
    NOR2X1 U18343 (.A1(n28747), .A2(N6534), .ZN(n31215));
    NANDX1 U18344 (.A1(n29675), .A2(n19706), .ZN(n31216));
    NOR2X1 U18345 (.A1(N6601), .A2(N5887), .ZN(n31217));
    NOR2X1 U18346 (.A1(N3525), .A2(N2017), .ZN(N31218));
    INVX1 U18347 (.I(N10268), .ZN(N31219));
    NANDX1 U18348 (.A1(n24207), .A2(n23604), .ZN(N31220));
    INVX1 U18349 (.I(N7742), .ZN(N31221));
    INVX1 U18350 (.I(n21642), .ZN(n31222));
    INVX1 U18351 (.I(N1906), .ZN(N31223));
    NOR2X1 U18352 (.A1(N4681), .A2(N3466), .ZN(N31224));
    NOR2X1 U18353 (.A1(N7973), .A2(n15395), .ZN(N31225));
    INVX1 U18354 (.I(n13573), .ZN(n31226));
    INVX1 U18355 (.I(n26908), .ZN(N31227));
    NANDX1 U18356 (.A1(n14882), .A2(n26445), .ZN(n31228));
    NANDX1 U18357 (.A1(n15218), .A2(n21606), .ZN(N31229));
    NOR2X1 U18358 (.A1(n22095), .A2(n25131), .ZN(N31230));
    NOR2X1 U18359 (.A1(N8722), .A2(n23959), .ZN(N31231));
    INVX1 U18360 (.I(n21489), .ZN(N31232));
    INVX1 U18361 (.I(N11631), .ZN(N31233));
    NOR2X1 U18362 (.A1(n13392), .A2(N3135), .ZN(n31234));
    NANDX1 U18363 (.A1(N3858), .A2(n14869), .ZN(N31235));
    NOR2X1 U18364 (.A1(N7323), .A2(N6609), .ZN(N31236));
    NANDX1 U18365 (.A1(N11279), .A2(n23469), .ZN(n31237));
    NANDX1 U18366 (.A1(n15764), .A2(n20239), .ZN(n31238));
    NOR2X1 U18367 (.A1(N509), .A2(N5108), .ZN(n31239));
    NANDX1 U18368 (.A1(N4287), .A2(n26713), .ZN(N31240));
    NANDX1 U18369 (.A1(n14942), .A2(N10267), .ZN(N31241));
    INVX1 U18370 (.I(N12224), .ZN(n31242));
    NANDX1 U18371 (.A1(n28738), .A2(N3575), .ZN(N31243));
    NOR2X1 U18372 (.A1(N10231), .A2(N2668), .ZN(n31244));
    NANDX1 U18373 (.A1(N1926), .A2(N6372), .ZN(n31245));
    NOR2X1 U18374 (.A1(N5355), .A2(N3317), .ZN(N31246));
    INVX1 U18375 (.I(N525), .ZN(n31247));
    NOR2X1 U18376 (.A1(n23045), .A2(n23993), .ZN(N31248));
    NANDX1 U18377 (.A1(N8671), .A2(n14094), .ZN(n31249));
    INVX1 U18378 (.I(n27877), .ZN(n31250));
    NANDX1 U18379 (.A1(N304), .A2(n20724), .ZN(N31251));
    NOR2X1 U18380 (.A1(n29819), .A2(N5528), .ZN(N31252));
    INVX1 U18381 (.I(N12456), .ZN(N31253));
    NOR2X1 U18382 (.A1(n18692), .A2(n29754), .ZN(n31254));
    INVX1 U18383 (.I(n28764), .ZN(N31255));
    NANDX1 U18384 (.A1(N12554), .A2(N10652), .ZN(n31256));
    NANDX1 U18385 (.A1(N7486), .A2(n15096), .ZN(n31257));
    NOR2X1 U18386 (.A1(N10802), .A2(n26862), .ZN(N31258));
    INVX1 U18387 (.I(N7598), .ZN(N31259));
    NANDX1 U18388 (.A1(n18765), .A2(N4186), .ZN(N31260));
    INVX1 U18389 (.I(n21419), .ZN(n31261));
    NOR2X1 U18390 (.A1(n26179), .A2(n29181), .ZN(N31262));
    NOR2X1 U18391 (.A1(N5326), .A2(N3381), .ZN(N31263));
    NANDX1 U18392 (.A1(N10854), .A2(N6545), .ZN(n31264));
    NANDX1 U18393 (.A1(n17165), .A2(n13797), .ZN(n31265));
    NANDX1 U18394 (.A1(n27051), .A2(N985), .ZN(N31266));
    NOR2X1 U18395 (.A1(N9467), .A2(N197), .ZN(n31267));
    NANDX1 U18396 (.A1(N5513), .A2(n15292), .ZN(n31268));
    INVX1 U18397 (.I(N4876), .ZN(N31269));
    NOR2X1 U18398 (.A1(n23568), .A2(N12473), .ZN(N31270));
    INVX1 U18399 (.I(N12195), .ZN(N31271));
    INVX1 U18400 (.I(n18647), .ZN(N31272));
    NOR2X1 U18401 (.A1(n14451), .A2(N3249), .ZN(N31273));
    INVX1 U18402 (.I(N12548), .ZN(N31274));
    NANDX1 U18403 (.A1(n24597), .A2(N10326), .ZN(N31275));
    NOR2X1 U18404 (.A1(n19703), .A2(N9121), .ZN(n31276));
    NOR2X1 U18405 (.A1(N3362), .A2(N7532), .ZN(N31277));
    INVX1 U18406 (.I(N4346), .ZN(n31278));
    NANDX1 U18407 (.A1(n20094), .A2(N4543), .ZN(n31279));
    NOR2X1 U18408 (.A1(n14167), .A2(n19834), .ZN(N31280));
    INVX1 U18409 (.I(n19042), .ZN(n31281));
    NANDX1 U18410 (.A1(N848), .A2(n20075), .ZN(N31282));
    NOR2X1 U18411 (.A1(N1603), .A2(n25293), .ZN(N31283));
    NANDX1 U18412 (.A1(N5079), .A2(N9607), .ZN(N31284));
    INVX1 U18413 (.I(n26295), .ZN(N31285));
    NOR2X1 U18414 (.A1(N10949), .A2(N9316), .ZN(N31286));
    NOR2X1 U18415 (.A1(n18936), .A2(n29018), .ZN(N31287));
    INVX1 U18416 (.I(n13951), .ZN(n31288));
    INVX1 U18417 (.I(n14814), .ZN(n31289));
    NOR2X1 U18418 (.A1(n25286), .A2(N7724), .ZN(N31290));
    NOR2X1 U18419 (.A1(n29828), .A2(n16484), .ZN(N31291));
    INVX1 U18420 (.I(N8085), .ZN(n31292));
    NANDX1 U18421 (.A1(n17605), .A2(n28495), .ZN(N31293));
    NANDX1 U18422 (.A1(n26240), .A2(N8976), .ZN(N31294));
    INVX1 U18423 (.I(n21396), .ZN(N31295));
    NOR2X1 U18424 (.A1(n27249), .A2(n19563), .ZN(n31296));
    INVX1 U18425 (.I(n23407), .ZN(N31297));
    NOR2X1 U18426 (.A1(n28684), .A2(n21283), .ZN(n31298));
    NANDX1 U18427 (.A1(N6043), .A2(n20163), .ZN(N31299));
    NOR2X1 U18428 (.A1(n19994), .A2(N10965), .ZN(n31300));
    NANDX1 U18429 (.A1(n14434), .A2(N6113), .ZN(N31301));
    NOR2X1 U18430 (.A1(n17528), .A2(N5803), .ZN(n31302));
    INVX1 U18431 (.I(n16090), .ZN(n31303));
    NOR2X1 U18432 (.A1(N8230), .A2(n22255), .ZN(n31304));
    INVX1 U18433 (.I(N10100), .ZN(n31305));
    INVX1 U18434 (.I(n17040), .ZN(n31306));
    NANDX1 U18435 (.A1(n28314), .A2(n13703), .ZN(n31307));
    NANDX1 U18436 (.A1(n17739), .A2(N1301), .ZN(N31308));
    INVX1 U18437 (.I(N6439), .ZN(N31309));
    INVX1 U18438 (.I(N2357), .ZN(N31310));
    NANDX1 U18439 (.A1(n24587), .A2(n22519), .ZN(n31311));
    NANDX1 U18440 (.A1(N3004), .A2(n22045), .ZN(N31312));
    INVX1 U18441 (.I(N5998), .ZN(N31313));
    NOR2X1 U18442 (.A1(n18366), .A2(n23525), .ZN(n31314));
    NOR2X1 U18443 (.A1(N2695), .A2(N9478), .ZN(N31315));
    NANDX1 U18444 (.A1(N10924), .A2(n20293), .ZN(n31316));
    NOR2X1 U18445 (.A1(N9585), .A2(N8513), .ZN(N31317));
    NANDX1 U18446 (.A1(N11718), .A2(N6689), .ZN(n31318));
    NOR2X1 U18447 (.A1(n29660), .A2(n12988), .ZN(N31319));
    NOR2X1 U18448 (.A1(N10735), .A2(n19427), .ZN(N31320));
    NOR2X1 U18449 (.A1(n13091), .A2(N5469), .ZN(N31321));
    INVX1 U18450 (.I(n24171), .ZN(n31322));
    NOR2X1 U18451 (.A1(n28057), .A2(n16078), .ZN(n31323));
    INVX1 U18452 (.I(n22615), .ZN(N31324));
    NOR2X1 U18453 (.A1(n24402), .A2(n16003), .ZN(N31325));
    NANDX1 U18454 (.A1(n27096), .A2(n14041), .ZN(N31326));
    INVX1 U18455 (.I(n26581), .ZN(n31327));
    NANDX1 U18456 (.A1(N11466), .A2(n24726), .ZN(N31328));
    NOR2X1 U18457 (.A1(N1264), .A2(n25004), .ZN(N31329));
    NOR2X1 U18458 (.A1(n23462), .A2(n24526), .ZN(n31330));
    NOR2X1 U18459 (.A1(N5384), .A2(N5123), .ZN(n31331));
    NOR2X1 U18460 (.A1(n17289), .A2(N6775), .ZN(N31332));
    NANDX1 U18461 (.A1(N765), .A2(N808), .ZN(N31333));
    NANDX1 U18462 (.A1(n28821), .A2(N5446), .ZN(n31334));
    NOR2X1 U18463 (.A1(n21299), .A2(N8103), .ZN(N31335));
    NANDX1 U18464 (.A1(n25862), .A2(N3144), .ZN(N31336));
    NOR2X1 U18465 (.A1(N9765), .A2(N274), .ZN(N31337));
    NOR2X1 U18466 (.A1(N2521), .A2(N11739), .ZN(N31338));
    NANDX1 U18467 (.A1(N3790), .A2(N1563), .ZN(N31339));
    NANDX1 U18468 (.A1(N309), .A2(n13585), .ZN(N31340));
    NANDX1 U18469 (.A1(n28513), .A2(n18968), .ZN(N31341));
    NOR2X1 U18470 (.A1(n15869), .A2(n24817), .ZN(N31342));
    INVX1 U18471 (.I(n27391), .ZN(N31343));
    NANDX1 U18472 (.A1(n13383), .A2(n17308), .ZN(n31344));
    NANDX1 U18473 (.A1(N7389), .A2(n13262), .ZN(n31345));
    NANDX1 U18474 (.A1(n15491), .A2(n22179), .ZN(N31346));
    NANDX1 U18475 (.A1(N7195), .A2(n16615), .ZN(n31347));
    INVX1 U18476 (.I(N7469), .ZN(n31348));
    NANDX1 U18477 (.A1(N7816), .A2(N7768), .ZN(n31349));
    NOR2X1 U18478 (.A1(N166), .A2(n28029), .ZN(N31350));
    NANDX1 U18479 (.A1(N474), .A2(N37), .ZN(n31351));
    INVX1 U18480 (.I(n28986), .ZN(N31352));
    INVX1 U18481 (.I(N9910), .ZN(n31353));
    NANDX1 U18482 (.A1(n20943), .A2(n22485), .ZN(n31354));
    NANDX1 U18483 (.A1(n16387), .A2(n24428), .ZN(N31355));
    INVX1 U18484 (.I(n17774), .ZN(N31356));
    NOR2X1 U18485 (.A1(n26920), .A2(n29019), .ZN(N31357));
    INVX1 U18486 (.I(N7522), .ZN(n31358));
    NOR2X1 U18487 (.A1(n24364), .A2(n24136), .ZN(n31359));
    NOR2X1 U18488 (.A1(n20393), .A2(N1492), .ZN(n31360));
    INVX1 U18489 (.I(n16722), .ZN(N31361));
    INVX1 U18490 (.I(N7688), .ZN(N31362));
    NOR2X1 U18491 (.A1(n23839), .A2(N8161), .ZN(n31363));
    NOR2X1 U18492 (.A1(n16509), .A2(n25708), .ZN(N31364));
    INVX1 U18493 (.I(n26418), .ZN(N31365));
    INVX1 U18494 (.I(N1581), .ZN(n31366));
    NOR2X1 U18495 (.A1(N6638), .A2(N6528), .ZN(N31367));
    INVX1 U18496 (.I(n20296), .ZN(N31368));
    NANDX1 U18497 (.A1(n14735), .A2(n17078), .ZN(n31369));
    NOR2X1 U18498 (.A1(n20465), .A2(n24600), .ZN(N31370));
    NOR2X1 U18499 (.A1(N3252), .A2(n18598), .ZN(N31371));
    NANDX1 U18500 (.A1(n23645), .A2(N8651), .ZN(N31372));
    INVX1 U18501 (.I(n28927), .ZN(n31373));
    NOR2X1 U18502 (.A1(n13812), .A2(n13402), .ZN(N31374));
    INVX1 U18503 (.I(N10533), .ZN(N31375));
    NANDX1 U18504 (.A1(n20571), .A2(n24801), .ZN(N31376));
    NOR2X1 U18505 (.A1(n16851), .A2(N12210), .ZN(N31377));
    INVX1 U18506 (.I(n24177), .ZN(N31378));
    NANDX1 U18507 (.A1(N5356), .A2(n25794), .ZN(N31379));
    NANDX1 U18508 (.A1(n18218), .A2(N10391), .ZN(n31380));
    NANDX1 U18509 (.A1(n29961), .A2(n19416), .ZN(n31381));
    NOR2X1 U18510 (.A1(n17418), .A2(n22667), .ZN(N31382));
    NANDX1 U18511 (.A1(N4581), .A2(N4735), .ZN(N31383));
    INVX1 U18512 (.I(n29403), .ZN(n31384));
    NOR2X1 U18513 (.A1(N5137), .A2(n13077), .ZN(N31385));
    INVX1 U18514 (.I(N9199), .ZN(N31386));
    NOR2X1 U18515 (.A1(n22097), .A2(n18330), .ZN(N31387));
    NOR2X1 U18516 (.A1(N7906), .A2(n23742), .ZN(N31388));
    INVX1 U18517 (.I(n25432), .ZN(N31389));
    INVX1 U18518 (.I(n26450), .ZN(N31390));
    NOR2X1 U18519 (.A1(N1998), .A2(n24015), .ZN(N31391));
    NOR2X1 U18520 (.A1(N949), .A2(n27219), .ZN(N31392));
    INVX1 U18521 (.I(n20364), .ZN(N31393));
    NOR2X1 U18522 (.A1(N1790), .A2(n12894), .ZN(n31394));
    INVX1 U18523 (.I(N6371), .ZN(N31395));
    NOR2X1 U18524 (.A1(n24484), .A2(N5636), .ZN(N31396));
    NOR2X1 U18525 (.A1(n29621), .A2(N7274), .ZN(N31397));
    INVX1 U18526 (.I(n27380), .ZN(N31398));
    NANDX1 U18527 (.A1(n18596), .A2(n15573), .ZN(n31399));
    NANDX1 U18528 (.A1(n15062), .A2(n27875), .ZN(n31400));
    NOR2X1 U18529 (.A1(N10356), .A2(N4079), .ZN(N31401));
    NANDX1 U18530 (.A1(n29704), .A2(N6077), .ZN(N31402));
    NOR2X1 U18531 (.A1(n25692), .A2(N7025), .ZN(N31403));
    NANDX1 U18532 (.A1(n21504), .A2(n27389), .ZN(N31404));
    NANDX1 U18533 (.A1(n23293), .A2(n28843), .ZN(N31405));
    NOR2X1 U18534 (.A1(n18224), .A2(n16333), .ZN(N31406));
    INVX1 U18535 (.I(n23860), .ZN(N31407));
    INVX1 U18536 (.I(N5118), .ZN(N31408));
    NOR2X1 U18537 (.A1(n22545), .A2(N2361), .ZN(N31409));
    NANDX1 U18538 (.A1(n29701), .A2(N6494), .ZN(n31410));
    NOR2X1 U18539 (.A1(n14626), .A2(N4231), .ZN(n31411));
    NOR2X1 U18540 (.A1(n24981), .A2(n27007), .ZN(N31412));
    NANDX1 U18541 (.A1(n13108), .A2(N2946), .ZN(n31413));
    NANDX1 U18542 (.A1(N8663), .A2(n28669), .ZN(N31414));
    INVX1 U18543 (.I(n18727), .ZN(N31415));
    INVX1 U18544 (.I(N11760), .ZN(N31416));
    NANDX1 U18545 (.A1(n13186), .A2(n23048), .ZN(N31417));
    INVX1 U18546 (.I(n18079), .ZN(N31418));
    INVX1 U18547 (.I(N12389), .ZN(n31419));
    INVX1 U18548 (.I(N3663), .ZN(N31420));
    NOR2X1 U18549 (.A1(N6394), .A2(n24721), .ZN(N31421));
    INVX1 U18550 (.I(n24655), .ZN(N31422));
    NANDX1 U18551 (.A1(n19161), .A2(N9143), .ZN(n31423));
    NOR2X1 U18552 (.A1(n23863), .A2(n22685), .ZN(N31424));
    NOR2X1 U18553 (.A1(N5742), .A2(n24353), .ZN(N31425));
    NOR2X1 U18554 (.A1(n18950), .A2(N2878), .ZN(n31426));
    INVX1 U18555 (.I(N7553), .ZN(n31427));
    NANDX1 U18556 (.A1(n25392), .A2(n19312), .ZN(N31428));
    INVX1 U18557 (.I(n27138), .ZN(n31429));
    NOR2X1 U18558 (.A1(N10576), .A2(n15080), .ZN(N31430));
    NOR2X1 U18559 (.A1(N11525), .A2(n29066), .ZN(N31431));
    NOR2X1 U18560 (.A1(n20728), .A2(n24020), .ZN(N31432));
    NOR2X1 U18561 (.A1(N8793), .A2(n18537), .ZN(N31433));
    NANDX1 U18562 (.A1(n16514), .A2(n16241), .ZN(N31434));
    NOR2X1 U18563 (.A1(N10239), .A2(n27486), .ZN(n31435));
    NOR2X1 U18564 (.A1(n15980), .A2(n21701), .ZN(n31436));
    NANDX1 U18565 (.A1(n23490), .A2(n13140), .ZN(n31437));
    INVX1 U18566 (.I(N905), .ZN(N31438));
    INVX1 U18567 (.I(N4881), .ZN(N31439));
    INVX1 U18568 (.I(N3774), .ZN(n31440));
    NANDX1 U18569 (.A1(N9561), .A2(N2910), .ZN(N31441));
    INVX1 U18570 (.I(N8889), .ZN(n31442));
    INVX1 U18571 (.I(N4450), .ZN(N31443));
    NANDX1 U18572 (.A1(n23722), .A2(n28469), .ZN(n31444));
    INVX1 U18573 (.I(n21075), .ZN(n31445));
    NANDX1 U18574 (.A1(N3924), .A2(N7452), .ZN(n31446));
    NANDX1 U18575 (.A1(N3701), .A2(n17690), .ZN(N31447));
    NANDX1 U18576 (.A1(n12913), .A2(n22231), .ZN(N31448));
    INVX1 U18577 (.I(n23066), .ZN(n31449));
    NANDX1 U18578 (.A1(N842), .A2(n13994), .ZN(N31450));
    NOR2X1 U18579 (.A1(n24145), .A2(N7436), .ZN(N31451));
    INVX1 U18580 (.I(n27919), .ZN(N31452));
    NANDX1 U18581 (.A1(N11947), .A2(n19389), .ZN(N31453));
    NOR2X1 U18582 (.A1(N9396), .A2(n22384), .ZN(n31454));
    INVX1 U18583 (.I(N9835), .ZN(n31455));
    INVX1 U18584 (.I(N6179), .ZN(n31456));
    NANDX1 U18585 (.A1(n25604), .A2(N168), .ZN(n31457));
    NANDX1 U18586 (.A1(N2918), .A2(N10398), .ZN(n31458));
    INVX1 U18587 (.I(N9168), .ZN(N31459));
    NANDX1 U18588 (.A1(N5506), .A2(n19959), .ZN(n31460));
    NOR2X1 U18589 (.A1(n28571), .A2(N5405), .ZN(n31461));
    NOR2X1 U18590 (.A1(N12428), .A2(n29151), .ZN(n31462));
    INVX1 U18591 (.I(n19863), .ZN(N31463));
    NOR2X1 U18592 (.A1(n17005), .A2(n17740), .ZN(N31464));
    NOR2X1 U18593 (.A1(N6256), .A2(n21138), .ZN(N31465));
    INVX1 U18594 (.I(n17200), .ZN(N31466));
    NOR2X1 U18595 (.A1(n21136), .A2(N3031), .ZN(N31467));
    NANDX1 U18596 (.A1(N6106), .A2(n17195), .ZN(n31468));
    NANDX1 U18597 (.A1(N6438), .A2(n20112), .ZN(N31469));
    NANDX1 U18598 (.A1(n29168), .A2(n17840), .ZN(n31470));
    NANDX1 U18599 (.A1(N4536), .A2(N7662), .ZN(N31471));
    INVX1 U18600 (.I(N2970), .ZN(N31472));
    INVX1 U18601 (.I(n22881), .ZN(N31473));
    INVX1 U18602 (.I(N640), .ZN(N31474));
    NANDX1 U18603 (.A1(N12381), .A2(n20737), .ZN(N31475));
    NANDX1 U18604 (.A1(n18681), .A2(n22643), .ZN(n31476));
    NANDX1 U18605 (.A1(N9681), .A2(N3807), .ZN(N31477));
    NOR2X1 U18606 (.A1(n27226), .A2(n13503), .ZN(N31478));
    NANDX1 U18607 (.A1(N9373), .A2(N8170), .ZN(N31479));
    INVX1 U18608 (.I(N3126), .ZN(n31480));
    INVX1 U18609 (.I(n28307), .ZN(N31481));
    INVX1 U18610 (.I(N2199), .ZN(N31482));
    INVX1 U18611 (.I(N6524), .ZN(N31483));
    NANDX1 U18612 (.A1(N12231), .A2(n22886), .ZN(N31484));
    NANDX1 U18613 (.A1(N2418), .A2(n15629), .ZN(N31485));
    NOR2X1 U18614 (.A1(n21755), .A2(n16156), .ZN(n31486));
    NANDX1 U18615 (.A1(N12354), .A2(N3550), .ZN(n31487));
    NOR2X1 U18616 (.A1(n23557), .A2(n27337), .ZN(N31488));
    INVX1 U18617 (.I(n15924), .ZN(N31489));
    NANDX1 U18618 (.A1(n24430), .A2(n17988), .ZN(N31490));
    INVX1 U18619 (.I(N3665), .ZN(N31491));
    NOR2X1 U18620 (.A1(n25943), .A2(N6791), .ZN(N31492));
    INVX1 U18621 (.I(N12673), .ZN(n31493));
    NOR2X1 U18622 (.A1(N1385), .A2(n17242), .ZN(n31494));
    INVX1 U18623 (.I(n26817), .ZN(N31495));
    NANDX1 U18624 (.A1(N9158), .A2(n13641), .ZN(N31496));
    INVX1 U18625 (.I(n24787), .ZN(N31497));
    NANDX1 U18626 (.A1(N630), .A2(n29503), .ZN(N31498));
    NOR2X1 U18627 (.A1(N1544), .A2(N2916), .ZN(N31499));
    INVX1 U18628 (.I(n25101), .ZN(n31500));
    NANDX1 U18629 (.A1(N3752), .A2(N10887), .ZN(N31501));
    NOR2X1 U18630 (.A1(n28182), .A2(n17435), .ZN(N31502));
    INVX1 U18631 (.I(N1709), .ZN(n31503));
    NOR2X1 U18632 (.A1(n17535), .A2(n27197), .ZN(n31504));
    INVX1 U18633 (.I(n18768), .ZN(N31505));
    INVX1 U18634 (.I(n14025), .ZN(N31506));
    INVX1 U18635 (.I(N4657), .ZN(N31507));
    NOR2X1 U18636 (.A1(N12466), .A2(n13815), .ZN(N31508));
    NANDX1 U18637 (.A1(n21478), .A2(n27162), .ZN(n31509));
    NOR2X1 U18638 (.A1(N10668), .A2(n26527), .ZN(n31510));
    NOR2X1 U18639 (.A1(N12211), .A2(n29442), .ZN(N31511));
    NOR2X1 U18640 (.A1(n25872), .A2(n18117), .ZN(N31512));
    NANDX1 U18641 (.A1(n25320), .A2(n22099), .ZN(N31513));
    INVX1 U18642 (.I(N12617), .ZN(N31514));
    INVX1 U18643 (.I(N7904), .ZN(n31515));
    NANDX1 U18644 (.A1(n19786), .A2(n23662), .ZN(N31516));
    NANDX1 U18645 (.A1(N8416), .A2(N470), .ZN(N31517));
    NANDX1 U18646 (.A1(N2849), .A2(N5127), .ZN(N31518));
    NOR2X1 U18647 (.A1(N3875), .A2(N7502), .ZN(N31519));
    INVX1 U18648 (.I(n25352), .ZN(N31520));
    INVX1 U18649 (.I(n17778), .ZN(N31521));
    NANDX1 U18650 (.A1(n19613), .A2(n19810), .ZN(N31522));
    INVX1 U18651 (.I(N7479), .ZN(n31523));
    NOR2X1 U18652 (.A1(N2388), .A2(n14156), .ZN(N31524));
    NANDX1 U18653 (.A1(n27707), .A2(n24816), .ZN(N31525));
    NOR2X1 U18654 (.A1(N10187), .A2(n27067), .ZN(n31526));
    NOR2X1 U18655 (.A1(N6120), .A2(N5277), .ZN(N31527));
    INVX1 U18656 (.I(N3254), .ZN(N31528));
    INVX1 U18657 (.I(n21755), .ZN(N31529));
    INVX1 U18658 (.I(n23799), .ZN(n31530));
    INVX1 U18659 (.I(N1957), .ZN(n31531));
    NANDX1 U18660 (.A1(N11504), .A2(n13846), .ZN(N31532));
    NOR2X1 U18661 (.A1(N4590), .A2(N1486), .ZN(N31533));
    NOR2X1 U18662 (.A1(N12763), .A2(N9857), .ZN(n31534));
    NOR2X1 U18663 (.A1(n20241), .A2(n15368), .ZN(N31535));
    INVX1 U18664 (.I(n22958), .ZN(N31536));
    NANDX1 U18665 (.A1(N12502), .A2(n17636), .ZN(N31537));
    INVX1 U18666 (.I(n22688), .ZN(N31538));
    NANDX1 U18667 (.A1(N9114), .A2(n17368), .ZN(n31539));
    NANDX1 U18668 (.A1(N262), .A2(N9182), .ZN(N31540));
    INVX1 U18669 (.I(N10577), .ZN(N31541));
    NANDX1 U18670 (.A1(n23014), .A2(n14579), .ZN(N31542));
    NOR2X1 U18671 (.A1(n20550), .A2(n26082), .ZN(N31543));
    NOR2X1 U18672 (.A1(N1862), .A2(N534), .ZN(N31544));
    INVX1 U18673 (.I(n19192), .ZN(n31545));
    NOR2X1 U18674 (.A1(N4981), .A2(N1599), .ZN(N31546));
    INVX1 U18675 (.I(N8909), .ZN(n31547));
    NANDX1 U18676 (.A1(n14918), .A2(n19240), .ZN(N31548));
    NOR2X1 U18677 (.A1(n21114), .A2(N593), .ZN(n31549));
    NANDX1 U18678 (.A1(N12800), .A2(n28404), .ZN(N31550));
    NANDX1 U18679 (.A1(n21202), .A2(n28665), .ZN(N31551));
    NOR2X1 U18680 (.A1(N8978), .A2(n27802), .ZN(n31552));
    NANDX1 U18681 (.A1(N1854), .A2(N12243), .ZN(N31553));
    NANDX1 U18682 (.A1(N10965), .A2(N8187), .ZN(N31554));
    INVX1 U18683 (.I(N12826), .ZN(n31555));
    NANDX1 U18684 (.A1(n28838), .A2(n20578), .ZN(N31556));
    NOR2X1 U18685 (.A1(n22379), .A2(N10737), .ZN(N31557));
    NOR2X1 U18686 (.A1(N1150), .A2(n27266), .ZN(n31558));
    INVX1 U18687 (.I(n20389), .ZN(n31559));
    NOR2X1 U18688 (.A1(N4250), .A2(N9542), .ZN(N31560));
    NANDX1 U18689 (.A1(n17049), .A2(N7809), .ZN(N31561));
    NANDX1 U18690 (.A1(n26811), .A2(N6336), .ZN(N31562));
    INVX1 U18691 (.I(N5651), .ZN(N31563));
    INVX1 U18692 (.I(N5916), .ZN(n31564));
    INVX1 U18693 (.I(N4804), .ZN(N31565));
    INVX1 U18694 (.I(N7030), .ZN(N31566));
    NOR2X1 U18695 (.A1(n19431), .A2(n19855), .ZN(N31567));
    INVX1 U18696 (.I(n18131), .ZN(N31568));
    INVX1 U18697 (.I(n28106), .ZN(n31569));
    NANDX1 U18698 (.A1(n21031), .A2(N7764), .ZN(N31570));
    NANDX1 U18699 (.A1(N6720), .A2(N2339), .ZN(N31571));
    NANDX1 U18700 (.A1(n21440), .A2(n25286), .ZN(n31572));
    INVX1 U18701 (.I(n16165), .ZN(N31573));
    NOR2X1 U18702 (.A1(n26382), .A2(N8261), .ZN(N31574));
    NOR2X1 U18703 (.A1(n21279), .A2(N6909), .ZN(N31575));
    NOR2X1 U18704 (.A1(n13840), .A2(N1386), .ZN(N31576));
    NOR2X1 U18705 (.A1(n18643), .A2(n17239), .ZN(n31577));
    INVX1 U18706 (.I(n20194), .ZN(n31578));
    INVX1 U18707 (.I(n14592), .ZN(N31579));
    NANDX1 U18708 (.A1(N1785), .A2(n13447), .ZN(N31580));
    INVX1 U18709 (.I(N718), .ZN(N31581));
    NANDX1 U18710 (.A1(n13319), .A2(N800), .ZN(N31582));
    NOR2X1 U18711 (.A1(N4218), .A2(N9832), .ZN(N31583));
    NANDX1 U18712 (.A1(n29504), .A2(n28406), .ZN(N31584));
    INVX1 U18713 (.I(N125), .ZN(n31585));
    INVX1 U18714 (.I(N3908), .ZN(N31586));
    NOR2X1 U18715 (.A1(n15791), .A2(n29514), .ZN(N31587));
    NOR2X1 U18716 (.A1(n18191), .A2(N762), .ZN(N31588));
    NANDX1 U18717 (.A1(N6697), .A2(N6562), .ZN(N31589));
    NOR2X1 U18718 (.A1(n15451), .A2(n20352), .ZN(n31590));
    INVX1 U18719 (.I(n23037), .ZN(N31591));
    NANDX1 U18720 (.A1(n29818), .A2(n17153), .ZN(n31592));
    NOR2X1 U18721 (.A1(n22718), .A2(n19032), .ZN(N31593));
    NOR2X1 U18722 (.A1(n22338), .A2(n23249), .ZN(N31594));
    NOR2X1 U18723 (.A1(N1821), .A2(N11176), .ZN(N31595));
    NOR2X1 U18724 (.A1(n27605), .A2(N11300), .ZN(N31596));
    NANDX1 U18725 (.A1(n20073), .A2(n27554), .ZN(N31597));
    INVX1 U18726 (.I(n19449), .ZN(N31598));
    INVX1 U18727 (.I(N3051), .ZN(n31599));
    INVX1 U18728 (.I(n23796), .ZN(N31600));
    INVX1 U18729 (.I(N3894), .ZN(n31601));
    NOR2X1 U18730 (.A1(N2319), .A2(n24245), .ZN(n31602));
    NANDX1 U18731 (.A1(n13917), .A2(N4805), .ZN(N31603));
    NOR2X1 U18732 (.A1(N932), .A2(n16218), .ZN(n31604));
    NANDX1 U18733 (.A1(n19963), .A2(n16992), .ZN(N31605));
    INVX1 U18734 (.I(N1635), .ZN(N31606));
    INVX1 U18735 (.I(n16790), .ZN(n31607));
    NANDX1 U18736 (.A1(N2154), .A2(N2818), .ZN(N31608));
    NOR2X1 U18737 (.A1(N12799), .A2(N11451), .ZN(n31609));
    INVX1 U18738 (.I(n27796), .ZN(N31610));
    NOR2X1 U18739 (.A1(n26839), .A2(N709), .ZN(n31611));
    NOR2X1 U18740 (.A1(n20497), .A2(n17714), .ZN(n31612));
    NANDX1 U18741 (.A1(n15935), .A2(n20032), .ZN(n31613));
    NANDX1 U18742 (.A1(n27745), .A2(N3811), .ZN(N31614));
    NOR2X1 U18743 (.A1(N9099), .A2(N4742), .ZN(N31615));
    NOR2X1 U18744 (.A1(N1731), .A2(n13265), .ZN(n31616));
    INVX1 U18745 (.I(n16700), .ZN(N31617));
    NANDX1 U18746 (.A1(n15949), .A2(n22050), .ZN(N31618));
    NOR2X1 U18747 (.A1(n18102), .A2(n13428), .ZN(N31619));
    NOR2X1 U18748 (.A1(N764), .A2(n24878), .ZN(N31620));
    INVX1 U18749 (.I(n17120), .ZN(N31621));
    INVX1 U18750 (.I(N12851), .ZN(N31622));
    INVX1 U18751 (.I(N855), .ZN(n31623));
    NANDX1 U18752 (.A1(n24102), .A2(n21539), .ZN(N31624));
    INVX1 U18753 (.I(n13996), .ZN(n31625));
    NANDX1 U18754 (.A1(n24011), .A2(n17807), .ZN(n31626));
    NANDX1 U18755 (.A1(n21670), .A2(N11109), .ZN(N31627));
    NANDX1 U18756 (.A1(n23400), .A2(n12935), .ZN(N31628));
    NOR2X1 U18757 (.A1(n28660), .A2(n16395), .ZN(N31629));
    INVX1 U18758 (.I(n20572), .ZN(N31630));
    NANDX1 U18759 (.A1(n23730), .A2(N3862), .ZN(n31631));
    INVX1 U18760 (.I(n13054), .ZN(N31632));
    NOR2X1 U18761 (.A1(N6041), .A2(N36), .ZN(n31633));
    INVX1 U18762 (.I(N7452), .ZN(n31634));
    INVX1 U18763 (.I(N9475), .ZN(n31635));
    NANDX1 U18764 (.A1(N388), .A2(n19575), .ZN(n31636));
    NOR2X1 U18765 (.A1(N2945), .A2(n25768), .ZN(N31637));
    NANDX1 U18766 (.A1(N9312), .A2(N9982), .ZN(N31638));
    NANDX1 U18767 (.A1(N8981), .A2(n18570), .ZN(n31639));
    INVX1 U18768 (.I(n21915), .ZN(n31640));
    NOR2X1 U18769 (.A1(n28771), .A2(n26870), .ZN(n31641));
    INVX1 U18770 (.I(N7766), .ZN(N31642));
    NANDX1 U18771 (.A1(n14729), .A2(N11627), .ZN(N31643));
    NOR2X1 U18772 (.A1(n16344), .A2(n17487), .ZN(n31644));
    INVX1 U18773 (.I(N4940), .ZN(N31645));
    INVX1 U18774 (.I(n17162), .ZN(n31646));
    NANDX1 U18775 (.A1(N5445), .A2(n16383), .ZN(N31647));
    NANDX1 U18776 (.A1(n25019), .A2(N431), .ZN(N31648));
    NOR2X1 U18777 (.A1(N9210), .A2(N8489), .ZN(N31649));
    INVX1 U18778 (.I(N7752), .ZN(n31650));
    NOR2X1 U18779 (.A1(n28807), .A2(n26321), .ZN(N31651));
    NOR2X1 U18780 (.A1(n20584), .A2(n23131), .ZN(N31652));
    NANDX1 U18781 (.A1(N5878), .A2(n14130), .ZN(N31653));
    NANDX1 U18782 (.A1(n23835), .A2(n28859), .ZN(N31654));
    NANDX1 U18783 (.A1(N8806), .A2(N3626), .ZN(N31655));
    NOR2X1 U18784 (.A1(n18516), .A2(N8565), .ZN(N31656));
    NANDX1 U18785 (.A1(N5540), .A2(n19928), .ZN(N31657));
    NOR2X1 U18786 (.A1(N10483), .A2(N8801), .ZN(N31658));
    NANDX1 U18787 (.A1(N10914), .A2(n19315), .ZN(N31659));
    INVX1 U18788 (.I(N7963), .ZN(N31660));
    NOR2X1 U18789 (.A1(n22639), .A2(N4603), .ZN(n31661));
    NOR2X1 U18790 (.A1(N7383), .A2(n20051), .ZN(n31662));
    NANDX1 U18791 (.A1(n19075), .A2(N3996), .ZN(n31663));
    NOR2X1 U18792 (.A1(N3067), .A2(n25842), .ZN(N31664));
    NANDX1 U18793 (.A1(n20486), .A2(n17739), .ZN(N31665));
    INVX1 U18794 (.I(n24111), .ZN(N31666));
    NOR2X1 U18795 (.A1(n20834), .A2(N2539), .ZN(N31667));
    INVX1 U18796 (.I(n14934), .ZN(N31668));
    INVX1 U18797 (.I(N1693), .ZN(n31669));
    NOR2X1 U18798 (.A1(N8388), .A2(N7370), .ZN(N31670));
    INVX1 U18799 (.I(n27703), .ZN(n31671));
    INVX1 U18800 (.I(n14155), .ZN(N31672));
    NANDX1 U18801 (.A1(N3319), .A2(N7318), .ZN(N31673));
    NANDX1 U18802 (.A1(n29399), .A2(n15930), .ZN(N31674));
    INVX1 U18803 (.I(n18336), .ZN(n31675));
    NOR2X1 U18804 (.A1(n23614), .A2(n21403), .ZN(n31676));
    INVX1 U18805 (.I(n28566), .ZN(N31677));
    NANDX1 U18806 (.A1(n21928), .A2(N12186), .ZN(n31678));
    NOR2X1 U18807 (.A1(N7473), .A2(n21581), .ZN(N31679));
    INVX1 U18808 (.I(n28506), .ZN(n31680));
    INVX1 U18809 (.I(n26548), .ZN(N31681));
    INVX1 U18810 (.I(N1656), .ZN(N31682));
    NANDX1 U18811 (.A1(n26129), .A2(n26546), .ZN(n31683));
    NOR2X1 U18812 (.A1(N6809), .A2(n29262), .ZN(N31684));
    INVX1 U18813 (.I(n28825), .ZN(N31685));
    INVX1 U18814 (.I(n23172), .ZN(N31686));
    NANDX1 U18815 (.A1(n22371), .A2(n24091), .ZN(N31687));
    INVX1 U18816 (.I(N719), .ZN(N31688));
    NOR2X1 U18817 (.A1(n26248), .A2(N4909), .ZN(N31689));
    NANDX1 U18818 (.A1(n26560), .A2(n15397), .ZN(n31690));
    NANDX1 U18819 (.A1(n20845), .A2(n22869), .ZN(N31691));
    INVX1 U18820 (.I(N6229), .ZN(N31692));
    INVX1 U18821 (.I(n14561), .ZN(N31693));
    NANDX1 U18822 (.A1(N9860), .A2(N4778), .ZN(N31694));
    INVX1 U18823 (.I(N5851), .ZN(N31695));
    NANDX1 U18824 (.A1(n28498), .A2(N12660), .ZN(N31696));
    INVX1 U18825 (.I(n25990), .ZN(N31697));
    NOR2X1 U18826 (.A1(n25450), .A2(N7585), .ZN(N31698));
    INVX1 U18827 (.I(N6244), .ZN(N31699));
    NOR2X1 U18828 (.A1(n14142), .A2(n25661), .ZN(N31700));
    NANDX1 U18829 (.A1(N10252), .A2(N432), .ZN(N31701));
    INVX1 U18830 (.I(n25372), .ZN(n31702));
    NOR2X1 U18831 (.A1(N6085), .A2(N4640), .ZN(N31703));
    INVX1 U18832 (.I(N2830), .ZN(N31704));
    NANDX1 U18833 (.A1(n18358), .A2(n17390), .ZN(N31705));
    NANDX1 U18834 (.A1(n28217), .A2(N10728), .ZN(N31706));
    NANDX1 U18835 (.A1(N3930), .A2(N11914), .ZN(N31707));
    NOR2X1 U18836 (.A1(n16589), .A2(N784), .ZN(N31708));
    INVX1 U18837 (.I(n16497), .ZN(n31709));
    NOR2X1 U18838 (.A1(N7122), .A2(n14353), .ZN(N31710));
    INVX1 U18839 (.I(n27358), .ZN(N31711));
    INVX1 U18840 (.I(n16561), .ZN(N31712));
    INVX1 U18841 (.I(N8609), .ZN(n31713));
    INVX1 U18842 (.I(n12927), .ZN(N31714));
    INVX1 U18843 (.I(n21380), .ZN(N31715));
    INVX1 U18844 (.I(n27181), .ZN(n31716));
    INVX1 U18845 (.I(n21840), .ZN(N31717));
    NANDX1 U18846 (.A1(n25418), .A2(n27791), .ZN(N31718));
    NOR2X1 U18847 (.A1(n23497), .A2(N8381), .ZN(N31719));
    NOR2X1 U18848 (.A1(n15988), .A2(N8855), .ZN(N31720));
    NOR2X1 U18849 (.A1(n21137), .A2(N9639), .ZN(n31721));
    NOR2X1 U18850 (.A1(N7496), .A2(n12993), .ZN(n31722));
    NOR2X1 U18851 (.A1(n21849), .A2(N3893), .ZN(n31723));
    NANDX1 U18852 (.A1(n20205), .A2(N9014), .ZN(N31724));
    INVX1 U18853 (.I(n17374), .ZN(N31725));
    NANDX1 U18854 (.A1(n17797), .A2(N9778), .ZN(n31726));
    NOR2X1 U18855 (.A1(n25369), .A2(n25519), .ZN(n31727));
    NOR2X1 U18856 (.A1(n17071), .A2(n21990), .ZN(N31728));
    NOR2X1 U18857 (.A1(n14724), .A2(n20529), .ZN(n31729));
    NANDX1 U18858 (.A1(n23105), .A2(n24391), .ZN(n31730));
    INVX1 U18859 (.I(N1822), .ZN(N31731));
    NANDX1 U18860 (.A1(n15755), .A2(N21), .ZN(n31732));
    INVX1 U18861 (.I(n23250), .ZN(n31733));
    INVX1 U18862 (.I(n15827), .ZN(N31734));
    NANDX1 U18863 (.A1(N5467), .A2(N8552), .ZN(n31735));
    INVX1 U18864 (.I(N3042), .ZN(N31736));
    INVX1 U18865 (.I(n29661), .ZN(N31737));
    NANDX1 U18866 (.A1(N8341), .A2(n27999), .ZN(N31738));
    INVX1 U18867 (.I(N3572), .ZN(n31739));
    NANDX1 U18868 (.A1(N9226), .A2(n20642), .ZN(N31740));
    NANDX1 U18869 (.A1(n24634), .A2(n23927), .ZN(n31741));
    NANDX1 U18870 (.A1(N3264), .A2(N5455), .ZN(N31742));
    NANDX1 U18871 (.A1(n28019), .A2(N7276), .ZN(n31743));
    NOR2X1 U18872 (.A1(N2197), .A2(n25995), .ZN(N31744));
    INVX1 U18873 (.I(n25446), .ZN(N31745));
    INVX1 U18874 (.I(n26383), .ZN(N31746));
    NOR2X1 U18875 (.A1(n21596), .A2(n23496), .ZN(n31747));
    INVX1 U18876 (.I(n24637), .ZN(n31748));
    INVX1 U18877 (.I(n29339), .ZN(N31749));
    NOR2X1 U18878 (.A1(n22379), .A2(n27201), .ZN(n31750));
    NOR2X1 U18879 (.A1(n25950), .A2(n20443), .ZN(n31751));
    INVX1 U18880 (.I(N5016), .ZN(N31752));
    NOR2X1 U18881 (.A1(N12184), .A2(n28942), .ZN(N31753));
    NANDX1 U18882 (.A1(N4009), .A2(N4259), .ZN(N31754));
    NOR2X1 U18883 (.A1(N1890), .A2(N95), .ZN(n31755));
    NOR2X1 U18884 (.A1(n22784), .A2(n14650), .ZN(n31756));
    INVX1 U18885 (.I(N6653), .ZN(N31757));
    NOR2X1 U18886 (.A1(N11154), .A2(n24181), .ZN(n31758));
    INVX1 U18887 (.I(n23210), .ZN(N31759));
    NOR2X1 U18888 (.A1(n16737), .A2(N7112), .ZN(N31760));
    NOR2X1 U18889 (.A1(N5965), .A2(n29490), .ZN(N31761));
    NOR2X1 U18890 (.A1(N2989), .A2(n13864), .ZN(N31762));
    NANDX1 U18891 (.A1(N9237), .A2(n18879), .ZN(N31763));
    NOR2X1 U18892 (.A1(N9982), .A2(N6244), .ZN(N31764));
    INVX1 U18893 (.I(n13990), .ZN(N31765));
    NOR2X1 U18894 (.A1(n18365), .A2(N4440), .ZN(N31766));
    NANDX1 U18895 (.A1(n22716), .A2(n27223), .ZN(N31767));
    NOR2X1 U18896 (.A1(n26185), .A2(N3738), .ZN(N31768));
    NOR2X1 U18897 (.A1(N7202), .A2(n27919), .ZN(n31769));
    NOR2X1 U18898 (.A1(n18972), .A2(n21640), .ZN(n31770));
    INVX1 U18899 (.I(n26083), .ZN(N31771));
    NANDX1 U18900 (.A1(N6371), .A2(n25436), .ZN(N31772));
    NANDX1 U18901 (.A1(n28057), .A2(n27860), .ZN(N31773));
    INVX1 U18902 (.I(N7157), .ZN(n31774));
    NOR2X1 U18903 (.A1(n19505), .A2(n17138), .ZN(N31775));
    NANDX1 U18904 (.A1(N12314), .A2(N990), .ZN(N31776));
    INVX1 U18905 (.I(n19239), .ZN(N31777));
    INVX1 U18906 (.I(n28321), .ZN(N31778));
    NOR2X1 U18907 (.A1(n21212), .A2(n19249), .ZN(n31779));
    NOR2X1 U18908 (.A1(n24949), .A2(n22258), .ZN(n31780));
    NOR2X1 U18909 (.A1(N11291), .A2(n17366), .ZN(N31781));
    NANDX1 U18910 (.A1(N2794), .A2(n17772), .ZN(n31782));
    NOR2X1 U18911 (.A1(n17356), .A2(N12704), .ZN(N31783));
    NOR2X1 U18912 (.A1(N3207), .A2(N10623), .ZN(n31784));
    NANDX1 U18913 (.A1(n18184), .A2(n17779), .ZN(N31785));
    NANDX1 U18914 (.A1(N7551), .A2(n23477), .ZN(n31786));
    INVX1 U18915 (.I(N8425), .ZN(N31787));
    NOR2X1 U18916 (.A1(n22976), .A2(n16225), .ZN(N31788));
    INVX1 U18917 (.I(N9721), .ZN(N31789));
    NOR2X1 U18918 (.A1(N9529), .A2(n28969), .ZN(N31790));
    NOR2X1 U18919 (.A1(n23039), .A2(n21089), .ZN(N31791));
    INVX1 U18920 (.I(N4192), .ZN(n31792));
    INVX1 U18921 (.I(N12195), .ZN(N31793));
    INVX1 U18922 (.I(N3211), .ZN(N31794));
    NANDX1 U18923 (.A1(n24341), .A2(N4475), .ZN(n31795));
    NOR2X1 U18924 (.A1(n16108), .A2(n15098), .ZN(n31796));
    NANDX1 U18925 (.A1(n22852), .A2(n21437), .ZN(N31797));
    INVX1 U18926 (.I(n18963), .ZN(n31798));
    NOR2X1 U18927 (.A1(N1124), .A2(n27387), .ZN(n31799));
    NOR2X1 U18928 (.A1(n24100), .A2(n13474), .ZN(n31800));
    INVX1 U18929 (.I(N3683), .ZN(N31801));
    NOR2X1 U18930 (.A1(n14210), .A2(N2514), .ZN(N31802));
    NOR2X1 U18931 (.A1(N7111), .A2(N12164), .ZN(N31803));
    INVX1 U18932 (.I(n30001), .ZN(n31804));
    INVX1 U18933 (.I(N3318), .ZN(N31805));
    NOR2X1 U18934 (.A1(N813), .A2(N11177), .ZN(N31806));
    NOR2X1 U18935 (.A1(N5288), .A2(n28698), .ZN(N31807));
    NOR2X1 U18936 (.A1(N8946), .A2(N12027), .ZN(N31808));
    NANDX1 U18937 (.A1(n18943), .A2(N641), .ZN(n31809));
    INVX1 U18938 (.I(N3582), .ZN(N31810));
    NANDX1 U18939 (.A1(n21904), .A2(n19946), .ZN(N31811));
    NOR2X1 U18940 (.A1(n23938), .A2(n24627), .ZN(N31812));
    NANDX1 U18941 (.A1(N12438), .A2(N8699), .ZN(N31813));
    INVX1 U18942 (.I(n21224), .ZN(N31814));
    NOR2X1 U18943 (.A1(n28603), .A2(N12347), .ZN(N31815));
    NANDX1 U18944 (.A1(n26205), .A2(N4225), .ZN(n31816));
    INVX1 U18945 (.I(n27017), .ZN(N31817));
    NANDX1 U18946 (.A1(n26650), .A2(n20865), .ZN(N31818));
    NOR2X1 U18947 (.A1(n20929), .A2(n29810), .ZN(N31819));
    NANDX1 U18948 (.A1(n26621), .A2(n18616), .ZN(N31820));
    NANDX1 U18949 (.A1(N2439), .A2(N10758), .ZN(N31821));
    INVX1 U18950 (.I(n12903), .ZN(N31822));
    INVX1 U18951 (.I(n15757), .ZN(N31823));
    NANDX1 U18952 (.A1(n13753), .A2(n22423), .ZN(N31824));
    NOR2X1 U18953 (.A1(N11013), .A2(N8725), .ZN(N31825));
    INVX1 U18954 (.I(N3944), .ZN(N31826));
    NOR2X1 U18955 (.A1(N11134), .A2(n26875), .ZN(N31827));
    NOR2X1 U18956 (.A1(n15358), .A2(n15077), .ZN(N31828));
    INVX1 U18957 (.I(n19319), .ZN(N31829));
    NOR2X1 U18958 (.A1(N9562), .A2(N10402), .ZN(N31830));
    INVX1 U18959 (.I(n27933), .ZN(N31831));
    NANDX1 U18960 (.A1(n17562), .A2(N4972), .ZN(n31832));
    INVX1 U18961 (.I(N8561), .ZN(N31833));
    INVX1 U18962 (.I(n18593), .ZN(N31834));
    NANDX1 U18963 (.A1(N4856), .A2(n22910), .ZN(n31835));
    NOR2X1 U18964 (.A1(N7169), .A2(n15195), .ZN(N31836));
    NOR2X1 U18965 (.A1(n18181), .A2(N12481), .ZN(N31837));
    INVX1 U18966 (.I(n22124), .ZN(n31838));
    INVX1 U18967 (.I(n15651), .ZN(n31839));
    INVX1 U18968 (.I(N11488), .ZN(N31840));
    INVX1 U18969 (.I(n22499), .ZN(N31841));
    NANDX1 U18970 (.A1(n27448), .A2(N11209), .ZN(N31842));
    NOR2X1 U18971 (.A1(n26411), .A2(N2150), .ZN(N31843));
    NANDX1 U18972 (.A1(N9784), .A2(N8272), .ZN(n31844));
    INVX1 U18973 (.I(N4166), .ZN(N31845));
    NANDX1 U18974 (.A1(n16802), .A2(n22758), .ZN(N31846));
    INVX1 U18975 (.I(N10218), .ZN(n31847));
    NANDX1 U18976 (.A1(n13447), .A2(n17386), .ZN(N31848));
    NOR2X1 U18977 (.A1(n19177), .A2(n24128), .ZN(N31849));
    NANDX1 U18978 (.A1(n23694), .A2(n16114), .ZN(N31850));
    NOR2X1 U18979 (.A1(n27905), .A2(n23536), .ZN(N31851));
    NANDX1 U18980 (.A1(N5897), .A2(N4458), .ZN(N31852));
    NOR2X1 U18981 (.A1(N3207), .A2(n15666), .ZN(n31853));
    NOR2X1 U18982 (.A1(n29617), .A2(N6377), .ZN(N31854));
    NANDX1 U18983 (.A1(n27962), .A2(n14648), .ZN(N31855));
    NANDX1 U18984 (.A1(N1990), .A2(n20041), .ZN(n31856));
    INVX1 U18985 (.I(n13308), .ZN(N31857));
    NANDX1 U18986 (.A1(N9711), .A2(n17398), .ZN(N31858));
    NOR2X1 U18987 (.A1(n15658), .A2(N6545), .ZN(N31859));
    NANDX1 U18988 (.A1(N9648), .A2(n15432), .ZN(N31860));
    INVX1 U18989 (.I(n14322), .ZN(n31861));
    NANDX1 U18990 (.A1(n17827), .A2(N7720), .ZN(n31862));
    NOR2X1 U18991 (.A1(n23723), .A2(N738), .ZN(n31863));
    NOR2X1 U18992 (.A1(n15491), .A2(N4965), .ZN(n31864));
    NANDX1 U18993 (.A1(n14970), .A2(n30039), .ZN(N31865));
    INVX1 U18994 (.I(N1355), .ZN(n31866));
    INVX1 U18995 (.I(n17995), .ZN(N31867));
    INVX1 U18996 (.I(n23151), .ZN(N31868));
    NANDX1 U18997 (.A1(n16651), .A2(n28471), .ZN(n31869));
    INVX1 U18998 (.I(N3911), .ZN(N31870));
    NOR2X1 U18999 (.A1(N1280), .A2(n29154), .ZN(N31871));
    INVX1 U19000 (.I(N10927), .ZN(N31872));
    INVX1 U19001 (.I(n14829), .ZN(N31873));
    NANDX1 U19002 (.A1(n28298), .A2(n21216), .ZN(n31874));
    NANDX1 U19003 (.A1(N10478), .A2(n14802), .ZN(N31875));
    NOR2X1 U19004 (.A1(N2748), .A2(N155), .ZN(N31876));
    INVX1 U19005 (.I(n22112), .ZN(n31877));
    NANDX1 U19006 (.A1(n15692), .A2(N4399), .ZN(n31878));
    NOR2X1 U19007 (.A1(n18802), .A2(n22393), .ZN(n31879));
    NOR2X1 U19008 (.A1(N11815), .A2(n28441), .ZN(N31880));
    NANDX1 U19009 (.A1(n28846), .A2(n14063), .ZN(N31881));
    NANDX1 U19010 (.A1(n15809), .A2(n15342), .ZN(N31882));
    INVX1 U19011 (.I(n29276), .ZN(N31883));
    INVX1 U19012 (.I(N8090), .ZN(N31884));
    NANDX1 U19013 (.A1(n21379), .A2(n24948), .ZN(N31885));
    NANDX1 U19014 (.A1(N1331), .A2(N5288), .ZN(n31886));
    INVX1 U19015 (.I(N12157), .ZN(N31887));
    NOR2X1 U19016 (.A1(n15820), .A2(n27948), .ZN(N31888));
    NOR2X1 U19017 (.A1(n19505), .A2(N2063), .ZN(n31889));
    INVX1 U19018 (.I(n13105), .ZN(N31890));
    NANDX1 U19019 (.A1(N3922), .A2(N10048), .ZN(N31891));
    NOR2X1 U19020 (.A1(n20923), .A2(n23642), .ZN(N31892));
    INVX1 U19021 (.I(N4849), .ZN(n31893));
    INVX1 U19022 (.I(n24317), .ZN(n31894));
    NOR2X1 U19023 (.A1(n23350), .A2(N12016), .ZN(N31895));
    NANDX1 U19024 (.A1(n20001), .A2(N3104), .ZN(N31896));
    NANDX1 U19025 (.A1(n14811), .A2(n15408), .ZN(n31897));
    NOR2X1 U19026 (.A1(N8660), .A2(N12375), .ZN(n31898));
    INVX1 U19027 (.I(N5255), .ZN(N31899));
    INVX1 U19028 (.I(n14678), .ZN(N31900));
    INVX1 U19029 (.I(N6123), .ZN(n31901));
    NOR2X1 U19030 (.A1(n24189), .A2(n19227), .ZN(n31902));
    NANDX1 U19031 (.A1(n28110), .A2(n29274), .ZN(N31903));
    NANDX1 U19032 (.A1(N7457), .A2(N11340), .ZN(N31904));
    NOR2X1 U19033 (.A1(N12305), .A2(N10910), .ZN(n31905));
    INVX1 U19034 (.I(n21055), .ZN(N31906));
    INVX1 U19035 (.I(N9092), .ZN(N31907));
    INVX1 U19036 (.I(N12683), .ZN(N31908));
    NOR2X1 U19037 (.A1(n29317), .A2(n16055), .ZN(n31909));
    INVX1 U19038 (.I(N3891), .ZN(N31910));
    INVX1 U19039 (.I(n28538), .ZN(N31911));
    INVX1 U19040 (.I(N7090), .ZN(N31912));
    INVX1 U19041 (.I(N5299), .ZN(N31913));
    NOR2X1 U19042 (.A1(n21278), .A2(N10600), .ZN(n31914));
    INVX1 U19043 (.I(N10367), .ZN(N31915));
    NOR2X1 U19044 (.A1(N198), .A2(n28201), .ZN(N31916));
    INVX1 U19045 (.I(N7654), .ZN(n31917));
    INVX1 U19046 (.I(N8092), .ZN(N31918));
    INVX1 U19047 (.I(N8873), .ZN(n31919));
    INVX1 U19048 (.I(n18134), .ZN(N31920));
    INVX1 U19049 (.I(n14258), .ZN(n31921));
    INVX1 U19050 (.I(N2799), .ZN(N31922));
    NOR2X1 U19051 (.A1(N1673), .A2(N7414), .ZN(n31923));
    INVX1 U19052 (.I(n24262), .ZN(N31924));
    NOR2X1 U19053 (.A1(N10878), .A2(n14883), .ZN(N31925));
    NANDX1 U19054 (.A1(n26033), .A2(n20181), .ZN(n31926));
    INVX1 U19055 (.I(n17173), .ZN(n31927));
    INVX1 U19056 (.I(N8038), .ZN(N31928));
    INVX1 U19057 (.I(n25969), .ZN(N31929));
    INVX1 U19058 (.I(n14164), .ZN(N31930));
    INVX1 U19059 (.I(N4449), .ZN(n31931));
    NANDX1 U19060 (.A1(n16377), .A2(N1528), .ZN(N31932));
    NANDX1 U19061 (.A1(n21543), .A2(n19662), .ZN(N31933));
    NOR2X1 U19062 (.A1(N5664), .A2(n22155), .ZN(n31934));
    NOR2X1 U19063 (.A1(n20677), .A2(N12388), .ZN(n31935));
    NOR2X1 U19064 (.A1(N3017), .A2(N6512), .ZN(n31936));
    NANDX1 U19065 (.A1(N2456), .A2(n21394), .ZN(N31937));
    NOR2X1 U19066 (.A1(n28488), .A2(n30136), .ZN(n31938));
    INVX1 U19067 (.I(n15524), .ZN(N31939));
    NANDX1 U19068 (.A1(N7750), .A2(N1486), .ZN(N31940));
    NANDX1 U19069 (.A1(N4545), .A2(n15649), .ZN(N31941));
    NANDX1 U19070 (.A1(n27692), .A2(n27776), .ZN(N31942));
    NOR2X1 U19071 (.A1(n29219), .A2(n18638), .ZN(n31943));
    NANDX1 U19072 (.A1(N7304), .A2(N11055), .ZN(N31944));
    NOR2X1 U19073 (.A1(n29458), .A2(n13529), .ZN(N31945));
    NANDX1 U19074 (.A1(N270), .A2(n23417), .ZN(N31946));
    NANDX1 U19075 (.A1(n25479), .A2(N978), .ZN(N31947));
    NANDX1 U19076 (.A1(n16736), .A2(n25013), .ZN(N31948));
    NOR2X1 U19077 (.A1(N5295), .A2(n24725), .ZN(N31949));
    NANDX1 U19078 (.A1(n13195), .A2(n21035), .ZN(N31950));
    INVX1 U19079 (.I(n16926), .ZN(n31951));
    NOR2X1 U19080 (.A1(n25421), .A2(n17503), .ZN(n31952));
    INVX1 U19081 (.I(N11620), .ZN(N31953));
    INVX1 U19082 (.I(N10776), .ZN(N31954));
    INVX1 U19083 (.I(N1238), .ZN(n31955));
    NOR2X1 U19084 (.A1(N11174), .A2(n22519), .ZN(N31956));
    INVX1 U19085 (.I(n13264), .ZN(N31957));
    NANDX1 U19086 (.A1(n24928), .A2(n25241), .ZN(n31958));
    NOR2X1 U19087 (.A1(n20269), .A2(n26218), .ZN(N31959));
    INVX1 U19088 (.I(n25565), .ZN(N31960));
    INVX1 U19089 (.I(n24912), .ZN(n31961));
    NOR2X1 U19090 (.A1(N4242), .A2(n14500), .ZN(N31962));
    NANDX1 U19091 (.A1(n25276), .A2(N12833), .ZN(N31963));
    NANDX1 U19092 (.A1(N9278), .A2(n26815), .ZN(N31964));
    NOR2X1 U19093 (.A1(n20972), .A2(N8297), .ZN(N31965));
    NOR2X1 U19094 (.A1(N1610), .A2(N8417), .ZN(N31966));
    NOR2X1 U19095 (.A1(N8249), .A2(N8151), .ZN(N31967));
    NOR2X1 U19096 (.A1(N2770), .A2(n21414), .ZN(n31968));
    INVX1 U19097 (.I(n27697), .ZN(N31969));
    NOR2X1 U19098 (.A1(n19581), .A2(n17829), .ZN(n31970));
    INVX1 U19099 (.I(N10152), .ZN(N31971));
    INVX1 U19100 (.I(n29511), .ZN(n31972));
    NOR2X1 U19101 (.A1(n21237), .A2(N3615), .ZN(N31973));
    INVX1 U19102 (.I(n23713), .ZN(N31974));
    NANDX1 U19103 (.A1(n20819), .A2(N1539), .ZN(n31975));
    INVX1 U19104 (.I(n17496), .ZN(N31976));
    INVX1 U19105 (.I(n17563), .ZN(N31977));
    NOR2X1 U19106 (.A1(n15210), .A2(N7733), .ZN(n31978));
    INVX1 U19107 (.I(N4654), .ZN(N31979));
    NANDX1 U19108 (.A1(N783), .A2(n23875), .ZN(n31980));
    NANDX1 U19109 (.A1(N10758), .A2(n17159), .ZN(N31981));
    INVX1 U19110 (.I(N4397), .ZN(N31982));
    NANDX1 U19111 (.A1(N11260), .A2(n24253), .ZN(N31983));
    INVX1 U19112 (.I(n13077), .ZN(N31984));
    NOR2X1 U19113 (.A1(N10240), .A2(N4176), .ZN(N31985));
    NOR2X1 U19114 (.A1(n18226), .A2(n16449), .ZN(n31986));
    NANDX1 U19115 (.A1(n27606), .A2(n17987), .ZN(n31987));
    NOR2X1 U19116 (.A1(N3525), .A2(N3414), .ZN(N31988));
    NOR2X1 U19117 (.A1(n17878), .A2(n18623), .ZN(N31989));
    NANDX1 U19118 (.A1(N10510), .A2(N11837), .ZN(N31990));
    NOR2X1 U19119 (.A1(n29991), .A2(N5574), .ZN(N31991));
    NANDX1 U19120 (.A1(n29309), .A2(N11293), .ZN(N31992));
    INVX1 U19121 (.I(N3568), .ZN(n31993));
    NANDX1 U19122 (.A1(n18666), .A2(n16381), .ZN(N31994));
    NANDX1 U19123 (.A1(n20303), .A2(n28568), .ZN(n31995));
    NANDX1 U19124 (.A1(n13039), .A2(n14233), .ZN(N31996));
    NOR2X1 U19125 (.A1(n18049), .A2(N5909), .ZN(n31997));
    INVX1 U19126 (.I(N5898), .ZN(N31998));
    NOR2X1 U19127 (.A1(n18349), .A2(n28009), .ZN(N31999));
    NOR2X1 U19128 (.A1(n24788), .A2(N5055), .ZN(N32000));
    INVX1 U19129 (.I(N5160), .ZN(N32001));
    INVX1 U19130 (.I(n16049), .ZN(N32002));
    NOR2X1 U19131 (.A1(n29723), .A2(n30024), .ZN(n32003));
    INVX1 U19132 (.I(N10879), .ZN(N32004));
    NOR2X1 U19133 (.A1(n15010), .A2(n17334), .ZN(n32005));
    INVX1 U19134 (.I(n19952), .ZN(n32006));
    NOR2X1 U19135 (.A1(n23383), .A2(n18382), .ZN(N32007));
    INVX1 U19136 (.I(N6284), .ZN(n32008));
    NANDX1 U19137 (.A1(n15452), .A2(n12893), .ZN(n32009));
    NANDX1 U19138 (.A1(n18837), .A2(N7352), .ZN(N32010));
    INVX1 U19139 (.I(n25747), .ZN(n32011));
    INVX1 U19140 (.I(N5643), .ZN(N32012));
    INVX1 U19141 (.I(N10278), .ZN(N32013));
    NOR2X1 U19142 (.A1(n14117), .A2(N4290), .ZN(N32014));
    NANDX1 U19143 (.A1(n26389), .A2(N3876), .ZN(N32015));
    INVX1 U19144 (.I(N7694), .ZN(n32016));
    NOR2X1 U19145 (.A1(n15377), .A2(N11265), .ZN(N32017));
    INVX1 U19146 (.I(n29895), .ZN(N32018));
    NOR2X1 U19147 (.A1(N8174), .A2(n23140), .ZN(N32019));
    INVX1 U19148 (.I(N6269), .ZN(N32020));
    INVX1 U19149 (.I(n29196), .ZN(N32021));
    INVX1 U19150 (.I(N740), .ZN(n32022));
    INVX1 U19151 (.I(n17679), .ZN(n32023));
    NOR2X1 U19152 (.A1(N1643), .A2(n13288), .ZN(n32024));
    INVX1 U19153 (.I(n25983), .ZN(n32025));
    INVX1 U19154 (.I(N713), .ZN(N32026));
    INVX1 U19155 (.I(n24923), .ZN(N32027));
    INVX1 U19156 (.I(n19072), .ZN(N32028));
    NOR2X1 U19157 (.A1(N8877), .A2(n27156), .ZN(n32029));
    NANDX1 U19158 (.A1(N12191), .A2(N12395), .ZN(N32030));
    INVX1 U19159 (.I(N2701), .ZN(n32031));
    NOR2X1 U19160 (.A1(n29770), .A2(N10874), .ZN(N32032));
    NOR2X1 U19161 (.A1(N7654), .A2(N5704), .ZN(n32033));
    INVX1 U19162 (.I(n25410), .ZN(N32034));
    INVX1 U19163 (.I(n19698), .ZN(n32035));
    NANDX1 U19164 (.A1(n22224), .A2(n16350), .ZN(N32036));
    NANDX1 U19165 (.A1(N5375), .A2(n18224), .ZN(N32037));
    NANDX1 U19166 (.A1(n16180), .A2(N7497), .ZN(N32038));
    NANDX1 U19167 (.A1(N10965), .A2(N12498), .ZN(n32039));
    INVX1 U19168 (.I(N2001), .ZN(N32040));
    NOR2X1 U19169 (.A1(N107), .A2(n19429), .ZN(N32041));
    NOR2X1 U19170 (.A1(N12501), .A2(n29422), .ZN(N32042));
    NANDX1 U19171 (.A1(n13213), .A2(n17616), .ZN(n32043));
    INVX1 U19172 (.I(N6928), .ZN(n32044));
    NOR2X1 U19173 (.A1(n29964), .A2(N7188), .ZN(N32045));
    INVX1 U19174 (.I(N4372), .ZN(n32046));
    NANDX1 U19175 (.A1(n19075), .A2(n26596), .ZN(N32047));
    INVX1 U19176 (.I(n19252), .ZN(N32048));
    NANDX1 U19177 (.A1(N8443), .A2(N3835), .ZN(n32049));
    NANDX1 U19178 (.A1(n15939), .A2(n17989), .ZN(N32050));
    INVX1 U19179 (.I(n16997), .ZN(N32051));
    NOR2X1 U19180 (.A1(N8099), .A2(n15493), .ZN(n32052));
    NANDX1 U19181 (.A1(n27527), .A2(N7482), .ZN(N32053));
    NOR2X1 U19182 (.A1(n15373), .A2(n20869), .ZN(N32054));
    INVX1 U19183 (.I(N2851), .ZN(N32055));
    INVX1 U19184 (.I(N12247), .ZN(N32056));
    INVX1 U19185 (.I(n22078), .ZN(N32057));
    INVX1 U19186 (.I(N7083), .ZN(N32058));
    INVX1 U19187 (.I(n23441), .ZN(N32059));
    NOR2X1 U19188 (.A1(N11468), .A2(n25099), .ZN(n32060));
    NANDX1 U19189 (.A1(n20559), .A2(N3404), .ZN(n32061));
    NOR2X1 U19190 (.A1(n27132), .A2(N7903), .ZN(N32062));
    NANDX1 U19191 (.A1(n21791), .A2(n24900), .ZN(n32063));
    INVX1 U19192 (.I(n29889), .ZN(N32064));
    NOR2X1 U19193 (.A1(n26336), .A2(n15840), .ZN(N32065));
    NANDX1 U19194 (.A1(n18442), .A2(n19773), .ZN(N32066));
    NANDX1 U19195 (.A1(n23761), .A2(n22623), .ZN(n32067));
    INVX1 U19196 (.I(N5870), .ZN(N32068));
    INVX1 U19197 (.I(n29917), .ZN(N32069));
    NOR2X1 U19198 (.A1(N4808), .A2(n14789), .ZN(N32070));
    NOR2X1 U19199 (.A1(n19525), .A2(n26257), .ZN(n32071));
    INVX1 U19200 (.I(N11918), .ZN(n32072));
    NANDX1 U19201 (.A1(N12792), .A2(N8144), .ZN(N32073));
    NOR2X1 U19202 (.A1(n20694), .A2(n22359), .ZN(n32074));
    NANDX1 U19203 (.A1(N4017), .A2(n16073), .ZN(N32075));
    NOR2X1 U19204 (.A1(N2833), .A2(N833), .ZN(N32076));
    INVX1 U19205 (.I(N9129), .ZN(N32077));
    NANDX1 U19206 (.A1(N6371), .A2(n13416), .ZN(N32078));
    NANDX1 U19207 (.A1(n17554), .A2(n21255), .ZN(N32079));
    NANDX1 U19208 (.A1(n15279), .A2(n21034), .ZN(N32080));
    NOR2X1 U19209 (.A1(N8647), .A2(n24383), .ZN(N32081));
    NANDX1 U19210 (.A1(n28171), .A2(N9063), .ZN(N32082));
    NOR2X1 U19211 (.A1(N9951), .A2(n14302), .ZN(N32083));
    NOR2X1 U19212 (.A1(n18095), .A2(n16534), .ZN(N32084));
    INVX1 U19213 (.I(n29014), .ZN(n32085));
    NOR2X1 U19214 (.A1(n29490), .A2(n14949), .ZN(n32086));
    NOR2X1 U19215 (.A1(N2185), .A2(n15781), .ZN(N32087));
    INVX1 U19216 (.I(N11314), .ZN(N32088));
    NANDX1 U19217 (.A1(N104), .A2(n13290), .ZN(N32089));
    INVX1 U19218 (.I(N6218), .ZN(N32090));
    INVX1 U19219 (.I(N2263), .ZN(n32091));
    NOR2X1 U19220 (.A1(n14001), .A2(N575), .ZN(N32092));
    NANDX1 U19221 (.A1(N8246), .A2(N6054), .ZN(N32093));
    INVX1 U19222 (.I(n17309), .ZN(n32094));
    NOR2X1 U19223 (.A1(n15248), .A2(N1473), .ZN(n32095));
    INVX1 U19224 (.I(n21903), .ZN(n32096));
    NANDX1 U19225 (.A1(N2338), .A2(n20779), .ZN(N32097));
    NANDX1 U19226 (.A1(N1690), .A2(n24288), .ZN(N32098));
    NANDX1 U19227 (.A1(N3875), .A2(n28630), .ZN(N32099));
    NANDX1 U19228 (.A1(N3749), .A2(n22108), .ZN(n32100));
    INVX1 U19229 (.I(N5599), .ZN(N32101));
    NOR2X1 U19230 (.A1(N12735), .A2(N10005), .ZN(n32102));
    NOR2X1 U19231 (.A1(n22791), .A2(N12566), .ZN(n32103));
    NANDX1 U19232 (.A1(N11356), .A2(n20811), .ZN(N32104));
    NOR2X1 U19233 (.A1(n16653), .A2(n26680), .ZN(N32105));
    INVX1 U19234 (.I(N1763), .ZN(N32106));
    NOR2X1 U19235 (.A1(N8097), .A2(n23665), .ZN(n32107));
    NANDX1 U19236 (.A1(N10434), .A2(N2867), .ZN(N32108));
    INVX1 U19237 (.I(N684), .ZN(N32109));
    NOR2X1 U19238 (.A1(n18630), .A2(n23256), .ZN(N32110));
    INVX1 U19239 (.I(n25044), .ZN(N32111));
    INVX1 U19240 (.I(n24875), .ZN(n32112));
    NOR2X1 U19241 (.A1(n21163), .A2(N342), .ZN(n32113));
    NOR2X1 U19242 (.A1(n19728), .A2(N8207), .ZN(N32114));
    INVX1 U19243 (.I(N2156), .ZN(n32115));
    INVX1 U19244 (.I(N6729), .ZN(n32116));
    NOR2X1 U19245 (.A1(n26959), .A2(n23381), .ZN(N32117));
    NANDX1 U19246 (.A1(N9356), .A2(n13704), .ZN(N32118));
    NANDX1 U19247 (.A1(N6013), .A2(n25929), .ZN(N32119));
    NOR2X1 U19248 (.A1(N5007), .A2(n28795), .ZN(n32120));
    NOR2X1 U19249 (.A1(n24389), .A2(N2934), .ZN(N32121));
    NOR2X1 U19250 (.A1(n17507), .A2(n17140), .ZN(n32122));
    NANDX1 U19251 (.A1(n21633), .A2(N11878), .ZN(n32123));
    INVX1 U19252 (.I(N1219), .ZN(N32124));
    NANDX1 U19253 (.A1(n30112), .A2(n20947), .ZN(n32125));
    NOR2X1 U19254 (.A1(n25485), .A2(N11663), .ZN(n32126));
    INVX1 U19255 (.I(n20775), .ZN(N32127));
    INVX1 U19256 (.I(n18274), .ZN(n32128));
    NANDX1 U19257 (.A1(n27080), .A2(n16190), .ZN(N32129));
    NANDX1 U19258 (.A1(N10286), .A2(n22203), .ZN(N32130));
    NANDX1 U19259 (.A1(N5332), .A2(n15770), .ZN(n32131));
    INVX1 U19260 (.I(N6325), .ZN(n32132));
    INVX1 U19261 (.I(N2226), .ZN(n32133));
    NANDX1 U19262 (.A1(n16089), .A2(N7926), .ZN(N32134));
    NOR2X1 U19263 (.A1(N7584), .A2(N8364), .ZN(N32135));
    INVX1 U19264 (.I(N8802), .ZN(N32136));
    NANDX1 U19265 (.A1(N3389), .A2(n18309), .ZN(N32137));
    NANDX1 U19266 (.A1(n28874), .A2(n18533), .ZN(N32138));
    NANDX1 U19267 (.A1(N8072), .A2(n18844), .ZN(n32139));
    INVX1 U19268 (.I(N10650), .ZN(n32140));
    NOR2X1 U19269 (.A1(n21028), .A2(n26932), .ZN(N32141));
    NANDX1 U19270 (.A1(N1654), .A2(n27567), .ZN(n32142));
    NOR2X1 U19271 (.A1(n17423), .A2(n15420), .ZN(N32143));
    NANDX1 U19272 (.A1(n27444), .A2(N6206), .ZN(N32144));
    INVX1 U19273 (.I(N1956), .ZN(N32145));
    NOR2X1 U19274 (.A1(N9559), .A2(N9539), .ZN(N32146));
    NANDX1 U19275 (.A1(n24412), .A2(N6901), .ZN(N32147));
    INVX1 U19276 (.I(n27800), .ZN(N32148));
    NANDX1 U19277 (.A1(N4009), .A2(n15097), .ZN(n32149));
    NOR2X1 U19278 (.A1(N2013), .A2(n23168), .ZN(N32150));
    NOR2X1 U19279 (.A1(n25548), .A2(n22379), .ZN(N32151));
    INVX1 U19280 (.I(N4999), .ZN(N32152));
    NOR2X1 U19281 (.A1(n28548), .A2(N6652), .ZN(N32153));
    NANDX1 U19282 (.A1(N6935), .A2(N12636), .ZN(N32154));
    NOR2X1 U19283 (.A1(n21783), .A2(n28640), .ZN(N32155));
    NANDX1 U19284 (.A1(N2304), .A2(N458), .ZN(n32156));
    NOR2X1 U19285 (.A1(N11862), .A2(N9996), .ZN(n32157));
    INVX1 U19286 (.I(N6136), .ZN(n32158));
    NOR2X1 U19287 (.A1(N7716), .A2(n22496), .ZN(n32159));
    INVX1 U19288 (.I(N11725), .ZN(N32160));
    NOR2X1 U19289 (.A1(N9953), .A2(N2298), .ZN(N32161));
    NOR2X1 U19290 (.A1(n19523), .A2(n16406), .ZN(N32162));
    NANDX1 U19291 (.A1(n22000), .A2(n21405), .ZN(n32163));
    NANDX1 U19292 (.A1(n20410), .A2(n28056), .ZN(N32164));
    NOR2X1 U19293 (.A1(n15905), .A2(N10554), .ZN(N32165));
    INVX1 U19294 (.I(N7550), .ZN(n32166));
    NANDX1 U19295 (.A1(N7235), .A2(n28551), .ZN(N32167));
    NANDX1 U19296 (.A1(n25274), .A2(N10275), .ZN(n32168));
    INVX1 U19297 (.I(N12792), .ZN(n32169));
    NOR2X1 U19298 (.A1(N2087), .A2(N9069), .ZN(n32170));
    INVX1 U19299 (.I(N9874), .ZN(N32171));
    NANDX1 U19300 (.A1(n23483), .A2(n19827), .ZN(n32172));
    INVX1 U19301 (.I(N12529), .ZN(N32173));
    INVX1 U19302 (.I(n16617), .ZN(N32174));
    INVX1 U19303 (.I(n19772), .ZN(N32175));
    INVX1 U19304 (.I(n12975), .ZN(N32176));
    NANDX1 U19305 (.A1(N5803), .A2(n25856), .ZN(N32177));
    NANDX1 U19306 (.A1(N4917), .A2(n17743), .ZN(n32178));
    NOR2X1 U19307 (.A1(n21232), .A2(n13539), .ZN(N32179));
    NOR2X1 U19308 (.A1(n19305), .A2(n27373), .ZN(n32180));
    INVX1 U19309 (.I(N4496), .ZN(n32181));
    NANDX1 U19310 (.A1(N12840), .A2(n25280), .ZN(N32182));
    NANDX1 U19311 (.A1(n28867), .A2(N5016), .ZN(N32183));
    NOR2X1 U19312 (.A1(N10773), .A2(n24842), .ZN(N32184));
    INVX1 U19313 (.I(n23301), .ZN(n32185));
    NOR2X1 U19314 (.A1(n15139), .A2(N5678), .ZN(N32186));
    NANDX1 U19315 (.A1(N11584), .A2(N7213), .ZN(N32187));
    INVX1 U19316 (.I(N5947), .ZN(n32188));
    NANDX1 U19317 (.A1(n21182), .A2(n29561), .ZN(N32189));
    INVX1 U19318 (.I(N1664), .ZN(N32190));
    NOR2X1 U19319 (.A1(N11334), .A2(N10697), .ZN(n32191));
    NOR2X1 U19320 (.A1(N8570), .A2(N7127), .ZN(N32192));
    NOR2X1 U19321 (.A1(N7158), .A2(N8527), .ZN(N32193));
    INVX1 U19322 (.I(n26253), .ZN(n32194));
    NANDX1 U19323 (.A1(n21734), .A2(n13125), .ZN(N32195));
    NANDX1 U19324 (.A1(N5000), .A2(N208), .ZN(n32196));
    INVX1 U19325 (.I(n16174), .ZN(n32197));
    INVX1 U19326 (.I(N12689), .ZN(n32198));
    NANDX1 U19327 (.A1(n15490), .A2(n19901), .ZN(N32199));
    NOR2X1 U19328 (.A1(n21436), .A2(N11393), .ZN(N32200));
    NANDX1 U19329 (.A1(n20860), .A2(N9189), .ZN(N32201));
    INVX1 U19330 (.I(n30075), .ZN(n32202));
    INVX1 U19331 (.I(n22879), .ZN(N32203));
    NOR2X1 U19332 (.A1(N6213), .A2(n30005), .ZN(n32204));
    NANDX1 U19333 (.A1(n13370), .A2(N8394), .ZN(n32205));
    NOR2X1 U19334 (.A1(n28183), .A2(N4210), .ZN(n32206));
    INVX1 U19335 (.I(n29868), .ZN(n32207));
    NANDX1 U19336 (.A1(n14513), .A2(n30075), .ZN(n32208));
    NANDX1 U19337 (.A1(N549), .A2(n22543), .ZN(N32209));
    NOR2X1 U19338 (.A1(n24790), .A2(N7895), .ZN(N32210));
    NOR2X1 U19339 (.A1(N6868), .A2(n17892), .ZN(n32211));
    INVX1 U19340 (.I(N10127), .ZN(N32212));
    INVX1 U19341 (.I(n17962), .ZN(n32213));
    INVX1 U19342 (.I(n27249), .ZN(N32214));
    NANDX1 U19343 (.A1(n15050), .A2(n25570), .ZN(n32215));
    INVX1 U19344 (.I(n14917), .ZN(N32216));
    NOR2X1 U19345 (.A1(N5051), .A2(n23310), .ZN(n32217));
    NOR2X1 U19346 (.A1(n21794), .A2(n16080), .ZN(N32218));
    NOR2X1 U19347 (.A1(n21525), .A2(n15438), .ZN(N32219));
    INVX1 U19348 (.I(N10023), .ZN(n32220));
    INVX1 U19349 (.I(n16243), .ZN(n32221));
    NANDX1 U19350 (.A1(n22165), .A2(N10896), .ZN(N32222));
    INVX1 U19351 (.I(N848), .ZN(N32223));
    NOR2X1 U19352 (.A1(N5336), .A2(n21060), .ZN(N32224));
    NOR2X1 U19353 (.A1(N2510), .A2(n27583), .ZN(N32225));
    NOR2X1 U19354 (.A1(n18319), .A2(n13051), .ZN(N32226));
    NANDX1 U19355 (.A1(n13751), .A2(N4731), .ZN(n32227));
    NANDX1 U19356 (.A1(n17641), .A2(n28479), .ZN(N32228));
    INVX1 U19357 (.I(n20749), .ZN(N32229));
    NANDX1 U19358 (.A1(n13521), .A2(n21931), .ZN(N32230));
    NOR2X1 U19359 (.A1(n28958), .A2(N7488), .ZN(n32231));
    NOR2X1 U19360 (.A1(n20626), .A2(N12291), .ZN(N32232));
    NANDX1 U19361 (.A1(N1214), .A2(N11747), .ZN(N32233));
    NANDX1 U19362 (.A1(N2061), .A2(n18071), .ZN(N32234));
    NANDX1 U19363 (.A1(N11682), .A2(n23082), .ZN(N32235));
    NOR2X1 U19364 (.A1(N9127), .A2(n20264), .ZN(N32236));
    INVX1 U19365 (.I(N10738), .ZN(N32237));
    INVX1 U19366 (.I(n28452), .ZN(N32238));
    NOR2X1 U19367 (.A1(N6627), .A2(n15955), .ZN(n32239));
    NOR2X1 U19368 (.A1(N4068), .A2(n25264), .ZN(N32240));
    NANDX1 U19369 (.A1(n17588), .A2(n17057), .ZN(n32241));
    INVX1 U19370 (.I(N4969), .ZN(n32242));
    NANDX1 U19371 (.A1(n21255), .A2(n14155), .ZN(N32243));
    NOR2X1 U19372 (.A1(N3651), .A2(n15369), .ZN(N32244));
    NANDX1 U19373 (.A1(N3628), .A2(n17429), .ZN(n32245));
    NANDX1 U19374 (.A1(N8940), .A2(n17671), .ZN(N32246));
    NANDX1 U19375 (.A1(N5322), .A2(n26797), .ZN(N32247));
    NOR2X1 U19376 (.A1(N1325), .A2(n26095), .ZN(n32248));
    INVX1 U19377 (.I(n18337), .ZN(N32249));
    NANDX1 U19378 (.A1(N1509), .A2(n22852), .ZN(N32250));
    INVX1 U19379 (.I(N5576), .ZN(N32251));
    NANDX1 U19380 (.A1(n13423), .A2(N11724), .ZN(N32252));
    NANDX1 U19381 (.A1(n24572), .A2(n16692), .ZN(N32253));
    INVX1 U19382 (.I(N4250), .ZN(n32254));
    NANDX1 U19383 (.A1(n20517), .A2(n26599), .ZN(N32255));
    NANDX1 U19384 (.A1(n16082), .A2(N89), .ZN(n32256));
    NOR2X1 U19385 (.A1(n18278), .A2(n27727), .ZN(N32257));
    NANDX1 U19386 (.A1(n13418), .A2(N2911), .ZN(n32258));
    INVX1 U19387 (.I(n17382), .ZN(N32259));
    INVX1 U19388 (.I(n20915), .ZN(N32260));
    INVX1 U19389 (.I(N11132), .ZN(n32261));
    NANDX1 U19390 (.A1(N2333), .A2(N3846), .ZN(N32262));
    NANDX1 U19391 (.A1(N7908), .A2(N10384), .ZN(N32263));
    INVX1 U19392 (.I(n19631), .ZN(N32264));
    INVX1 U19393 (.I(N8235), .ZN(N32265));
    NOR2X1 U19394 (.A1(n29100), .A2(N12485), .ZN(N32266));
    NANDX1 U19395 (.A1(N8041), .A2(N8946), .ZN(N32267));
    INVX1 U19396 (.I(N12683), .ZN(n32268));
    NANDX1 U19397 (.A1(n22158), .A2(N824), .ZN(N32269));
    INVX1 U19398 (.I(N1621), .ZN(n32270));
    INVX1 U19399 (.I(n16793), .ZN(n32271));
    NANDX1 U19400 (.A1(n20184), .A2(N9588), .ZN(N32272));
    NANDX1 U19401 (.A1(N2310), .A2(n20720), .ZN(N32273));
    INVX1 U19402 (.I(N4643), .ZN(N32274));
    NANDX1 U19403 (.A1(n19936), .A2(N1111), .ZN(N32275));
    NANDX1 U19404 (.A1(n15039), .A2(N9303), .ZN(N32276));
    NOR2X1 U19405 (.A1(N11834), .A2(N4048), .ZN(N32277));
    NANDX1 U19406 (.A1(n24318), .A2(n29639), .ZN(N32278));
    NOR2X1 U19407 (.A1(n21824), .A2(n18292), .ZN(N32279));
    NOR2X1 U19408 (.A1(N7980), .A2(N10312), .ZN(N32280));
    NANDX1 U19409 (.A1(N3163), .A2(N493), .ZN(n32281));
    NOR2X1 U19410 (.A1(n19955), .A2(n27070), .ZN(N32282));
    NANDX1 U19411 (.A1(n18104), .A2(N2849), .ZN(N32283));
    INVX1 U19412 (.I(n27384), .ZN(n32284));
    NANDX1 U19413 (.A1(N9160), .A2(N10372), .ZN(n32285));
    NANDX1 U19414 (.A1(N10271), .A2(n22442), .ZN(n32286));
    NOR2X1 U19415 (.A1(N8134), .A2(N8216), .ZN(N32287));
    INVX1 U19416 (.I(N12181), .ZN(N32288));
    NOR2X1 U19417 (.A1(N6198), .A2(N244), .ZN(n32289));
    NOR2X1 U19418 (.A1(n28022), .A2(n18535), .ZN(N32290));
    NOR2X1 U19419 (.A1(N5864), .A2(n28846), .ZN(N32291));
    NANDX1 U19420 (.A1(n27724), .A2(n29339), .ZN(N32292));
    NANDX1 U19421 (.A1(N6103), .A2(n14832), .ZN(N32293));
    INVX1 U19422 (.I(n24206), .ZN(N32294));
    NOR2X1 U19423 (.A1(N736), .A2(N10013), .ZN(N32295));
    NANDX1 U19424 (.A1(N9896), .A2(n20384), .ZN(N32296));
    INVX1 U19425 (.I(N8727), .ZN(n32297));
    NOR2X1 U19426 (.A1(n13975), .A2(n16860), .ZN(N32298));
    NANDX1 U19427 (.A1(n25992), .A2(n29040), .ZN(n32299));
    NANDX1 U19428 (.A1(N2053), .A2(n17844), .ZN(n32300));
    NANDX1 U19429 (.A1(n18635), .A2(N6241), .ZN(N32301));
    INVX1 U19430 (.I(n13059), .ZN(N32302));
    NOR2X1 U19431 (.A1(N7809), .A2(n29343), .ZN(N32303));
    INVX1 U19432 (.I(n27776), .ZN(N32304));
    INVX1 U19433 (.I(n14802), .ZN(N32305));
    NANDX1 U19434 (.A1(n18074), .A2(n21043), .ZN(n32306));
    NOR2X1 U19435 (.A1(n28086), .A2(n15371), .ZN(n32307));
    NANDX1 U19436 (.A1(N6894), .A2(N6284), .ZN(N32308));
    INVX1 U19437 (.I(n19582), .ZN(N32309));
    NANDX1 U19438 (.A1(n25893), .A2(n17607), .ZN(N32310));
    NANDX1 U19439 (.A1(n24795), .A2(n27281), .ZN(N32311));
    NOR2X1 U19440 (.A1(N12502), .A2(N7063), .ZN(N32312));
    INVX1 U19441 (.I(N7303), .ZN(N32313));
    NANDX1 U19442 (.A1(n26979), .A2(N813), .ZN(N32314));
    NANDX1 U19443 (.A1(n26185), .A2(N783), .ZN(N32315));
    NOR2X1 U19444 (.A1(n20053), .A2(n15585), .ZN(N32316));
    NANDX1 U19445 (.A1(N7990), .A2(N6490), .ZN(N32317));
    INVX1 U19446 (.I(n24636), .ZN(N32318));
    NOR2X1 U19447 (.A1(n19967), .A2(N1392), .ZN(N32319));
    NANDX1 U19448 (.A1(N10302), .A2(N9534), .ZN(N32320));
    INVX1 U19449 (.I(N6057), .ZN(N32321));
    NOR2X1 U19450 (.A1(N60), .A2(n19412), .ZN(n32322));
    NANDX1 U19451 (.A1(n25484), .A2(n20474), .ZN(n32323));
    NOR2X1 U19452 (.A1(N9267), .A2(n27777), .ZN(n32324));
    NANDX1 U19453 (.A1(N6109), .A2(n17150), .ZN(N32325));
    NOR2X1 U19454 (.A1(N2156), .A2(n17933), .ZN(n32326));
    NANDX1 U19455 (.A1(n22208), .A2(N3380), .ZN(N32327));
    INVX1 U19456 (.I(n18758), .ZN(N32328));
    NOR2X1 U19457 (.A1(n20112), .A2(N1818), .ZN(N32329));
    NOR2X1 U19458 (.A1(N9941), .A2(n21907), .ZN(N32330));
    NANDX1 U19459 (.A1(N8803), .A2(N1304), .ZN(n32331));
    NANDX1 U19460 (.A1(N3420), .A2(N5565), .ZN(n32332));
    NOR2X1 U19461 (.A1(n22832), .A2(n18409), .ZN(N32333));
    NOR2X1 U19462 (.A1(N1729), .A2(n15436), .ZN(n32334));
    INVX1 U19463 (.I(n18066), .ZN(n32335));
    NANDX1 U19464 (.A1(n27540), .A2(n23777), .ZN(N32336));
    NANDX1 U19465 (.A1(n18256), .A2(N11572), .ZN(N32337));
    NANDX1 U19466 (.A1(n29025), .A2(N3512), .ZN(n32338));
    NANDX1 U19467 (.A1(N6206), .A2(n20639), .ZN(N32339));
    INVX1 U19468 (.I(N8023), .ZN(N32340));
    NOR2X1 U19469 (.A1(N11170), .A2(n29930), .ZN(N32341));
    NOR2X1 U19470 (.A1(N8534), .A2(n19794), .ZN(N32342));
    INVX1 U19471 (.I(N11953), .ZN(N32343));
    NOR2X1 U19472 (.A1(N12727), .A2(N4647), .ZN(n32344));
    INVX1 U19473 (.I(n24892), .ZN(N32345));
    INVX1 U19474 (.I(n17626), .ZN(N32346));
    INVX1 U19475 (.I(n13002), .ZN(N32347));
    INVX1 U19476 (.I(N2150), .ZN(N32348));
    NOR2X1 U19477 (.A1(N12297), .A2(N8967), .ZN(N32349));
    NOR2X1 U19478 (.A1(N221), .A2(N7854), .ZN(N32350));
    INVX1 U19479 (.I(N11475), .ZN(N32351));
    INVX1 U19480 (.I(n19483), .ZN(N32352));
    INVX1 U19481 (.I(N10643), .ZN(N32353));
    NANDX1 U19482 (.A1(N996), .A2(N10435), .ZN(N32354));
    INVX1 U19483 (.I(N9529), .ZN(N32355));
    INVX1 U19484 (.I(N1148), .ZN(N32356));
    INVX1 U19485 (.I(n14009), .ZN(N32357));
    NOR2X1 U19486 (.A1(n14689), .A2(n16199), .ZN(n32358));
    NANDX1 U19487 (.A1(N9625), .A2(N3687), .ZN(N32359));
    NOR2X1 U19488 (.A1(N11187), .A2(N10703), .ZN(n32360));
    NANDX1 U19489 (.A1(n17828), .A2(N11560), .ZN(N32361));
    NANDX1 U19490 (.A1(n13161), .A2(N11780), .ZN(N32362));
    NOR2X1 U19491 (.A1(N12006), .A2(n23255), .ZN(N32363));
    INVX1 U19492 (.I(N1351), .ZN(n32364));
    NOR2X1 U19493 (.A1(N4030), .A2(n16004), .ZN(N32365));
    NANDX1 U19494 (.A1(N3025), .A2(n21244), .ZN(n32366));
    INVX1 U19495 (.I(N3115), .ZN(N32367));
    INVX1 U19496 (.I(N3508), .ZN(n32368));
    NOR2X1 U19497 (.A1(N6129), .A2(N6757), .ZN(N32369));
    INVX1 U19498 (.I(N3318), .ZN(N32370));
    NANDX1 U19499 (.A1(n14130), .A2(N5255), .ZN(n32371));
    NOR2X1 U19500 (.A1(n13393), .A2(N9341), .ZN(N32372));
    NANDX1 U19501 (.A1(n24953), .A2(n22393), .ZN(N32373));
    INVX1 U19502 (.I(N6595), .ZN(N32374));
    NANDX1 U19503 (.A1(n17545), .A2(n18410), .ZN(n32375));
    NANDX1 U19504 (.A1(N7456), .A2(N1353), .ZN(n32376));
    INVX1 U19505 (.I(n23460), .ZN(N32377));
    NANDX1 U19506 (.A1(n20861), .A2(n14566), .ZN(N32378));
    NOR2X1 U19507 (.A1(N12537), .A2(n25518), .ZN(N32379));
    NANDX1 U19508 (.A1(n18221), .A2(n20207), .ZN(N32380));
    INVX1 U19509 (.I(n28664), .ZN(n32381));
    INVX1 U19510 (.I(N8478), .ZN(N32382));
    INVX1 U19511 (.I(n17340), .ZN(N32383));
    INVX1 U19512 (.I(n14609), .ZN(N32384));
    NOR2X1 U19513 (.A1(N5545), .A2(N9424), .ZN(N32385));
    INVX1 U19514 (.I(N11084), .ZN(N32386));
    NOR2X1 U19515 (.A1(N9217), .A2(n28628), .ZN(N32387));
    NANDX1 U19516 (.A1(N4325), .A2(N5946), .ZN(N32388));
    NANDX1 U19517 (.A1(N10722), .A2(n29405), .ZN(N32389));
    INVX1 U19518 (.I(N1446), .ZN(n32390));
    INVX1 U19519 (.I(n21602), .ZN(n32391));
    NANDX1 U19520 (.A1(n27912), .A2(n18382), .ZN(N32392));
    INVX1 U19521 (.I(N6543), .ZN(N32393));
    NOR2X1 U19522 (.A1(n19289), .A2(n18628), .ZN(N32394));
    NANDX1 U19523 (.A1(n20505), .A2(N5830), .ZN(n32395));
    NOR2X1 U19524 (.A1(n23674), .A2(N2372), .ZN(N32396));
    NOR2X1 U19525 (.A1(N2961), .A2(N9867), .ZN(N32397));
    NOR2X1 U19526 (.A1(N7540), .A2(n19083), .ZN(n32398));
    NOR2X1 U19527 (.A1(n19089), .A2(N11968), .ZN(N32399));
    NANDX1 U19528 (.A1(N1854), .A2(n22690), .ZN(N32400));
    NANDX1 U19529 (.A1(N7304), .A2(n24135), .ZN(N32401));
    NOR2X1 U19530 (.A1(n17466), .A2(n26677), .ZN(n32402));
    INVX1 U19531 (.I(n24408), .ZN(n32403));
    NANDX1 U19532 (.A1(n13406), .A2(n16188), .ZN(N32404));
    INVX1 U19533 (.I(N1896), .ZN(N32405));
    NANDX1 U19534 (.A1(n15518), .A2(n26423), .ZN(N32406));
    NANDX1 U19535 (.A1(N9054), .A2(n28794), .ZN(N32407));
    NANDX1 U19536 (.A1(N575), .A2(n27221), .ZN(N32408));
    INVX1 U19537 (.I(n26812), .ZN(N32409));
    INVX1 U19538 (.I(n15911), .ZN(N32410));
    NANDX1 U19539 (.A1(n16694), .A2(n27518), .ZN(N32411));
    NANDX1 U19540 (.A1(N9246), .A2(n15514), .ZN(N32412));
    NOR2X1 U19541 (.A1(n21941), .A2(N5905), .ZN(n32413));
    INVX1 U19542 (.I(n18480), .ZN(n32414));
    NOR2X1 U19543 (.A1(n13777), .A2(N5644), .ZN(n32415));
    NOR2X1 U19544 (.A1(n18525), .A2(N657), .ZN(N32416));
    NOR2X1 U19545 (.A1(N12091), .A2(N4735), .ZN(n32417));
    INVX1 U19546 (.I(N7640), .ZN(N32418));
    INVX1 U19547 (.I(N131), .ZN(N32419));
    INVX1 U19548 (.I(N2924), .ZN(N32420));
    NOR2X1 U19549 (.A1(n20966), .A2(n18297), .ZN(N32421));
    INVX1 U19550 (.I(N6739), .ZN(N32422));
    NOR2X1 U19551 (.A1(n18633), .A2(n22817), .ZN(n32423));
    INVX1 U19552 (.I(n16440), .ZN(N32424));
    NOR2X1 U19553 (.A1(n19400), .A2(N8243), .ZN(N32425));
    INVX1 U19554 (.I(N8769), .ZN(N32426));
    NANDX1 U19555 (.A1(N3986), .A2(N11106), .ZN(N32427));
    INVX1 U19556 (.I(n18719), .ZN(N32428));
    NOR2X1 U19557 (.A1(N10145), .A2(N5210), .ZN(N32429));
    INVX1 U19558 (.I(n14879), .ZN(N32430));
    NOR2X1 U19559 (.A1(n26481), .A2(n17228), .ZN(N32431));
    NOR2X1 U19560 (.A1(n25759), .A2(N8713), .ZN(N32432));
    NANDX1 U19561 (.A1(N5148), .A2(n27009), .ZN(N32433));
    NOR2X1 U19562 (.A1(N447), .A2(n19492), .ZN(N32434));
    NOR2X1 U19563 (.A1(n23263), .A2(N6713), .ZN(N32435));
    INVX1 U19564 (.I(N8577), .ZN(n32436));
    INVX1 U19565 (.I(n14963), .ZN(N32437));
    NANDX1 U19566 (.A1(n23441), .A2(N109), .ZN(N32438));
    NOR2X1 U19567 (.A1(n23107), .A2(N9597), .ZN(N32439));
    INVX1 U19568 (.I(N11160), .ZN(N32440));
    INVX1 U19569 (.I(n27709), .ZN(N32441));
    NANDX1 U19570 (.A1(N11741), .A2(N4256), .ZN(N32442));
    NOR2X1 U19571 (.A1(n17530), .A2(N11069), .ZN(n32443));
    NANDX1 U19572 (.A1(n26242), .A2(N3657), .ZN(N32444));
    NANDX1 U19573 (.A1(N11674), .A2(n28320), .ZN(N32445));
    NANDX1 U19574 (.A1(n19726), .A2(n30040), .ZN(N32446));
    NOR2X1 U19575 (.A1(n26438), .A2(n18062), .ZN(N32447));
    INVX1 U19576 (.I(N10973), .ZN(N32448));
    NOR2X1 U19577 (.A1(n24875), .A2(N4276), .ZN(N32449));
    INVX1 U19578 (.I(n28655), .ZN(n32450));
    NOR2X1 U19579 (.A1(N1153), .A2(n21017), .ZN(N32451));
    NOR2X1 U19580 (.A1(N9454), .A2(N7150), .ZN(n32452));
    NANDX1 U19581 (.A1(N9756), .A2(n30103), .ZN(n32453));
    INVX1 U19582 (.I(n27285), .ZN(N32454));
    INVX1 U19583 (.I(n29517), .ZN(N32455));
    NANDX1 U19584 (.A1(N3251), .A2(N3613), .ZN(N32456));
    NOR2X1 U19585 (.A1(n20132), .A2(N8293), .ZN(n32457));
    NANDX1 U19586 (.A1(n20034), .A2(n24795), .ZN(n32458));
    INVX1 U19587 (.I(N7959), .ZN(N32459));
    INVX1 U19588 (.I(n27742), .ZN(N32460));
    NOR2X1 U19589 (.A1(N3035), .A2(n20578), .ZN(N32461));
    NOR2X1 U19590 (.A1(N1553), .A2(N6383), .ZN(n32462));
    NANDX1 U19591 (.A1(N11130), .A2(n22045), .ZN(n32463));
    NANDX1 U19592 (.A1(N6840), .A2(N7433), .ZN(N32464));
    NANDX1 U19593 (.A1(N6805), .A2(N7725), .ZN(N32465));
    NOR2X1 U19594 (.A1(N6400), .A2(N7104), .ZN(N32466));
    INVX1 U19595 (.I(n28348), .ZN(n32467));
    NOR2X1 U19596 (.A1(n21164), .A2(n18342), .ZN(n32468));
    INVX1 U19597 (.I(n22935), .ZN(N32469));
    NANDX1 U19598 (.A1(n20925), .A2(N9567), .ZN(n32470));
    NANDX1 U19599 (.A1(n29223), .A2(N7171), .ZN(N32471));
    INVX1 U19600 (.I(N2120), .ZN(N32472));
    NANDX1 U19601 (.A1(N6565), .A2(n22370), .ZN(N32473));
    INVX1 U19602 (.I(n17378), .ZN(N32474));
    NANDX1 U19603 (.A1(n14598), .A2(N7508), .ZN(N32475));
    NANDX1 U19604 (.A1(N10591), .A2(N7392), .ZN(N32476));
    INVX1 U19605 (.I(n18316), .ZN(n32477));
    INVX1 U19606 (.I(n19226), .ZN(n32478));
    NOR2X1 U19607 (.A1(n13404), .A2(n17436), .ZN(n32479));
    NANDX1 U19608 (.A1(N4431), .A2(N5641), .ZN(N32480));
    NOR2X1 U19609 (.A1(n27365), .A2(n13879), .ZN(N32481));
    INVX1 U19610 (.I(n25493), .ZN(N32482));
    NANDX1 U19611 (.A1(N10699), .A2(n21224), .ZN(N32483));
    NANDX1 U19612 (.A1(N1379), .A2(N7396), .ZN(n32484));
    NANDX1 U19613 (.A1(N12310), .A2(n30086), .ZN(n32485));
    INVX1 U19614 (.I(n22931), .ZN(n32486));
    INVX1 U19615 (.I(N1233), .ZN(n32487));
    NANDX1 U19616 (.A1(n13698), .A2(N8624), .ZN(n32488));
    NANDX1 U19617 (.A1(n20574), .A2(n13047), .ZN(N32489));
    INVX1 U19618 (.I(N4417), .ZN(N32490));
    INVX1 U19619 (.I(n29604), .ZN(N32491));
    NANDX1 U19620 (.A1(N8003), .A2(N5107), .ZN(N32492));
    NANDX1 U19621 (.A1(n23928), .A2(N7546), .ZN(n32493));
    NOR2X1 U19622 (.A1(n19283), .A2(n14742), .ZN(N32494));
    NANDX1 U19623 (.A1(N10370), .A2(n26101), .ZN(n32495));
    INVX1 U19624 (.I(n17765), .ZN(N32496));
    INVX1 U19625 (.I(N10043), .ZN(n32497));
    NANDX1 U19626 (.A1(n26310), .A2(n21534), .ZN(N32498));
    NOR2X1 U19627 (.A1(n16103), .A2(N1651), .ZN(n32499));
    NANDX1 U19628 (.A1(n24727), .A2(n24730), .ZN(N32500));
    INVX1 U19629 (.I(n26334), .ZN(N32501));
    NANDX1 U19630 (.A1(n13751), .A2(n29906), .ZN(N32502));
    INVX1 U19631 (.I(n19985), .ZN(n32503));
    INVX1 U19632 (.I(N11333), .ZN(n32504));
    NOR2X1 U19633 (.A1(N1562), .A2(N7439), .ZN(N32505));
    NANDX1 U19634 (.A1(n20844), .A2(n22180), .ZN(N32506));
    NOR2X1 U19635 (.A1(n19774), .A2(N6704), .ZN(N32507));
    INVX1 U19636 (.I(n26099), .ZN(N32508));
    INVX1 U19637 (.I(N10875), .ZN(n32509));
    INVX1 U19638 (.I(N12583), .ZN(n32510));
    INVX1 U19639 (.I(n18875), .ZN(N32511));
    NANDX1 U19640 (.A1(n22619), .A2(n19075), .ZN(n32512));
    INVX1 U19641 (.I(n17212), .ZN(N32513));
    NOR2X1 U19642 (.A1(N8032), .A2(n23972), .ZN(N32514));
    NOR2X1 U19643 (.A1(N7800), .A2(n18759), .ZN(n32515));
    INVX1 U19644 (.I(N4132), .ZN(n32516));
    INVX1 U19645 (.I(N7337), .ZN(N32517));
    NANDX1 U19646 (.A1(n26090), .A2(N2641), .ZN(n32518));
    INVX1 U19647 (.I(N6693), .ZN(N32519));
    NOR2X1 U19648 (.A1(n23432), .A2(N1957), .ZN(n32520));
    NANDX1 U19649 (.A1(n19393), .A2(n29805), .ZN(N32521));
    NANDX1 U19650 (.A1(N10189), .A2(N12250), .ZN(N32522));
    NOR2X1 U19651 (.A1(n29064), .A2(n29496), .ZN(n32523));
    NANDX1 U19652 (.A1(N6562), .A2(N11193), .ZN(n32524));
    INVX1 U19653 (.I(n23532), .ZN(N32525));
    INVX1 U19654 (.I(N7623), .ZN(N32526));
    NOR2X1 U19655 (.A1(N4146), .A2(n26381), .ZN(N32527));
    NOR2X1 U19656 (.A1(N8277), .A2(n14895), .ZN(N32528));
    NOR2X1 U19657 (.A1(N2530), .A2(n29545), .ZN(n32529));
    INVX1 U19658 (.I(N6187), .ZN(n32530));
    NOR2X1 U19659 (.A1(n18823), .A2(n29618), .ZN(N32531));
    NANDX1 U19660 (.A1(N2515), .A2(n18874), .ZN(N32532));
    INVX1 U19661 (.I(n27218), .ZN(n32533));
    NANDX1 U19662 (.A1(N8534), .A2(N12615), .ZN(n32534));
    NOR2X1 U19663 (.A1(n26590), .A2(n20631), .ZN(N32535));
    NANDX1 U19664 (.A1(N7645), .A2(N4282), .ZN(n32536));
    INVX1 U19665 (.I(N3991), .ZN(n32537));
    INVX1 U19666 (.I(n17742), .ZN(n32538));
    NANDX1 U19667 (.A1(n15406), .A2(N2151), .ZN(N32539));
    NANDX1 U19668 (.A1(N163), .A2(N12594), .ZN(N32540));
    NOR2X1 U19669 (.A1(n18268), .A2(n25677), .ZN(n32541));
    NANDX1 U19670 (.A1(n24367), .A2(N2923), .ZN(N32542));
    NOR2X1 U19671 (.A1(n20983), .A2(N5437), .ZN(N32543));
    NOR2X1 U19672 (.A1(n17267), .A2(N2517), .ZN(N32544));
    NANDX1 U19673 (.A1(n25800), .A2(n15132), .ZN(n32545));
    NANDX1 U19674 (.A1(n22252), .A2(n24323), .ZN(n32546));
    INVX1 U19675 (.I(n18457), .ZN(N32547));
    NANDX1 U19676 (.A1(n14315), .A2(n22447), .ZN(N32548));
    NOR2X1 U19677 (.A1(N1920), .A2(N7704), .ZN(n32549));
    INVX1 U19678 (.I(n22768), .ZN(N32550));
    INVX1 U19679 (.I(n21759), .ZN(n32551));
    NOR2X1 U19680 (.A1(n27436), .A2(N9890), .ZN(N32552));
    NOR2X1 U19681 (.A1(n18246), .A2(N4119), .ZN(N32553));
    INVX1 U19682 (.I(n27234), .ZN(N32554));
    INVX1 U19683 (.I(n27820), .ZN(n32555));
    NANDX1 U19684 (.A1(N12231), .A2(n18898), .ZN(n32556));
    INVX1 U19685 (.I(n26591), .ZN(N32557));
    INVX1 U19686 (.I(N486), .ZN(N32558));
    NANDX1 U19687 (.A1(n16775), .A2(n21174), .ZN(N32559));
    NOR2X1 U19688 (.A1(n15242), .A2(n24050), .ZN(N32560));
    NANDX1 U19689 (.A1(N2735), .A2(n14530), .ZN(n32561));
    INVX1 U19690 (.I(n24331), .ZN(N32562));
    NANDX1 U19691 (.A1(n15533), .A2(n15952), .ZN(N32563));
    NANDX1 U19692 (.A1(N1392), .A2(n25841), .ZN(N32564));
    NANDX1 U19693 (.A1(N8198), .A2(n18521), .ZN(N32565));
    NANDX1 U19694 (.A1(N5294), .A2(N2046), .ZN(n32566));
    NOR2X1 U19695 (.A1(N114), .A2(n14276), .ZN(N32567));
    INVX1 U19696 (.I(N10281), .ZN(N32568));
    NOR2X1 U19697 (.A1(n17502), .A2(n29464), .ZN(n32569));
    INVX1 U19698 (.I(N4139), .ZN(N32570));
    NOR2X1 U19699 (.A1(n20837), .A2(N7942), .ZN(n32571));
    NOR2X1 U19700 (.A1(n15990), .A2(n29374), .ZN(n32572));
    INVX1 U19701 (.I(N149), .ZN(N32573));
    NANDX1 U19702 (.A1(n13223), .A2(N4242), .ZN(n32574));
    NANDX1 U19703 (.A1(N2727), .A2(n24331), .ZN(N32575));
    NOR2X1 U19704 (.A1(N11691), .A2(n21090), .ZN(N32576));
    NOR2X1 U19705 (.A1(n12902), .A2(n14944), .ZN(N32577));
    NOR2X1 U19706 (.A1(n19054), .A2(n15058), .ZN(n32578));
    NANDX1 U19707 (.A1(n13966), .A2(n13899), .ZN(N32579));
    INVX1 U19708 (.I(N1330), .ZN(n32580));
    INVX1 U19709 (.I(N11451), .ZN(N32581));
    NANDX1 U19710 (.A1(N10847), .A2(N2150), .ZN(N32582));
    NOR2X1 U19711 (.A1(N2381), .A2(n18140), .ZN(N32583));
    NANDX1 U19712 (.A1(n19883), .A2(N6849), .ZN(N32584));
    NOR2X1 U19713 (.A1(n21666), .A2(n29788), .ZN(N32585));
    NANDX1 U19714 (.A1(n24392), .A2(N12542), .ZN(N32586));
    NANDX1 U19715 (.A1(N5946), .A2(N3494), .ZN(N32587));
    INVX1 U19716 (.I(N7408), .ZN(n32588));
    INVX1 U19717 (.I(n24036), .ZN(N32589));
    INVX1 U19718 (.I(N10617), .ZN(N32590));
    INVX1 U19719 (.I(n28987), .ZN(n32591));
    NANDX1 U19720 (.A1(n15841), .A2(N179), .ZN(N32592));
    NANDX1 U19721 (.A1(n27291), .A2(n24344), .ZN(N32593));
    NOR2X1 U19722 (.A1(n18001), .A2(n26314), .ZN(n32594));
    NANDX1 U19723 (.A1(n24701), .A2(n27519), .ZN(N32595));
    NOR2X1 U19724 (.A1(N1412), .A2(N10715), .ZN(n32596));
    NANDX1 U19725 (.A1(n19760), .A2(n14730), .ZN(N32597));
    NOR2X1 U19726 (.A1(N2165), .A2(N951), .ZN(N32598));
    INVX1 U19727 (.I(n24356), .ZN(N32599));
    NOR2X1 U19728 (.A1(N1350), .A2(N1217), .ZN(N32600));
    NANDX1 U19729 (.A1(n27810), .A2(N11833), .ZN(n32601));
    NOR2X1 U19730 (.A1(n15220), .A2(n13469), .ZN(N32602));
    INVX1 U19731 (.I(N3959), .ZN(N32603));
    NOR2X1 U19732 (.A1(n24431), .A2(n28302), .ZN(N32604));
    NANDX1 U19733 (.A1(N12294), .A2(n13039), .ZN(n32605));
    NOR2X1 U19734 (.A1(N6858), .A2(n29119), .ZN(N32606));
    NANDX1 U19735 (.A1(n26967), .A2(N9696), .ZN(N32607));
    NANDX1 U19736 (.A1(n16590), .A2(n12986), .ZN(N32608));
    NANDX1 U19737 (.A1(N7315), .A2(N2497), .ZN(n32609));
    NANDX1 U19738 (.A1(n20231), .A2(N1833), .ZN(N32610));
    NANDX1 U19739 (.A1(N10009), .A2(n13765), .ZN(n32611));
    NOR2X1 U19740 (.A1(N10402), .A2(n25202), .ZN(n32612));
    INVX1 U19741 (.I(n23871), .ZN(N32613));
    NANDX1 U19742 (.A1(n29383), .A2(n22063), .ZN(n32614));
    NANDX1 U19743 (.A1(n16108), .A2(n23084), .ZN(N32615));
    INVX1 U19744 (.I(n29147), .ZN(N32616));
    INVX1 U19745 (.I(n24346), .ZN(N32617));
    INVX1 U19746 (.I(N4543), .ZN(N32618));
    INVX1 U19747 (.I(n14945), .ZN(N32619));
    NOR2X1 U19748 (.A1(n14887), .A2(n27930), .ZN(n32620));
    INVX1 U19749 (.I(n22201), .ZN(N32621));
    INVX1 U19750 (.I(n13379), .ZN(N32622));
    NOR2X1 U19751 (.A1(n20819), .A2(N7214), .ZN(N32623));
    NOR2X1 U19752 (.A1(N4446), .A2(n17419), .ZN(N32624));
    NOR2X1 U19753 (.A1(n29647), .A2(N12706), .ZN(N32625));
    NOR2X1 U19754 (.A1(n21851), .A2(N11951), .ZN(N32626));
    NOR2X1 U19755 (.A1(N8348), .A2(n28058), .ZN(n32627));
    INVX1 U19756 (.I(n14397), .ZN(N32628));
    NOR2X1 U19757 (.A1(n29182), .A2(n27304), .ZN(N32629));
    INVX1 U19758 (.I(n22285), .ZN(n32630));
    INVX1 U19759 (.I(N5684), .ZN(N32631));
    NANDX1 U19760 (.A1(n21789), .A2(N3476), .ZN(n32632));
    NANDX1 U19761 (.A1(N2413), .A2(n22462), .ZN(N32633));
    NANDX1 U19762 (.A1(n21965), .A2(n13143), .ZN(N32634));
    NOR2X1 U19763 (.A1(N2691), .A2(N6149), .ZN(N32635));
    INVX1 U19764 (.I(n23955), .ZN(n32636));
    NANDX1 U19765 (.A1(n14389), .A2(n27513), .ZN(N32637));
    NANDX1 U19766 (.A1(n14900), .A2(n22996), .ZN(N32638));
    INVX1 U19767 (.I(N1382), .ZN(N32639));
    INVX1 U19768 (.I(n27374), .ZN(N32640));
    INVX1 U19769 (.I(n29167), .ZN(N32641));
    NANDX1 U19770 (.A1(N7749), .A2(n21315), .ZN(N32642));
    NANDX1 U19771 (.A1(N1993), .A2(N5673), .ZN(N32643));
    NOR2X1 U19772 (.A1(N5469), .A2(n29622), .ZN(N32644));
    NOR2X1 U19773 (.A1(n16491), .A2(N6674), .ZN(N32645));
    NOR2X1 U19774 (.A1(n18195), .A2(N9638), .ZN(n32646));
    NANDX1 U19775 (.A1(n24343), .A2(N11321), .ZN(n32647));
    INVX1 U19776 (.I(n30001), .ZN(n32648));
    NOR2X1 U19777 (.A1(n25732), .A2(n15932), .ZN(n32649));
    INVX1 U19778 (.I(N7151), .ZN(N32650));
    NANDX1 U19779 (.A1(N414), .A2(n18575), .ZN(n32651));
    NOR2X1 U19780 (.A1(N5984), .A2(N6166), .ZN(N32652));
    NANDX1 U19781 (.A1(N2293), .A2(n27480), .ZN(N32653));
    INVX1 U19782 (.I(N4285), .ZN(N32654));
    NOR2X1 U19783 (.A1(n29324), .A2(n28451), .ZN(N32655));
    INVX1 U19784 (.I(n20511), .ZN(N32656));
    NOR2X1 U19785 (.A1(n27871), .A2(N3525), .ZN(N32657));
    NANDX1 U19786 (.A1(n26069), .A2(n19367), .ZN(N32658));
    INVX1 U19787 (.I(N7252), .ZN(n32659));
    NOR2X1 U19788 (.A1(n15628), .A2(N10083), .ZN(n32660));
    NANDX1 U19789 (.A1(n20121), .A2(N9116), .ZN(N32661));
    NANDX1 U19790 (.A1(N7453), .A2(n28227), .ZN(N32662));
    NANDX1 U19791 (.A1(n22158), .A2(N4073), .ZN(N32663));
    NOR2X1 U19792 (.A1(N1128), .A2(N6365), .ZN(n32664));
    NANDX1 U19793 (.A1(n18798), .A2(N10650), .ZN(N32665));
    INVX1 U19794 (.I(n17984), .ZN(N32666));
    INVX1 U19795 (.I(n20868), .ZN(N32667));
    NOR2X1 U19796 (.A1(N12328), .A2(N7162), .ZN(N32668));
    NANDX1 U19797 (.A1(N3750), .A2(N3093), .ZN(N32669));
    INVX1 U19798 (.I(n19515), .ZN(N32670));
    NOR2X1 U19799 (.A1(n25955), .A2(n23703), .ZN(N32671));
    NOR2X1 U19800 (.A1(n16257), .A2(N2247), .ZN(n32672));
    NANDX1 U19801 (.A1(n13709), .A2(N9699), .ZN(N32673));
    NOR2X1 U19802 (.A1(n18297), .A2(n20417), .ZN(N32674));
    NOR2X1 U19803 (.A1(n29050), .A2(n21544), .ZN(n32675));
    NOR2X1 U19804 (.A1(N7008), .A2(N10204), .ZN(N32676));
    INVX1 U19805 (.I(N6679), .ZN(N32677));
    NANDX1 U19806 (.A1(N11924), .A2(n27546), .ZN(N32678));
    INVX1 U19807 (.I(n24251), .ZN(N32679));
    NOR2X1 U19808 (.A1(n25546), .A2(n16562), .ZN(n32680));
    INVX1 U19809 (.I(n15216), .ZN(n32681));
    INVX1 U19810 (.I(N6566), .ZN(N32682));
    NANDX1 U19811 (.A1(n18202), .A2(n15553), .ZN(n32683));
    INVX1 U19812 (.I(n20449), .ZN(n32684));
    NANDX1 U19813 (.A1(n29559), .A2(N10), .ZN(N32685));
    NOR2X1 U19814 (.A1(n17718), .A2(N8988), .ZN(N32686));
    NANDX1 U19815 (.A1(N5192), .A2(n19092), .ZN(n32687));
    NANDX1 U19816 (.A1(N12199), .A2(n17857), .ZN(n32688));
    INVX1 U19817 (.I(n18877), .ZN(N32689));
    NANDX1 U19818 (.A1(n24291), .A2(N4846), .ZN(N32690));
    INVX1 U19819 (.I(N6965), .ZN(N32691));
    INVX1 U19820 (.I(n13540), .ZN(n32692));
    NOR2X1 U19821 (.A1(N5637), .A2(n17316), .ZN(N32693));
    INVX1 U19822 (.I(N764), .ZN(N32694));
    INVX1 U19823 (.I(N6090), .ZN(N32695));
    NOR2X1 U19824 (.A1(n21320), .A2(n15099), .ZN(N32696));
    NOR2X1 U19825 (.A1(n20741), .A2(N3669), .ZN(n32697));
    NANDX1 U19826 (.A1(n27020), .A2(N12656), .ZN(N32698));
    NOR2X1 U19827 (.A1(N2074), .A2(N1611), .ZN(n32699));
    NANDX1 U19828 (.A1(N2833), .A2(n19467), .ZN(N32700));
    NANDX1 U19829 (.A1(N10271), .A2(n23933), .ZN(n32701));
    NANDX1 U19830 (.A1(n15116), .A2(N488), .ZN(N32702));
    NANDX1 U19831 (.A1(n13092), .A2(n14027), .ZN(N32703));
    NANDX1 U19832 (.A1(N7289), .A2(n19904), .ZN(N32704));
    INVX1 U19833 (.I(N8052), .ZN(N32705));
    NOR2X1 U19834 (.A1(N12778), .A2(n24368), .ZN(N32706));
    INVX1 U19835 (.I(n27876), .ZN(N32707));
    NANDX1 U19836 (.A1(N7160), .A2(N1407), .ZN(n32708));
    INVX1 U19837 (.I(n22740), .ZN(N32709));
    NANDX1 U19838 (.A1(N3112), .A2(n13374), .ZN(N32710));
    NOR2X1 U19839 (.A1(n19219), .A2(n16206), .ZN(n32711));
    NOR2X1 U19840 (.A1(n28996), .A2(n26476), .ZN(N32712));
    NANDX1 U19841 (.A1(n21486), .A2(N16), .ZN(N32713));
    NANDX1 U19842 (.A1(N9502), .A2(N1668), .ZN(N32714));
    NANDX1 U19843 (.A1(N9605), .A2(N8956), .ZN(n32715));
    INVX1 U19844 (.I(n16293), .ZN(N32716));
    INVX1 U19845 (.I(N5572), .ZN(n32717));
    NOR2X1 U19846 (.A1(n29936), .A2(n22128), .ZN(N32718));
    NOR2X1 U19847 (.A1(n21121), .A2(n17848), .ZN(N32719));
    INVX1 U19848 (.I(n13351), .ZN(N32720));
    INVX1 U19849 (.I(n19398), .ZN(n32721));
    NANDX1 U19850 (.A1(n23823), .A2(n23631), .ZN(N32722));
    NOR2X1 U19851 (.A1(n28589), .A2(N5754), .ZN(N32723));
    INVX1 U19852 (.I(n13489), .ZN(n32724));
    INVX1 U19853 (.I(N3009), .ZN(N32725));
    NOR2X1 U19854 (.A1(n18353), .A2(N12510), .ZN(N32726));
    INVX1 U19855 (.I(n27483), .ZN(n32727));
    NANDX1 U19856 (.A1(n24126), .A2(n26380), .ZN(N32728));
    NOR2X1 U19857 (.A1(n29694), .A2(n20512), .ZN(n32729));
    NOR2X1 U19858 (.A1(n29492), .A2(N1063), .ZN(N32730));
    NANDX1 U19859 (.A1(N9036), .A2(n18910), .ZN(N32731));
    NOR2X1 U19860 (.A1(n22386), .A2(n29359), .ZN(N32732));
    NOR2X1 U19861 (.A1(n27408), .A2(n23044), .ZN(N32733));
    NANDX1 U19862 (.A1(n21512), .A2(n21496), .ZN(n32734));
    NOR2X1 U19863 (.A1(n14473), .A2(n23545), .ZN(N32735));
    INVX1 U19864 (.I(n17481), .ZN(N32736));
    NANDX1 U19865 (.A1(N817), .A2(n18552), .ZN(N32737));
    NOR2X1 U19866 (.A1(n16861), .A2(n29226), .ZN(N32738));
    INVX1 U19867 (.I(n13103), .ZN(n32739));
    NOR2X1 U19868 (.A1(n22885), .A2(n22175), .ZN(N32740));
    NANDX1 U19869 (.A1(N10800), .A2(n23238), .ZN(N32741));
    NANDX1 U19870 (.A1(n19836), .A2(N12010), .ZN(N32742));
    NANDX1 U19871 (.A1(N12084), .A2(n29930), .ZN(N32743));
    INVX1 U19872 (.I(n28053), .ZN(N32744));
    INVX1 U19873 (.I(N4420), .ZN(N32745));
    INVX1 U19874 (.I(n21453), .ZN(n32746));
    INVX1 U19875 (.I(N3762), .ZN(N32747));
    NOR2X1 U19876 (.A1(N10555), .A2(n21243), .ZN(N32748));
    NANDX1 U19877 (.A1(N11372), .A2(N9657), .ZN(N32749));
    INVX1 U19878 (.I(n28232), .ZN(N32750));
    INVX1 U19879 (.I(n14163), .ZN(n32751));
    NANDX1 U19880 (.A1(n23361), .A2(n25608), .ZN(N32752));
    INVX1 U19881 (.I(n22300), .ZN(n32753));
    NOR2X1 U19882 (.A1(n22291), .A2(n20929), .ZN(N32754));
    NANDX1 U19883 (.A1(n22862), .A2(n13145), .ZN(N32755));
    NANDX1 U19884 (.A1(n22654), .A2(N11086), .ZN(N32756));
    NOR2X1 U19885 (.A1(N3913), .A2(n15506), .ZN(n32757));
    NOR2X1 U19886 (.A1(n13927), .A2(N2020), .ZN(N32758));
    NOR2X1 U19887 (.A1(n28786), .A2(N1135), .ZN(N32759));
    NOR2X1 U19888 (.A1(N8980), .A2(N12506), .ZN(N32760));
    INVX1 U19889 (.I(n29951), .ZN(n32761));
    NANDX1 U19890 (.A1(N11602), .A2(N2537), .ZN(N32762));
    INVX1 U19891 (.I(N4825), .ZN(N32763));
    INVX1 U19892 (.I(n28109), .ZN(N32764));
    INVX1 U19893 (.I(n22975), .ZN(N32765));
    INVX1 U19894 (.I(n25174), .ZN(n32766));
    NOR2X1 U19895 (.A1(n12986), .A2(N8181), .ZN(n32767));
    NANDX1 U19896 (.A1(N5502), .A2(N7828), .ZN(n32768));
    NANDX1 U19897 (.A1(n28113), .A2(n23333), .ZN(N32769));
    NANDX1 U19898 (.A1(N11902), .A2(n13913), .ZN(N32770));
    NANDX1 U19899 (.A1(n29248), .A2(N3608), .ZN(N32771));
    NANDX1 U19900 (.A1(N8090), .A2(N4675), .ZN(N32772));
    NOR2X1 U19901 (.A1(n26602), .A2(N3835), .ZN(N32773));
    INVX1 U19902 (.I(n17699), .ZN(N32774));
    NOR2X1 U19903 (.A1(N8475), .A2(N4267), .ZN(n32775));
    INVX1 U19904 (.I(n24160), .ZN(n32776));
    NANDX1 U19905 (.A1(n28244), .A2(N7757), .ZN(N32777));
    NANDX1 U19906 (.A1(N11093), .A2(N4499), .ZN(N32778));
    INVX1 U19907 (.I(N5155), .ZN(N32779));
    NANDX1 U19908 (.A1(n29139), .A2(N3130), .ZN(n32780));
    NOR2X1 U19909 (.A1(n26115), .A2(N3592), .ZN(N32781));
    NOR2X1 U19910 (.A1(n29366), .A2(N2703), .ZN(N32782));
    NANDX1 U19911 (.A1(n18558), .A2(n29490), .ZN(n32783));
    NANDX1 U19912 (.A1(n22046), .A2(n25954), .ZN(N32784));
    INVX1 U19913 (.I(N6998), .ZN(N32785));
    INVX1 U19914 (.I(n18682), .ZN(N32786));
    NANDX1 U19915 (.A1(N6343), .A2(n26664), .ZN(N32787));
    NANDX1 U19916 (.A1(n22144), .A2(n24770), .ZN(N32788));
    NOR2X1 U19917 (.A1(N3871), .A2(N5725), .ZN(N32789));
    NOR2X1 U19918 (.A1(n27109), .A2(n29578), .ZN(N32790));
    INVX1 U19919 (.I(n14672), .ZN(n32791));
    NANDX1 U19920 (.A1(N5277), .A2(N10649), .ZN(N32792));
    NOR2X1 U19921 (.A1(N1831), .A2(N9877), .ZN(N32793));
    NOR2X1 U19922 (.A1(N1993), .A2(n28434), .ZN(N32794));
    NOR2X1 U19923 (.A1(n25526), .A2(N8904), .ZN(N32795));
    NANDX1 U19924 (.A1(n22757), .A2(N4462), .ZN(N32796));
    NANDX1 U19925 (.A1(N11301), .A2(N8495), .ZN(N32797));
    INVX1 U19926 (.I(N7827), .ZN(N32798));
    NOR2X1 U19927 (.A1(N11716), .A2(n21158), .ZN(N32799));
    NOR2X1 U19928 (.A1(N4147), .A2(n15443), .ZN(N32800));
    NOR2X1 U19929 (.A1(n19817), .A2(n14883), .ZN(N32801));
    NANDX1 U19930 (.A1(N4351), .A2(N6014), .ZN(N32802));
    INVX1 U19931 (.I(n14999), .ZN(n32803));
    NANDX1 U19932 (.A1(N2477), .A2(n24875), .ZN(N32804));
    NANDX1 U19933 (.A1(n23167), .A2(N11732), .ZN(n32805));
    NANDX1 U19934 (.A1(n18555), .A2(n20635), .ZN(n32806));
    NOR2X1 U19935 (.A1(N11175), .A2(n13658), .ZN(N32807));
    NANDX1 U19936 (.A1(N11036), .A2(n22152), .ZN(n32808));
    NANDX1 U19937 (.A1(n18863), .A2(n17263), .ZN(N32809));
    NANDX1 U19938 (.A1(n28581), .A2(n25444), .ZN(N32810));
    NOR2X1 U19939 (.A1(n13886), .A2(n21056), .ZN(N32811));
    NOR2X1 U19940 (.A1(n28769), .A2(n27864), .ZN(N32812));
    NANDX1 U19941 (.A1(N4645), .A2(n28510), .ZN(N32813));
    NOR2X1 U19942 (.A1(n24078), .A2(n19547), .ZN(N32814));
    NOR2X1 U19943 (.A1(N10798), .A2(N12576), .ZN(n32815));
    INVX1 U19944 (.I(N1553), .ZN(n32816));
    NOR2X1 U19945 (.A1(n22661), .A2(n15039), .ZN(N32817));
    NOR2X1 U19946 (.A1(N6181), .A2(N315), .ZN(N32818));
    NANDX1 U19947 (.A1(n16893), .A2(n16740), .ZN(N32819));
    INVX1 U19948 (.I(n22716), .ZN(N32820));
    INVX1 U19949 (.I(N6191), .ZN(N32821));
    NOR2X1 U19950 (.A1(N12711), .A2(n20076), .ZN(N32822));
    NOR2X1 U19951 (.A1(N11798), .A2(N7268), .ZN(N32823));
    INVX1 U19952 (.I(n26674), .ZN(N32824));
    NOR2X1 U19953 (.A1(N859), .A2(N3533), .ZN(N32825));
    INVX1 U19954 (.I(n20405), .ZN(n32826));
    NOR2X1 U19955 (.A1(N5210), .A2(n21541), .ZN(n32827));
    NANDX1 U19956 (.A1(N6763), .A2(n29793), .ZN(N32828));
    INVX1 U19957 (.I(N10362), .ZN(N32829));
    INVX1 U19958 (.I(n13254), .ZN(N32830));
    NOR2X1 U19959 (.A1(N7966), .A2(N9), .ZN(n32831));
    NANDX1 U19960 (.A1(n15713), .A2(n22725), .ZN(N32832));
    NOR2X1 U19961 (.A1(N10464), .A2(n17868), .ZN(N32833));
    NOR2X1 U19962 (.A1(n19101), .A2(N3930), .ZN(N32834));
    NOR2X1 U19963 (.A1(n26368), .A2(n17856), .ZN(n32835));
    INVX1 U19964 (.I(n26841), .ZN(n32836));
    INVX1 U19965 (.I(N9539), .ZN(N32837));
    NANDX1 U19966 (.A1(n27680), .A2(N3365), .ZN(N32838));
    NANDX1 U19967 (.A1(n19083), .A2(N10656), .ZN(n32839));
    NANDX1 U19968 (.A1(N7299), .A2(n29168), .ZN(n32840));
    NANDX1 U19969 (.A1(n26380), .A2(N845), .ZN(N32841));
    NANDX1 U19970 (.A1(n22906), .A2(N854), .ZN(N32842));
    NANDX1 U19971 (.A1(N8482), .A2(N12139), .ZN(n32843));
    NANDX1 U19972 (.A1(N7506), .A2(n30006), .ZN(n32844));
    INVX1 U19973 (.I(n26606), .ZN(n32845));
    NOR2X1 U19974 (.A1(N9323), .A2(n22837), .ZN(N32846));
    INVX1 U19975 (.I(n15329), .ZN(n32847));
    NOR2X1 U19976 (.A1(n17489), .A2(n13428), .ZN(N32848));
    INVX1 U19977 (.I(n15031), .ZN(N32849));
    NANDX1 U19978 (.A1(N2800), .A2(n22675), .ZN(N32850));
    NOR2X1 U19979 (.A1(n13146), .A2(n29973), .ZN(N32851));
    NOR2X1 U19980 (.A1(n22414), .A2(n14776), .ZN(N32852));
    INVX1 U19981 (.I(N12221), .ZN(N32853));
    NANDX1 U19982 (.A1(n23996), .A2(n25262), .ZN(N32854));
    NOR2X1 U19983 (.A1(n24695), .A2(n16005), .ZN(n32855));
    NOR2X1 U19984 (.A1(n24563), .A2(N4419), .ZN(n32856));
    NOR2X1 U19985 (.A1(n16922), .A2(N2303), .ZN(n32857));
    INVX1 U19986 (.I(n15697), .ZN(N32858));
    INVX1 U19987 (.I(n16619), .ZN(N32859));
    NANDX1 U19988 (.A1(n19619), .A2(N4395), .ZN(N32860));
    NOR2X1 U19989 (.A1(n24971), .A2(N7195), .ZN(n32861));
    INVX1 U19990 (.I(N10842), .ZN(N32862));
    NANDX1 U19991 (.A1(n29150), .A2(N3003), .ZN(N32863));
    NANDX1 U19992 (.A1(n13788), .A2(n26145), .ZN(n32864));
    INVX1 U19993 (.I(N9893), .ZN(n32865));
    NANDX1 U19994 (.A1(n27220), .A2(n14479), .ZN(N32866));
    INVX1 U19995 (.I(N1648), .ZN(N32867));
    NANDX1 U19996 (.A1(n27683), .A2(N6066), .ZN(N32868));
    NANDX1 U19997 (.A1(N3029), .A2(n27066), .ZN(N32869));
    NOR2X1 U19998 (.A1(n18725), .A2(N3120), .ZN(n32870));
    NOR2X1 U19999 (.A1(N10334), .A2(n22738), .ZN(N32871));
    INVX1 U20000 (.I(n16974), .ZN(N32872));
    NOR2X1 U20001 (.A1(N142), .A2(n16150), .ZN(N32873));
    NANDX1 U20002 (.A1(N9043), .A2(N3723), .ZN(N32874));
    INVX1 U20003 (.I(N10220), .ZN(N32875));
    INVX1 U20004 (.I(N4544), .ZN(N32876));
    INVX1 U20005 (.I(n27403), .ZN(N32877));
    NOR2X1 U20006 (.A1(N9260), .A2(N306), .ZN(N32878));
    NOR2X1 U20007 (.A1(N10907), .A2(n26876), .ZN(N32879));
    NOR2X1 U20008 (.A1(N5533), .A2(n20430), .ZN(N32880));
    NOR2X1 U20009 (.A1(N2462), .A2(N11063), .ZN(N32881));
    INVX1 U20010 (.I(N5581), .ZN(N32882));
    INVX1 U20011 (.I(N4283), .ZN(N32883));
    NOR2X1 U20012 (.A1(N11261), .A2(n21256), .ZN(N32884));
    NANDX1 U20013 (.A1(n30101), .A2(N7268), .ZN(N32885));
    NOR2X1 U20014 (.A1(N9006), .A2(N10991), .ZN(N32886));
    NANDX1 U20015 (.A1(n19225), .A2(n17062), .ZN(N32887));
    NANDX1 U20016 (.A1(N1265), .A2(N2888), .ZN(N32888));
    NANDX1 U20017 (.A1(n29222), .A2(N3193), .ZN(n32889));
    NANDX1 U20018 (.A1(N9991), .A2(n30068), .ZN(N32890));
    NANDX1 U20019 (.A1(n15523), .A2(N8921), .ZN(n32891));
    INVX1 U20020 (.I(n17984), .ZN(N32892));
    NOR2X1 U20021 (.A1(n23767), .A2(n23565), .ZN(N32893));
    NOR2X1 U20022 (.A1(n28049), .A2(N10307), .ZN(n32894));
    NOR2X1 U20023 (.A1(n19167), .A2(n21879), .ZN(n32895));
    INVX1 U20024 (.I(n14995), .ZN(N32896));
    NOR2X1 U20025 (.A1(N5510), .A2(n25985), .ZN(n32897));
    INVX1 U20026 (.I(n13295), .ZN(n32898));
    NANDX1 U20027 (.A1(N4404), .A2(N3120), .ZN(N32899));
    NANDX1 U20028 (.A1(N6121), .A2(N2204), .ZN(N32900));
    NOR2X1 U20029 (.A1(N5366), .A2(N12194), .ZN(N32901));
    NOR2X1 U20030 (.A1(n18384), .A2(n16277), .ZN(n32902));
    INVX1 U20031 (.I(N6625), .ZN(n32903));
    INVX1 U20032 (.I(N2067), .ZN(n32904));
    NOR2X1 U20033 (.A1(n16249), .A2(n28923), .ZN(N32905));
    NANDX1 U20034 (.A1(n15116), .A2(N6766), .ZN(N32906));
    INVX1 U20035 (.I(N6857), .ZN(N32907));
    INVX1 U20036 (.I(N9448), .ZN(N32908));
    NANDX1 U20037 (.A1(n27477), .A2(n23993), .ZN(N32909));
    INVX1 U20038 (.I(N10634), .ZN(n32910));
    NOR2X1 U20039 (.A1(n24461), .A2(N2314), .ZN(N32911));
    NANDX1 U20040 (.A1(N444), .A2(N4517), .ZN(N32912));
    NANDX1 U20041 (.A1(n24507), .A2(N5271), .ZN(n32913));
    INVX1 U20042 (.I(N1314), .ZN(n32914));
    INVX1 U20043 (.I(n22753), .ZN(n32915));
    NANDX1 U20044 (.A1(N2793), .A2(n24819), .ZN(N32916));
    NANDX1 U20045 (.A1(N7602), .A2(n23604), .ZN(N32917));
    INVX1 U20046 (.I(N11278), .ZN(N32918));
    INVX1 U20047 (.I(N8068), .ZN(n32919));
    NANDX1 U20048 (.A1(N10761), .A2(N6076), .ZN(N32920));
    NOR2X1 U20049 (.A1(N8101), .A2(n30069), .ZN(n32921));
    NOR2X1 U20050 (.A1(N7295), .A2(n13955), .ZN(n32922));
    INVX1 U20051 (.I(N9609), .ZN(N32923));
    NANDX1 U20052 (.A1(n25782), .A2(N2686), .ZN(N32924));
    NOR2X1 U20053 (.A1(N8713), .A2(n26655), .ZN(n32925));
    INVX1 U20054 (.I(N10026), .ZN(N32926));
    NANDX1 U20055 (.A1(n19835), .A2(n17964), .ZN(n32927));
    NANDX1 U20056 (.A1(N3077), .A2(n14717), .ZN(n32928));
    NANDX1 U20057 (.A1(n15241), .A2(n16893), .ZN(n32929));
    NANDX1 U20058 (.A1(N4034), .A2(n24960), .ZN(N32930));
    NOR2X1 U20059 (.A1(N3356), .A2(N899), .ZN(N32931));
    NANDX1 U20060 (.A1(N11456), .A2(n19528), .ZN(n32932));
    NOR2X1 U20061 (.A1(N7311), .A2(N3345), .ZN(n32933));
    NOR2X1 U20062 (.A1(N5480), .A2(N5542), .ZN(n32934));
    INVX1 U20063 (.I(N8166), .ZN(N32935));
    INVX1 U20064 (.I(n23507), .ZN(N32936));
    NANDX1 U20065 (.A1(N7872), .A2(N3395), .ZN(N32937));
    NOR2X1 U20066 (.A1(n16267), .A2(N9920), .ZN(n32938));
    NANDX1 U20067 (.A1(n19343), .A2(n24636), .ZN(N32939));
    INVX1 U20068 (.I(n23145), .ZN(N32940));
    NANDX1 U20069 (.A1(N4663), .A2(n15739), .ZN(n32941));
    NANDX1 U20070 (.A1(n16774), .A2(n19094), .ZN(N32942));
    NANDX1 U20071 (.A1(N9706), .A2(n19110), .ZN(N32943));
    NANDX1 U20072 (.A1(n14956), .A2(n26421), .ZN(N32944));
    NANDX1 U20073 (.A1(N3969), .A2(N1763), .ZN(n32945));
    INVX1 U20074 (.I(n18763), .ZN(N32946));
    NANDX1 U20075 (.A1(N557), .A2(N693), .ZN(N32947));
    INVX1 U20076 (.I(n27126), .ZN(N32948));
    NANDX1 U20077 (.A1(n17557), .A2(n13256), .ZN(N32949));
    NANDX1 U20078 (.A1(n22662), .A2(n21159), .ZN(N32950));
    INVX1 U20079 (.I(n21907), .ZN(n32951));
    NOR2X1 U20080 (.A1(n15714), .A2(n15130), .ZN(N32952));
    NANDX1 U20081 (.A1(n29186), .A2(N1766), .ZN(N32953));
    NOR2X1 U20082 (.A1(N1979), .A2(N33), .ZN(n32954));
    INVX1 U20083 (.I(n24437), .ZN(n32955));
    NOR2X1 U20084 (.A1(n22815), .A2(N8662), .ZN(N32956));
    NOR2X1 U20085 (.A1(n13138), .A2(n28566), .ZN(N32957));
    NOR2X1 U20086 (.A1(N11627), .A2(n17683), .ZN(N32958));
    INVX1 U20087 (.I(N10617), .ZN(n32959));
    NANDX1 U20088 (.A1(n26878), .A2(n28174), .ZN(N32960));
    NANDX1 U20089 (.A1(n29444), .A2(N9259), .ZN(n32961));
    NANDX1 U20090 (.A1(n15070), .A2(N1029), .ZN(n32962));
    NANDX1 U20091 (.A1(N646), .A2(N4719), .ZN(n32963));
    INVX1 U20092 (.I(n18392), .ZN(n32964));
    INVX1 U20093 (.I(N5985), .ZN(N32965));
    INVX1 U20094 (.I(n25215), .ZN(N32966));
    INVX1 U20095 (.I(N3231), .ZN(n32967));
    NANDX1 U20096 (.A1(n13754), .A2(N11892), .ZN(N32968));
    NANDX1 U20097 (.A1(n15452), .A2(n29018), .ZN(N32969));
    NANDX1 U20098 (.A1(n15639), .A2(n16563), .ZN(N32970));
    INVX1 U20099 (.I(n26256), .ZN(N32971));
    INVX1 U20100 (.I(N10376), .ZN(N32972));
    NOR2X1 U20101 (.A1(n17583), .A2(N9682), .ZN(N32973));
    INVX1 U20102 (.I(n13652), .ZN(n32974));
    NANDX1 U20103 (.A1(n23139), .A2(N12448), .ZN(n32975));
    NOR2X1 U20104 (.A1(n27858), .A2(N11010), .ZN(n32976));
    INVX1 U20105 (.I(N11464), .ZN(N32977));
    NOR2X1 U20106 (.A1(N11143), .A2(N6541), .ZN(N32978));
    INVX1 U20107 (.I(n14373), .ZN(N32979));
    NANDX1 U20108 (.A1(N10247), .A2(n26265), .ZN(N32980));
    NOR2X1 U20109 (.A1(n25699), .A2(n13706), .ZN(n32981));
    NOR2X1 U20110 (.A1(N11200), .A2(N132), .ZN(N32982));
    NOR2X1 U20111 (.A1(n26016), .A2(n19926), .ZN(N32983));
    NOR2X1 U20112 (.A1(n20170), .A2(n26069), .ZN(n32984));
    NANDX1 U20113 (.A1(N12144), .A2(n28282), .ZN(N32985));
    INVX1 U20114 (.I(N5145), .ZN(N32986));
    INVX1 U20115 (.I(N5918), .ZN(N32987));
    NANDX1 U20116 (.A1(n21601), .A2(N8129), .ZN(N32988));
    INVX1 U20117 (.I(n27156), .ZN(n32989));
    INVX1 U20118 (.I(n28127), .ZN(N32990));
    NANDX1 U20119 (.A1(n22205), .A2(N10415), .ZN(N32991));
    NANDX1 U20120 (.A1(N6893), .A2(n28981), .ZN(n32992));
    NANDX1 U20121 (.A1(n20599), .A2(n26953), .ZN(N32993));
    NOR2X1 U20122 (.A1(N9291), .A2(N8423), .ZN(N32994));
    NANDX1 U20123 (.A1(n29216), .A2(n18966), .ZN(N32995));
    NANDX1 U20124 (.A1(n13708), .A2(N9054), .ZN(n32996));
    NANDX1 U20125 (.A1(N11852), .A2(N12453), .ZN(n32997));
    INVX1 U20126 (.I(n22443), .ZN(N32998));
    NOR2X1 U20127 (.A1(n26920), .A2(n13907), .ZN(N32999));
    INVX1 U20128 (.I(n18370), .ZN(N33000));
    NANDX1 U20129 (.A1(n22891), .A2(N4920), .ZN(N33001));
    INVX1 U20130 (.I(N3520), .ZN(N33002));
    NOR2X1 U20131 (.A1(N4014), .A2(N10412), .ZN(n33003));
    NOR2X1 U20132 (.A1(N10592), .A2(N873), .ZN(n33004));
    INVX1 U20133 (.I(n16931), .ZN(N33005));
    INVX1 U20134 (.I(n19416), .ZN(N33006));
    INVX1 U20135 (.I(n27939), .ZN(N33007));
    NOR2X1 U20136 (.A1(n30095), .A2(N71), .ZN(n33008));
    NANDX1 U20137 (.A1(n23049), .A2(N11922), .ZN(N33009));
    NANDX1 U20138 (.A1(N9708), .A2(N4228), .ZN(N33010));
    INVX1 U20139 (.I(N6490), .ZN(n33011));
    INVX1 U20140 (.I(n28860), .ZN(N33012));
    INVX1 U20141 (.I(n24878), .ZN(N33013));
    INVX1 U20142 (.I(n18340), .ZN(n33014));
    NOR2X1 U20143 (.A1(n13693), .A2(N3536), .ZN(n33015));
    NOR2X1 U20144 (.A1(n24105), .A2(n17713), .ZN(N33016));
    NANDX1 U20145 (.A1(n13538), .A2(n28706), .ZN(n33017));
    NANDX1 U20146 (.A1(N12262), .A2(N6545), .ZN(N33018));
    NOR2X1 U20147 (.A1(n28761), .A2(N3349), .ZN(n33019));
    NOR2X1 U20148 (.A1(n28831), .A2(n27905), .ZN(N33020));
    NANDX1 U20149 (.A1(N10616), .A2(N4638), .ZN(N33021));
    INVX1 U20150 (.I(N3404), .ZN(N33022));
    NOR2X1 U20151 (.A1(N8987), .A2(n28796), .ZN(n33023));
    NANDX1 U20152 (.A1(n22407), .A2(N12097), .ZN(N33024));
    NANDX1 U20153 (.A1(N10609), .A2(n18531), .ZN(N33025));
    NANDX1 U20154 (.A1(N2705), .A2(n17540), .ZN(N33026));
    NANDX1 U20155 (.A1(n20418), .A2(n15702), .ZN(N33027));
    NANDX1 U20156 (.A1(n18986), .A2(N656), .ZN(N33028));
    NOR2X1 U20157 (.A1(n14091), .A2(N12017), .ZN(N33029));
    NANDX1 U20158 (.A1(N6000), .A2(n23335), .ZN(n33030));
    NANDX1 U20159 (.A1(N3767), .A2(n27564), .ZN(N33031));
    NOR2X1 U20160 (.A1(N8405), .A2(n30061), .ZN(N33032));
    NANDX1 U20161 (.A1(n26843), .A2(n27608), .ZN(n33033));
    INVX1 U20162 (.I(N2427), .ZN(N33034));
    NANDX1 U20163 (.A1(N6988), .A2(n18321), .ZN(N33035));
    INVX1 U20164 (.I(n14080), .ZN(N33036));
    NANDX1 U20165 (.A1(N10312), .A2(N1482), .ZN(N33037));
    INVX1 U20166 (.I(N592), .ZN(N33038));
    INVX1 U20167 (.I(n25402), .ZN(n33039));
    NOR2X1 U20168 (.A1(n25098), .A2(N3041), .ZN(N33040));
    INVX1 U20169 (.I(N6977), .ZN(n33041));
    INVX1 U20170 (.I(n16788), .ZN(n33042));
    NANDX1 U20171 (.A1(n21794), .A2(n20555), .ZN(n33043));
    NOR2X1 U20172 (.A1(n26063), .A2(n17520), .ZN(N33044));
    INVX1 U20173 (.I(N10858), .ZN(N33045));
    NANDX1 U20174 (.A1(N2252), .A2(N5749), .ZN(N33046));
    NOR2X1 U20175 (.A1(n29388), .A2(N1298), .ZN(N33047));
    NOR2X1 U20176 (.A1(n25555), .A2(n15377), .ZN(n33048));
    NANDX1 U20177 (.A1(N5729), .A2(N5419), .ZN(N33049));
    NANDX1 U20178 (.A1(n25018), .A2(N11163), .ZN(n33050));
    NANDX1 U20179 (.A1(n21716), .A2(n24821), .ZN(n33051));
    NANDX1 U20180 (.A1(N2367), .A2(n20358), .ZN(n33052));
    NANDX1 U20181 (.A1(n19155), .A2(n20531), .ZN(n33053));
    NOR2X1 U20182 (.A1(n28270), .A2(n25389), .ZN(N33054));
    INVX1 U20183 (.I(n15652), .ZN(N33055));
    NOR2X1 U20184 (.A1(n20177), .A2(n18437), .ZN(N33056));
    NANDX1 U20185 (.A1(n25925), .A2(N12209), .ZN(N33057));
    NOR2X1 U20186 (.A1(n15783), .A2(N5603), .ZN(N33058));
    NOR2X1 U20187 (.A1(N1022), .A2(N5329), .ZN(n33059));
    INVX1 U20188 (.I(N6441), .ZN(n33060));
    NOR2X1 U20189 (.A1(n23518), .A2(N6164), .ZN(N33061));
    INVX1 U20190 (.I(n15096), .ZN(n33062));
    NANDX1 U20191 (.A1(n16019), .A2(N6024), .ZN(N33063));
    NOR2X1 U20192 (.A1(n19059), .A2(n13739), .ZN(N33064));
    NANDX1 U20193 (.A1(n13754), .A2(N11871), .ZN(n33065));
    INVX1 U20194 (.I(n23073), .ZN(n33066));
    INVX1 U20195 (.I(n14139), .ZN(n33067));
    INVX1 U20196 (.I(n23080), .ZN(N33068));
    NANDX1 U20197 (.A1(n16159), .A2(N5151), .ZN(n33069));
    NOR2X1 U20198 (.A1(N1804), .A2(n29451), .ZN(n33070));
    NOR2X1 U20199 (.A1(N2826), .A2(n23341), .ZN(n33071));
    INVX1 U20200 (.I(n27964), .ZN(N33072));
    NANDX1 U20201 (.A1(N9865), .A2(n22688), .ZN(N33073));
    NOR2X1 U20202 (.A1(n13522), .A2(N12095), .ZN(n33074));
    NANDX1 U20203 (.A1(n19545), .A2(n21859), .ZN(N33075));
    INVX1 U20204 (.I(N3146), .ZN(n33076));
    NOR2X1 U20205 (.A1(N12061), .A2(N3577), .ZN(N33077));
    INVX1 U20206 (.I(n23695), .ZN(N33078));
    NANDX1 U20207 (.A1(N8684), .A2(n25367), .ZN(N33079));
    INVX1 U20208 (.I(N2227), .ZN(n33080));
    INVX1 U20209 (.I(n17751), .ZN(n33081));
    NANDX1 U20210 (.A1(n13192), .A2(N5625), .ZN(N33082));
    INVX1 U20211 (.I(N4578), .ZN(N33083));
    NANDX1 U20212 (.A1(n20335), .A2(n21102), .ZN(N33084));
    NOR2X1 U20213 (.A1(n18760), .A2(n13652), .ZN(N33085));
    INVX1 U20214 (.I(N2144), .ZN(n33086));
    NOR2X1 U20215 (.A1(N3768), .A2(N10249), .ZN(N33087));
    NOR2X1 U20216 (.A1(N2075), .A2(n13394), .ZN(N33088));
    NANDX1 U20217 (.A1(n14135), .A2(n16970), .ZN(n33089));
    NOR2X1 U20218 (.A1(N7692), .A2(N6491), .ZN(n33090));
    NOR2X1 U20219 (.A1(n21620), .A2(N7652), .ZN(N33091));
    NOR2X1 U20220 (.A1(N2870), .A2(n25402), .ZN(N33092));
    NANDX1 U20221 (.A1(N4622), .A2(n19588), .ZN(N33093));
    NOR2X1 U20222 (.A1(N9199), .A2(n18415), .ZN(n33094));
    NANDX1 U20223 (.A1(n18861), .A2(N3810), .ZN(n33095));
    INVX1 U20224 (.I(N2375), .ZN(N33096));
    NANDX1 U20225 (.A1(n25951), .A2(n16681), .ZN(n33097));
    INVX1 U20226 (.I(N6063), .ZN(N33098));
    NOR2X1 U20227 (.A1(n29989), .A2(N8017), .ZN(N33099));
    NANDX1 U20228 (.A1(N2547), .A2(n24987), .ZN(n33100));
    INVX1 U20229 (.I(N10239), .ZN(N33101));
    INVX1 U20230 (.I(n13095), .ZN(n33102));
    INVX1 U20231 (.I(n27690), .ZN(n33103));
    INVX1 U20232 (.I(n23288), .ZN(n33104));
    NANDX1 U20233 (.A1(n16017), .A2(n27910), .ZN(N33105));
    NANDX1 U20234 (.A1(n23608), .A2(n25669), .ZN(n33106));
    NOR2X1 U20235 (.A1(n28656), .A2(n14393), .ZN(N33107));
    INVX1 U20236 (.I(n22326), .ZN(N33108));
    INVX1 U20237 (.I(n17199), .ZN(N33109));
    NANDX1 U20238 (.A1(n22009), .A2(n14976), .ZN(N33110));
    NOR2X1 U20239 (.A1(n21838), .A2(N3388), .ZN(N33111));
    NOR2X1 U20240 (.A1(N8134), .A2(N5934), .ZN(N33112));
    NOR2X1 U20241 (.A1(N12836), .A2(n16172), .ZN(N33113));
    INVX1 U20242 (.I(n14492), .ZN(N33114));
    INVX1 U20243 (.I(n29037), .ZN(N33115));
    NOR2X1 U20244 (.A1(n29741), .A2(n29113), .ZN(N33116));
    NOR2X1 U20245 (.A1(n16074), .A2(n18638), .ZN(N33117));
    NANDX1 U20246 (.A1(N11605), .A2(n26578), .ZN(n33118));
    NOR2X1 U20247 (.A1(n14558), .A2(n26888), .ZN(N33119));
    NANDX1 U20248 (.A1(n19886), .A2(n13949), .ZN(N33120));
    NANDX1 U20249 (.A1(N318), .A2(n17485), .ZN(n33121));
    NANDX1 U20250 (.A1(n22155), .A2(n20872), .ZN(N33122));
    NANDX1 U20251 (.A1(n18849), .A2(n26806), .ZN(n33123));
    INVX1 U20252 (.I(n20246), .ZN(N33124));
    NANDX1 U20253 (.A1(n26977), .A2(N4600), .ZN(N33125));
    INVX1 U20254 (.I(n25876), .ZN(N33126));
    NANDX1 U20255 (.A1(n26155), .A2(n13412), .ZN(N33127));
    INVX1 U20256 (.I(N652), .ZN(n33128));
    NOR2X1 U20257 (.A1(N4367), .A2(N817), .ZN(N33129));
    INVX1 U20258 (.I(n16259), .ZN(n33130));
    INVX1 U20259 (.I(n13802), .ZN(N33131));
    INVX1 U20260 (.I(N5123), .ZN(N33132));
    NOR2X1 U20261 (.A1(N8239), .A2(N5440), .ZN(N33133));
    NOR2X1 U20262 (.A1(n20341), .A2(n16155), .ZN(n33134));
    NANDX1 U20263 (.A1(N11644), .A2(N4867), .ZN(n33135));
    INVX1 U20264 (.I(n25834), .ZN(N33136));
    INVX1 U20265 (.I(n29858), .ZN(n33137));
    NANDX1 U20266 (.A1(n18272), .A2(n26272), .ZN(N33138));
    INVX1 U20267 (.I(N8060), .ZN(n33139));
    NANDX1 U20268 (.A1(N8945), .A2(n29190), .ZN(n33140));
    INVX1 U20269 (.I(N10857), .ZN(N33141));
    NANDX1 U20270 (.A1(N12317), .A2(n16468), .ZN(N33142));
    INVX1 U20271 (.I(n16252), .ZN(N33143));
    NOR2X1 U20272 (.A1(N5698), .A2(n21374), .ZN(N33144));
    NOR2X1 U20273 (.A1(n13936), .A2(n15374), .ZN(N33145));
    NANDX1 U20274 (.A1(n22837), .A2(N1392), .ZN(N33146));
    INVX1 U20275 (.I(N4344), .ZN(n33147));
    NANDX1 U20276 (.A1(n15892), .A2(n18738), .ZN(n33148));
    NOR2X1 U20277 (.A1(n15612), .A2(n29971), .ZN(N33149));
    NANDX1 U20278 (.A1(N307), .A2(n25503), .ZN(N33150));
    NOR2X1 U20279 (.A1(n29854), .A2(N4310), .ZN(N33151));
    NOR2X1 U20280 (.A1(n29915), .A2(N3727), .ZN(N33152));
    NANDX1 U20281 (.A1(N655), .A2(n20195), .ZN(n33153));
    INVX1 U20282 (.I(n16907), .ZN(n33154));
    NANDX1 U20283 (.A1(n16909), .A2(n26841), .ZN(n33155));
    NANDX1 U20284 (.A1(n19405), .A2(N12078), .ZN(N33156));
    INVX1 U20285 (.I(N12105), .ZN(N33157));
    NANDX1 U20286 (.A1(N5806), .A2(N5009), .ZN(N33158));
    INVX1 U20287 (.I(n21697), .ZN(N33159));
    INVX1 U20288 (.I(N12597), .ZN(N33160));
    INVX1 U20289 (.I(N12140), .ZN(n33161));
    NOR2X1 U20290 (.A1(n26175), .A2(n26203), .ZN(N33162));
    NANDX1 U20291 (.A1(n14452), .A2(n19074), .ZN(N33163));
    NANDX1 U20292 (.A1(n14229), .A2(n22800), .ZN(N33164));
    NOR2X1 U20293 (.A1(N3444), .A2(N1418), .ZN(N33165));
    INVX1 U20294 (.I(n20350), .ZN(n33166));
    INVX1 U20295 (.I(N2975), .ZN(N33167));
    NANDX1 U20296 (.A1(N1316), .A2(N10941), .ZN(N33168));
    INVX1 U20297 (.I(N8248), .ZN(n33169));
    NANDX1 U20298 (.A1(N8282), .A2(n14053), .ZN(N33170));
    NOR2X1 U20299 (.A1(n23827), .A2(N5612), .ZN(N33171));
    NOR2X1 U20300 (.A1(n24984), .A2(N1343), .ZN(n33172));
    INVX1 U20301 (.I(n22765), .ZN(N33173));
    NOR2X1 U20302 (.A1(n25685), .A2(N2351), .ZN(N33174));
    NOR2X1 U20303 (.A1(n14621), .A2(N4370), .ZN(N33175));
    NOR2X1 U20304 (.A1(n25982), .A2(N9362), .ZN(n33176));
    INVX1 U20305 (.I(n27399), .ZN(N33177));
    INVX1 U20306 (.I(n15535), .ZN(N33178));
    NOR2X1 U20307 (.A1(n28540), .A2(n21149), .ZN(N33179));
    NOR2X1 U20308 (.A1(n28041), .A2(N8703), .ZN(N33180));
    NOR2X1 U20309 (.A1(n20948), .A2(N5545), .ZN(N33181));
    NOR2X1 U20310 (.A1(N7424), .A2(n17932), .ZN(N33182));
    INVX1 U20311 (.I(n24904), .ZN(N33183));
    NOR2X1 U20312 (.A1(N11076), .A2(n24386), .ZN(n33184));
    NOR2X1 U20313 (.A1(n27153), .A2(n19934), .ZN(N33185));
    INVX1 U20314 (.I(N4666), .ZN(N33186));
    INVX1 U20315 (.I(n19383), .ZN(n33187));
    NOR2X1 U20316 (.A1(n18959), .A2(n28744), .ZN(N33188));
    INVX1 U20317 (.I(N4782), .ZN(N33189));
    NOR2X1 U20318 (.A1(N7125), .A2(n19606), .ZN(N33190));
    INVX1 U20319 (.I(n28273), .ZN(N33191));
    NOR2X1 U20320 (.A1(N9039), .A2(n25536), .ZN(N33192));
    NOR2X1 U20321 (.A1(n18548), .A2(N943), .ZN(N33193));
    NANDX1 U20322 (.A1(n14532), .A2(n18874), .ZN(N33194));
    NANDX1 U20323 (.A1(N9299), .A2(n20212), .ZN(N33195));
    NOR2X1 U20324 (.A1(N3547), .A2(n14177), .ZN(N33196));
    INVX1 U20325 (.I(N12041), .ZN(N33197));
    NANDX1 U20326 (.A1(N7771), .A2(n23717), .ZN(N33198));
    NANDX1 U20327 (.A1(N4177), .A2(N1099), .ZN(n33199));
    NANDX1 U20328 (.A1(n25905), .A2(N5880), .ZN(n33200));
    NANDX1 U20329 (.A1(N2892), .A2(n25486), .ZN(n33201));
    NANDX1 U20330 (.A1(N1028), .A2(n19655), .ZN(N33202));
    NOR2X1 U20331 (.A1(n15124), .A2(N8075), .ZN(N33203));
    INVX1 U20332 (.I(n16067), .ZN(n33204));
    NANDX1 U20333 (.A1(N11313), .A2(n23501), .ZN(n33205));
    NANDX1 U20334 (.A1(N9172), .A2(N2137), .ZN(N33206));
    INVX1 U20335 (.I(N1280), .ZN(n33207));
    NANDX1 U20336 (.A1(n27706), .A2(N1881), .ZN(N33208));
    NANDX1 U20337 (.A1(n24037), .A2(n25597), .ZN(N33209));
    INVX1 U20338 (.I(n28214), .ZN(n33210));
    INVX1 U20339 (.I(n27963), .ZN(N33211));
    NANDX1 U20340 (.A1(n21136), .A2(n16161), .ZN(n33212));
    NANDX1 U20341 (.A1(N5045), .A2(n15493), .ZN(n33213));
    INVX1 U20342 (.I(n24700), .ZN(n33214));
    NOR2X1 U20343 (.A1(N8706), .A2(n21335), .ZN(N33215));
    INVX1 U20344 (.I(n24772), .ZN(N33216));
    INVX1 U20345 (.I(N9080), .ZN(N33217));
    NOR2X1 U20346 (.A1(N3063), .A2(n18251), .ZN(n33218));
    INVX1 U20347 (.I(n27663), .ZN(n33219));
    INVX1 U20348 (.I(n13706), .ZN(N33220));
    INVX1 U20349 (.I(N9972), .ZN(N33221));
    NANDX1 U20350 (.A1(N7691), .A2(n24129), .ZN(n33222));
    NANDX1 U20351 (.A1(n24465), .A2(N9248), .ZN(N33223));
    NANDX1 U20352 (.A1(N6869), .A2(n18945), .ZN(N33224));
    INVX1 U20353 (.I(N10863), .ZN(n33225));
    NOR2X1 U20354 (.A1(N5016), .A2(N4444), .ZN(N33226));
    NANDX1 U20355 (.A1(n17441), .A2(n13149), .ZN(N33227));
    INVX1 U20356 (.I(n26646), .ZN(n33228));
    INVX1 U20357 (.I(N1561), .ZN(N33229));
    NANDX1 U20358 (.A1(n21738), .A2(n23321), .ZN(n33230));
    INVX1 U20359 (.I(N432), .ZN(N33231));
    NOR2X1 U20360 (.A1(n20490), .A2(N2698), .ZN(N33232));
    NOR2X1 U20361 (.A1(N324), .A2(N8890), .ZN(N33233));
    NANDX1 U20362 (.A1(n24453), .A2(n26004), .ZN(N33234));
    INVX1 U20363 (.I(n22261), .ZN(n33235));
    INVX1 U20364 (.I(N9207), .ZN(N33236));
    NANDX1 U20365 (.A1(n19027), .A2(N8630), .ZN(n33237));
    NANDX1 U20366 (.A1(n24042), .A2(N1634), .ZN(N33238));
    INVX1 U20367 (.I(N11345), .ZN(n33239));
    NOR2X1 U20368 (.A1(n29038), .A2(n26552), .ZN(N33240));
    INVX1 U20369 (.I(n19159), .ZN(N33241));
    NOR2X1 U20370 (.A1(n21424), .A2(N12342), .ZN(N33242));
    INVX1 U20371 (.I(N10417), .ZN(n33243));
    NOR2X1 U20372 (.A1(n23452), .A2(n13114), .ZN(N33244));
    NANDX1 U20373 (.A1(N12336), .A2(N10565), .ZN(N33245));
    INVX1 U20374 (.I(n25349), .ZN(n33246));
    NANDX1 U20375 (.A1(N6459), .A2(n17473), .ZN(N33247));
    NANDX1 U20376 (.A1(N4226), .A2(n28540), .ZN(N33248));
    NANDX1 U20377 (.A1(N1416), .A2(n22020), .ZN(N33249));
    NOR2X1 U20378 (.A1(N3049), .A2(N11173), .ZN(N33250));
    NOR2X1 U20379 (.A1(N6392), .A2(N10073), .ZN(n33251));
    INVX1 U20380 (.I(N6079), .ZN(n33252));
    NOR2X1 U20381 (.A1(n24307), .A2(n16063), .ZN(N33253));
    NOR2X1 U20382 (.A1(n27269), .A2(n26479), .ZN(N33254));
    NANDX1 U20383 (.A1(N9144), .A2(n28154), .ZN(n33255));
    NANDX1 U20384 (.A1(n21479), .A2(N8581), .ZN(N33256));
    NANDX1 U20385 (.A1(N5252), .A2(n15011), .ZN(N33257));
    INVX1 U20386 (.I(N11285), .ZN(n33258));
    NANDX1 U20387 (.A1(N5600), .A2(n28385), .ZN(N33259));
    INVX1 U20388 (.I(N7015), .ZN(n33260));
    NANDX1 U20389 (.A1(n30038), .A2(N10064), .ZN(n33261));
    NOR2X1 U20390 (.A1(n25792), .A2(N5016), .ZN(N33262));
    NANDX1 U20391 (.A1(n29399), .A2(n29792), .ZN(N33263));
    INVX1 U20392 (.I(n23569), .ZN(N33264));
    NANDX1 U20393 (.A1(N6283), .A2(N9261), .ZN(N33265));
    NANDX1 U20394 (.A1(n28027), .A2(n18404), .ZN(N33266));
    NOR2X1 U20395 (.A1(n23003), .A2(n28443), .ZN(N33267));
    NANDX1 U20396 (.A1(n29358), .A2(N3557), .ZN(n33268));
    NANDX1 U20397 (.A1(N12035), .A2(N3402), .ZN(N33269));
    NOR2X1 U20398 (.A1(n17634), .A2(N1650), .ZN(n33270));
    NOR2X1 U20399 (.A1(n13210), .A2(N10478), .ZN(n33271));
    NOR2X1 U20400 (.A1(n23273), .A2(N341), .ZN(n33272));
    NOR2X1 U20401 (.A1(n16849), .A2(n18974), .ZN(n33273));
    NOR2X1 U20402 (.A1(n16504), .A2(n25261), .ZN(N33274));
    INVX1 U20403 (.I(N2084), .ZN(n33275));
    INVX1 U20404 (.I(n24793), .ZN(n33276));
    NANDX1 U20405 (.A1(n29432), .A2(n13059), .ZN(N33277));
    NOR2X1 U20406 (.A1(N10858), .A2(n30062), .ZN(n33278));
    INVX1 U20407 (.I(N10079), .ZN(N33279));
    NOR2X1 U20408 (.A1(n15161), .A2(N10674), .ZN(n33280));
    NOR2X1 U20409 (.A1(N12436), .A2(n28307), .ZN(n33281));
    NOR2X1 U20410 (.A1(n13764), .A2(N11379), .ZN(N33282));
    NANDX1 U20411 (.A1(N3553), .A2(n23212), .ZN(n33283));
    NOR2X1 U20412 (.A1(n19133), .A2(N9924), .ZN(N33284));
    NANDX1 U20413 (.A1(n22536), .A2(n14988), .ZN(N33285));
    NANDX1 U20414 (.A1(n19370), .A2(n17071), .ZN(n33286));
    NOR2X1 U20415 (.A1(n14025), .A2(N8334), .ZN(N33287));
    NOR2X1 U20416 (.A1(n15644), .A2(n16931), .ZN(N33288));
    INVX1 U20417 (.I(n15569), .ZN(N33289));
    NOR2X1 U20418 (.A1(n20764), .A2(n26309), .ZN(n33290));
    NOR2X1 U20419 (.A1(N1300), .A2(n21752), .ZN(N33291));
    NANDX1 U20420 (.A1(n18167), .A2(N7406), .ZN(N33292));
    NANDX1 U20421 (.A1(n18107), .A2(n14975), .ZN(N33293));
    INVX1 U20422 (.I(N11181), .ZN(N33294));
    NANDX1 U20423 (.A1(N2196), .A2(N9665), .ZN(N33295));
    INVX1 U20424 (.I(n24731), .ZN(n33296));
    NOR2X1 U20425 (.A1(n18758), .A2(n13964), .ZN(N33297));
    NOR2X1 U20426 (.A1(N593), .A2(n16549), .ZN(n33298));
    NOR2X1 U20427 (.A1(N420), .A2(N2056), .ZN(N33299));
    INVX1 U20428 (.I(N11105), .ZN(N33300));
    NANDX1 U20429 (.A1(N5138), .A2(N1731), .ZN(N33301));
    NANDX1 U20430 (.A1(N26), .A2(n21728), .ZN(N33302));
    NOR2X1 U20431 (.A1(N7350), .A2(N9758), .ZN(n33303));
    NOR2X1 U20432 (.A1(n28436), .A2(n16425), .ZN(N33304));
    NANDX1 U20433 (.A1(n22938), .A2(n27605), .ZN(N33305));
    NOR2X1 U20434 (.A1(n25133), .A2(n25831), .ZN(N33306));
    NOR2X1 U20435 (.A1(n19726), .A2(N8906), .ZN(N33307));
    NOR2X1 U20436 (.A1(n22250), .A2(n27750), .ZN(n33308));
    NOR2X1 U20437 (.A1(n27360), .A2(n13351), .ZN(N33309));
    NOR2X1 U20438 (.A1(n17976), .A2(n27321), .ZN(N33310));
    NOR2X1 U20439 (.A1(n24160), .A2(n21020), .ZN(N33311));
    NOR2X1 U20440 (.A1(N3637), .A2(n21045), .ZN(n33312));
    NANDX1 U20441 (.A1(n16304), .A2(n16955), .ZN(N33313));
    INVX1 U20442 (.I(n13499), .ZN(n33314));
    INVX1 U20443 (.I(n24985), .ZN(N33315));
    NOR2X1 U20444 (.A1(n26752), .A2(N11014), .ZN(N33316));
    NANDX1 U20445 (.A1(N10308), .A2(n25405), .ZN(N33317));
    NANDX1 U20446 (.A1(n18594), .A2(N4173), .ZN(N33318));
    NANDX1 U20447 (.A1(n29405), .A2(n20483), .ZN(N33319));
    NANDX1 U20448 (.A1(n26627), .A2(N3696), .ZN(N33320));
    INVX1 U20449 (.I(n14465), .ZN(N33321));
    NOR2X1 U20450 (.A1(N4919), .A2(n27185), .ZN(n33322));
    NOR2X1 U20451 (.A1(n23571), .A2(N684), .ZN(n33323));
    INVX1 U20452 (.I(n22374), .ZN(N33324));
    INVX1 U20453 (.I(N6883), .ZN(N33325));
    INVX1 U20454 (.I(n19046), .ZN(n33326));
    INVX1 U20455 (.I(N2904), .ZN(N33327));
    INVX1 U20456 (.I(N7311), .ZN(n33328));
    NANDX1 U20457 (.A1(N3583), .A2(N6179), .ZN(N33329));
    INVX1 U20458 (.I(n20215), .ZN(N33330));
    NOR2X1 U20459 (.A1(n20616), .A2(n15695), .ZN(N33331));
    INVX1 U20460 (.I(N10961), .ZN(N33332));
    INVX1 U20461 (.I(n20528), .ZN(n33333));
    INVX1 U20462 (.I(n23267), .ZN(n33334));
    NOR2X1 U20463 (.A1(n22795), .A2(n28185), .ZN(N33335));
    INVX1 U20464 (.I(n21815), .ZN(N33336));
    NANDX1 U20465 (.A1(n21283), .A2(N11742), .ZN(N33337));
    INVX1 U20466 (.I(n26831), .ZN(N33338));
    NOR2X1 U20467 (.A1(N10471), .A2(n15739), .ZN(N33339));
    INVX1 U20468 (.I(N1936), .ZN(N33340));
    INVX1 U20469 (.I(n13752), .ZN(N33341));
    NOR2X1 U20470 (.A1(n22458), .A2(N8491), .ZN(N33342));
    NANDX1 U20471 (.A1(N12535), .A2(N3126), .ZN(N33343));
    NOR2X1 U20472 (.A1(n16790), .A2(n15725), .ZN(N33344));
    NOR2X1 U20473 (.A1(n21923), .A2(N6116), .ZN(N33345));
    INVX1 U20474 (.I(N3613), .ZN(N33346));
    NANDX1 U20475 (.A1(n25427), .A2(N1660), .ZN(N33347));
    NOR2X1 U20476 (.A1(n17104), .A2(N11838), .ZN(N33348));
    NANDX1 U20477 (.A1(n17407), .A2(n21511), .ZN(N33349));
    NOR2X1 U20478 (.A1(n13152), .A2(N1845), .ZN(n33350));
    NANDX1 U20479 (.A1(n19594), .A2(N3780), .ZN(N33351));
    NOR2X1 U20480 (.A1(n21906), .A2(n26890), .ZN(N33352));
    INVX1 U20481 (.I(N260), .ZN(N33353));
    INVX1 U20482 (.I(N1682), .ZN(N33354));
    NANDX1 U20483 (.A1(n17502), .A2(N7032), .ZN(N33355));
    NANDX1 U20484 (.A1(n16918), .A2(n17515), .ZN(N33356));
    INVX1 U20485 (.I(n19550), .ZN(n33357));
    NANDX1 U20486 (.A1(n20575), .A2(N3401), .ZN(N33358));
    NOR2X1 U20487 (.A1(n29266), .A2(n20504), .ZN(N33359));
    NOR2X1 U20488 (.A1(n17663), .A2(n26471), .ZN(N33360));
    INVX1 U20489 (.I(N2754), .ZN(N33361));
    INVX1 U20490 (.I(N4963), .ZN(N33362));
    NOR2X1 U20491 (.A1(n17640), .A2(n27440), .ZN(N33363));
    NANDX1 U20492 (.A1(N9408), .A2(N12753), .ZN(N33364));
    NOR2X1 U20493 (.A1(n28365), .A2(n18922), .ZN(N33365));
    NANDX1 U20494 (.A1(n20310), .A2(N6286), .ZN(N33366));
    INVX1 U20495 (.I(n27980), .ZN(N33367));
    INVX1 U20496 (.I(n23041), .ZN(N33368));
    NOR2X1 U20497 (.A1(n19875), .A2(n14031), .ZN(N33369));
    NANDX1 U20498 (.A1(n23275), .A2(n25377), .ZN(n33370));
    INVX1 U20499 (.I(N2202), .ZN(n33371));
    NANDX1 U20500 (.A1(n14675), .A2(n28673), .ZN(N33372));
    NOR2X1 U20501 (.A1(N5989), .A2(n26719), .ZN(N33373));
    NANDX1 U20502 (.A1(n28269), .A2(n14221), .ZN(N33374));
    NANDX1 U20503 (.A1(n28677), .A2(N12189), .ZN(n33375));
    INVX1 U20504 (.I(N6792), .ZN(n33376));
    NOR2X1 U20505 (.A1(N2464), .A2(n16726), .ZN(N33377));
    NANDX1 U20506 (.A1(n27448), .A2(n22252), .ZN(N33378));
    INVX1 U20507 (.I(n27772), .ZN(N33379));
    INVX1 U20508 (.I(N5878), .ZN(N33380));
    NOR2X1 U20509 (.A1(n29185), .A2(N3761), .ZN(n33381));
    NANDX1 U20510 (.A1(n24425), .A2(n19471), .ZN(n33382));
    INVX1 U20511 (.I(N1272), .ZN(n33383));
    NOR2X1 U20512 (.A1(n18642), .A2(N11374), .ZN(N33384));
    NANDX1 U20513 (.A1(n15223), .A2(n14999), .ZN(N33385));
    INVX1 U20514 (.I(n18004), .ZN(N33386));
    NANDX1 U20515 (.A1(n25364), .A2(N55), .ZN(N33387));
    NOR2X1 U20516 (.A1(N2018), .A2(N10471), .ZN(N33388));
    NANDX1 U20517 (.A1(N7304), .A2(n29758), .ZN(n33389));
    INVX1 U20518 (.I(n29555), .ZN(n33390));
    NOR2X1 U20519 (.A1(N4135), .A2(n14573), .ZN(n33391));
    INVX1 U20520 (.I(n21644), .ZN(N33392));
    INVX1 U20521 (.I(N3509), .ZN(n33393));
    NANDX1 U20522 (.A1(N7907), .A2(N11540), .ZN(n33394));
    NANDX1 U20523 (.A1(n27876), .A2(n15547), .ZN(n33395));
    NANDX1 U20524 (.A1(n27810), .A2(n14103), .ZN(N33396));
    NOR2X1 U20525 (.A1(N12671), .A2(N10790), .ZN(n33397));
    NOR2X1 U20526 (.A1(n17157), .A2(n24714), .ZN(N33398));
    NOR2X1 U20527 (.A1(N5186), .A2(n26731), .ZN(n33399));
    NANDX1 U20528 (.A1(n14376), .A2(n22596), .ZN(N33400));
    INVX1 U20529 (.I(n20876), .ZN(N33401));
    NOR2X1 U20530 (.A1(N2247), .A2(n25010), .ZN(n33402));
    NOR2X1 U20531 (.A1(N1994), .A2(N5077), .ZN(n33403));
    INVX1 U20532 (.I(n24200), .ZN(N33404));
    INVX1 U20533 (.I(n16535), .ZN(N33405));
    NANDX1 U20534 (.A1(n25306), .A2(N2835), .ZN(N33406));
    INVX1 U20535 (.I(n24629), .ZN(N33407));
    NOR2X1 U20536 (.A1(n23811), .A2(n27734), .ZN(N33408));
    NANDX1 U20537 (.A1(N4463), .A2(n18706), .ZN(n33409));
    NANDX1 U20538 (.A1(n29176), .A2(n28430), .ZN(N33410));
    NANDX1 U20539 (.A1(n14331), .A2(N7048), .ZN(N33411));
    NOR2X1 U20540 (.A1(N6789), .A2(n15424), .ZN(n33412));
    NANDX1 U20541 (.A1(n28801), .A2(n17670), .ZN(N33413));
    INVX1 U20542 (.I(n23810), .ZN(N33414));
    NANDX1 U20543 (.A1(n13523), .A2(n13740), .ZN(N33415));
    NANDX1 U20544 (.A1(n28010), .A2(n18835), .ZN(N33416));
    INVX1 U20545 (.I(n23179), .ZN(n33417));
    NOR2X1 U20546 (.A1(N6158), .A2(N6231), .ZN(N33418));
    INVX1 U20547 (.I(n29968), .ZN(N33419));
    INVX1 U20548 (.I(N12475), .ZN(n33420));
    INVX1 U20549 (.I(N11093), .ZN(n33421));
    INVX1 U20550 (.I(n22030), .ZN(N33422));
    INVX1 U20551 (.I(N9693), .ZN(N33423));
    NANDX1 U20552 (.A1(n16433), .A2(n25269), .ZN(N33424));
    NANDX1 U20553 (.A1(n20417), .A2(N8706), .ZN(n33425));
    NOR2X1 U20554 (.A1(n26647), .A2(n17152), .ZN(n33426));
    NOR2X1 U20555 (.A1(N4733), .A2(n19235), .ZN(N33427));
    INVX1 U20556 (.I(n25717), .ZN(n33428));
    NANDX1 U20557 (.A1(N3603), .A2(n22166), .ZN(n33429));
    NOR2X1 U20558 (.A1(n13833), .A2(n16884), .ZN(n33430));
    NANDX1 U20559 (.A1(n24569), .A2(n16714), .ZN(N33431));
    NOR2X1 U20560 (.A1(n25604), .A2(N9568), .ZN(N33432));
    NOR2X1 U20561 (.A1(N3957), .A2(n20159), .ZN(N33433));
    NOR2X1 U20562 (.A1(n13649), .A2(n14942), .ZN(N33434));
    NANDX1 U20563 (.A1(n27479), .A2(N5075), .ZN(n33435));
    NANDX1 U20564 (.A1(N6047), .A2(N12569), .ZN(N33436));
    NANDX1 U20565 (.A1(N11759), .A2(n25174), .ZN(N33437));
    NANDX1 U20566 (.A1(N856), .A2(n28640), .ZN(n33438));
    NOR2X1 U20567 (.A1(N6524), .A2(N2105), .ZN(n33439));
    NANDX1 U20568 (.A1(N12492), .A2(n15937), .ZN(n33440));
    NANDX1 U20569 (.A1(N5992), .A2(n29066), .ZN(N33441));
    INVX1 U20570 (.I(n22017), .ZN(N33442));
    NOR2X1 U20571 (.A1(n18031), .A2(n18997), .ZN(N33443));
    INVX1 U20572 (.I(n26750), .ZN(n33444));
    NOR2X1 U20573 (.A1(n19259), .A2(N11555), .ZN(n33445));
    NANDX1 U20574 (.A1(n16600), .A2(N5190), .ZN(N33446));
    NOR2X1 U20575 (.A1(N11207), .A2(n17758), .ZN(N33447));
    NOR2X1 U20576 (.A1(n22965), .A2(N12794), .ZN(N33448));
    NANDX1 U20577 (.A1(N12382), .A2(N11296), .ZN(n33449));
    INVX1 U20578 (.I(N7466), .ZN(N33450));
    NOR2X1 U20579 (.A1(N4343), .A2(n19958), .ZN(N33451));
    INVX1 U20580 (.I(N7531), .ZN(N33452));
    INVX1 U20581 (.I(n24085), .ZN(N33453));
    NOR2X1 U20582 (.A1(n25087), .A2(N7041), .ZN(n33454));
    INVX1 U20583 (.I(n13946), .ZN(N33455));
    NOR2X1 U20584 (.A1(n19198), .A2(n16429), .ZN(n33456));
    NOR2X1 U20585 (.A1(N615), .A2(N11571), .ZN(N33457));
    INVX1 U20586 (.I(N5804), .ZN(N33458));
    NANDX1 U20587 (.A1(n18139), .A2(N12122), .ZN(n33459));
    NANDX1 U20588 (.A1(n29665), .A2(n24915), .ZN(n33460));
    INVX1 U20589 (.I(N11909), .ZN(n33461));
    INVX1 U20590 (.I(N10752), .ZN(N33462));
    NANDX1 U20591 (.A1(n15293), .A2(n15094), .ZN(N33463));
    NANDX1 U20592 (.A1(n21751), .A2(n22624), .ZN(N33464));
    NOR2X1 U20593 (.A1(N4259), .A2(n27179), .ZN(n33465));
    INVX1 U20594 (.I(N11299), .ZN(N33466));
    NANDX1 U20595 (.A1(n28419), .A2(N5251), .ZN(N33467));
    NANDX1 U20596 (.A1(n14710), .A2(N7023), .ZN(N33468));
    NOR2X1 U20597 (.A1(n26280), .A2(n13955), .ZN(N33469));
    INVX1 U20598 (.I(n23189), .ZN(n33470));
    NOR2X1 U20599 (.A1(N4349), .A2(n22282), .ZN(n33471));
    NOR2X1 U20600 (.A1(n17824), .A2(n14996), .ZN(n33472));
    INVX1 U20601 (.I(N1019), .ZN(n33473));
    INVX1 U20602 (.I(n28585), .ZN(N33474));
    NOR2X1 U20603 (.A1(N10703), .A2(n14900), .ZN(n33475));
    INVX1 U20604 (.I(n21888), .ZN(N33476));
    INVX1 U20605 (.I(n19441), .ZN(N33477));
    INVX1 U20606 (.I(N61), .ZN(n33478));
    INVX1 U20607 (.I(n27116), .ZN(N33479));
    NOR2X1 U20608 (.A1(n24551), .A2(n24363), .ZN(n33480));
    NOR2X1 U20609 (.A1(n20134), .A2(N10786), .ZN(N33481));
    NOR2X1 U20610 (.A1(N3951), .A2(n21711), .ZN(n33482));
    NANDX1 U20611 (.A1(n24605), .A2(n26059), .ZN(n33483));
    NOR2X1 U20612 (.A1(N3209), .A2(N2306), .ZN(n33484));
    NANDX1 U20613 (.A1(n23859), .A2(n22022), .ZN(N33485));
    NOR2X1 U20614 (.A1(n22306), .A2(n26893), .ZN(N33486));
    INVX1 U20615 (.I(N7068), .ZN(N33487));
    INVX1 U20616 (.I(N10525), .ZN(n33488));
    NOR2X1 U20617 (.A1(N1242), .A2(n18014), .ZN(N33489));
    NOR2X1 U20618 (.A1(N1844), .A2(N3553), .ZN(N33490));
    NANDX1 U20619 (.A1(n14955), .A2(n16476), .ZN(N33491));
    NANDX1 U20620 (.A1(N4952), .A2(n27262), .ZN(N33492));
    INVX1 U20621 (.I(n27600), .ZN(N33493));
    NANDX1 U20622 (.A1(n21700), .A2(N10628), .ZN(n33494));
    NOR2X1 U20623 (.A1(N469), .A2(n13837), .ZN(n33495));
    NOR2X1 U20624 (.A1(n24370), .A2(N7558), .ZN(N33496));
    NANDX1 U20625 (.A1(n13743), .A2(n18424), .ZN(N33497));
    INVX1 U20626 (.I(N2380), .ZN(n33498));
    NANDX1 U20627 (.A1(n13459), .A2(N1465), .ZN(n33499));
    NANDX1 U20628 (.A1(N3261), .A2(N8039), .ZN(N33500));
    INVX1 U20629 (.I(n23802), .ZN(N33501));
    NANDX1 U20630 (.A1(N816), .A2(N8619), .ZN(N33502));
    NANDX1 U20631 (.A1(N8001), .A2(N2131), .ZN(N33503));
    INVX1 U20632 (.I(n20198), .ZN(N33504));
    INVX1 U20633 (.I(n21147), .ZN(n33505));
    INVX1 U20634 (.I(n28919), .ZN(N33506));
    NOR2X1 U20635 (.A1(N790), .A2(N12618), .ZN(n33507));
    NOR2X1 U20636 (.A1(n25159), .A2(N8736), .ZN(N33508));
    INVX1 U20637 (.I(n27462), .ZN(N33509));
    NANDX1 U20638 (.A1(N2053), .A2(n29842), .ZN(N33510));
    NANDX1 U20639 (.A1(N4072), .A2(N1169), .ZN(N33511));
    INVX1 U20640 (.I(n26030), .ZN(n33512));
    NOR2X1 U20641 (.A1(N8842), .A2(n19694), .ZN(N33513));
    INVX1 U20642 (.I(N9657), .ZN(N33514));
    NOR2X1 U20643 (.A1(n25986), .A2(N6219), .ZN(N33515));
    NOR2X1 U20644 (.A1(n28298), .A2(n26416), .ZN(N33516));
    INVX1 U20645 (.I(N7868), .ZN(N33517));
    NOR2X1 U20646 (.A1(N5939), .A2(N9452), .ZN(N33518));
    NOR2X1 U20647 (.A1(N7118), .A2(N5219), .ZN(N33519));
    NANDX1 U20648 (.A1(N4414), .A2(n24448), .ZN(n33520));
    NANDX1 U20649 (.A1(N1436), .A2(n15061), .ZN(N33521));
    NANDX1 U20650 (.A1(N1070), .A2(n19132), .ZN(N33522));
    NANDX1 U20651 (.A1(n14669), .A2(N3585), .ZN(n33523));
    INVX1 U20652 (.I(n23510), .ZN(N33524));
    NANDX1 U20653 (.A1(n23691), .A2(n21728), .ZN(n33525));
    NANDX1 U20654 (.A1(N8100), .A2(n27946), .ZN(N33526));
    NANDX1 U20655 (.A1(n24959), .A2(n24224), .ZN(N33527));
    NANDX1 U20656 (.A1(n21387), .A2(N9385), .ZN(N33528));
    NANDX1 U20657 (.A1(N702), .A2(N6773), .ZN(N33529));
    INVX1 U20658 (.I(n24618), .ZN(N33530));
    NANDX1 U20659 (.A1(N7887), .A2(n18928), .ZN(N33531));
    INVX1 U20660 (.I(N9322), .ZN(N33532));
    NOR2X1 U20661 (.A1(N11571), .A2(n29089), .ZN(n33533));
    NOR2X1 U20662 (.A1(N9436), .A2(n13620), .ZN(N33534));
    NANDX1 U20663 (.A1(n23768), .A2(n25691), .ZN(n33535));
    NOR2X1 U20664 (.A1(N5882), .A2(n17281), .ZN(N33536));
    INVX1 U20665 (.I(n13981), .ZN(N33537));
    NOR2X1 U20666 (.A1(N8801), .A2(n27500), .ZN(N33538));
    NANDX1 U20667 (.A1(N10657), .A2(n18750), .ZN(N33539));
    NOR2X1 U20668 (.A1(n18452), .A2(N8012), .ZN(N33540));
    INVX1 U20669 (.I(n21924), .ZN(n33541));
    NOR2X1 U20670 (.A1(n27593), .A2(n29810), .ZN(n33542));
    NOR2X1 U20671 (.A1(N12329), .A2(n27692), .ZN(N33543));
    NOR2X1 U20672 (.A1(n23899), .A2(n15204), .ZN(n33544));
    INVX1 U20673 (.I(n21895), .ZN(n33545));
    INVX1 U20674 (.I(N6186), .ZN(N33546));
    NANDX1 U20675 (.A1(n12938), .A2(n21713), .ZN(N33547));
    INVX1 U20676 (.I(N81), .ZN(N33548));
    NOR2X1 U20677 (.A1(n23948), .A2(N3730), .ZN(n33549));
    NANDX1 U20678 (.A1(n21310), .A2(n20163), .ZN(N33550));
    INVX1 U20679 (.I(n28620), .ZN(N33551));
    NANDX1 U20680 (.A1(n20708), .A2(N6494), .ZN(N33552));
    NANDX1 U20681 (.A1(N1055), .A2(n27683), .ZN(N33553));
    INVX1 U20682 (.I(N728), .ZN(N33554));
    INVX1 U20683 (.I(N5202), .ZN(N33555));
    NANDX1 U20684 (.A1(n28615), .A2(n29100), .ZN(N33556));
    NOR2X1 U20685 (.A1(N974), .A2(n20857), .ZN(N33557));
    INVX1 U20686 (.I(n25857), .ZN(n33558));
    INVX1 U20687 (.I(N2231), .ZN(N33559));
    INVX1 U20688 (.I(N4772), .ZN(N33560));
    NANDX1 U20689 (.A1(N232), .A2(n28719), .ZN(N33561));
    INVX1 U20690 (.I(n21968), .ZN(N33562));
    NANDX1 U20691 (.A1(N3324), .A2(n24224), .ZN(N33563));
    NANDX1 U20692 (.A1(N7728), .A2(n14794), .ZN(N33564));
    NOR2X1 U20693 (.A1(N3146), .A2(N4410), .ZN(N33565));
    NOR2X1 U20694 (.A1(n26156), .A2(N5137), .ZN(n33566));
    INVX1 U20695 (.I(N1220), .ZN(n33567));
    INVX1 U20696 (.I(N5538), .ZN(N33568));
    NOR2X1 U20697 (.A1(N1284), .A2(n25209), .ZN(n33569));
    NANDX1 U20698 (.A1(n20714), .A2(N9490), .ZN(N33570));
    NANDX1 U20699 (.A1(N11505), .A2(n26922), .ZN(n33571));
    NOR2X1 U20700 (.A1(N2376), .A2(n15714), .ZN(n33572));
    NANDX1 U20701 (.A1(n27113), .A2(N7544), .ZN(N33573));
    NOR2X1 U20702 (.A1(n18998), .A2(n20329), .ZN(N33574));
    NANDX1 U20703 (.A1(n26725), .A2(n23683), .ZN(n33575));
    INVX1 U20704 (.I(n29871), .ZN(N33576));
    NANDX1 U20705 (.A1(n13229), .A2(n25889), .ZN(N33577));
    INVX1 U20706 (.I(n20288), .ZN(N33578));
    INVX1 U20707 (.I(N2329), .ZN(N33579));
    INVX1 U20708 (.I(n15851), .ZN(n33580));
    NANDX1 U20709 (.A1(n28156), .A2(n25450), .ZN(n33581));
    INVX1 U20710 (.I(N7508), .ZN(n33582));
    NOR2X1 U20711 (.A1(n24391), .A2(n22990), .ZN(N33583));
    NOR2X1 U20712 (.A1(n26767), .A2(n27264), .ZN(N33584));
    INVX1 U20713 (.I(N12303), .ZN(n33585));
    NOR2X1 U20714 (.A1(n17240), .A2(n19861), .ZN(N33586));
    NANDX1 U20715 (.A1(n17505), .A2(n16449), .ZN(N33587));
    INVX1 U20716 (.I(n19760), .ZN(N33588));
    NANDX1 U20717 (.A1(N5059), .A2(N2851), .ZN(n33589));
    NOR2X1 U20718 (.A1(n26848), .A2(N11699), .ZN(N33590));
    NOR2X1 U20719 (.A1(n17737), .A2(n14646), .ZN(n33591));
    INVX1 U20720 (.I(n21348), .ZN(n33592));
    NANDX1 U20721 (.A1(n23146), .A2(n22795), .ZN(N33593));
    NOR2X1 U20722 (.A1(N11424), .A2(n17049), .ZN(N33594));
    NOR2X1 U20723 (.A1(N8877), .A2(N2239), .ZN(n33595));
    INVX1 U20724 (.I(n21346), .ZN(n33596));
    NOR2X1 U20725 (.A1(N10638), .A2(n27146), .ZN(n33597));
    NOR2X1 U20726 (.A1(N12758), .A2(N3074), .ZN(n33598));
    NANDX1 U20727 (.A1(n19862), .A2(n22833), .ZN(N33599));
    INVX1 U20728 (.I(n24920), .ZN(n33600));
    INVX1 U20729 (.I(N10329), .ZN(n33601));
    INVX1 U20730 (.I(n25943), .ZN(n33602));
    INVX1 U20731 (.I(n27927), .ZN(n33603));
    NANDX1 U20732 (.A1(N12749), .A2(N7699), .ZN(n33604));
    NOR2X1 U20733 (.A1(N5757), .A2(N356), .ZN(n33605));
    NOR2X1 U20734 (.A1(n17180), .A2(N5965), .ZN(N33606));
    NOR2X1 U20735 (.A1(n14617), .A2(N8203), .ZN(n33607));
    NOR2X1 U20736 (.A1(n24523), .A2(N11305), .ZN(n33608));
    NOR2X1 U20737 (.A1(n21531), .A2(N4130), .ZN(N33609));
    NANDX1 U20738 (.A1(n13166), .A2(N1964), .ZN(N33610));
    INVX1 U20739 (.I(N5861), .ZN(N33611));
    INVX1 U20740 (.I(N8800), .ZN(n33612));
    NANDX1 U20741 (.A1(n14868), .A2(N7551), .ZN(N33613));
    INVX1 U20742 (.I(n18481), .ZN(N33614));
    NOR2X1 U20743 (.A1(n22180), .A2(N1092), .ZN(n33615));
    NOR2X1 U20744 (.A1(n22415), .A2(n25547), .ZN(N33616));
    NANDX1 U20745 (.A1(N8503), .A2(N12589), .ZN(n33617));
    NANDX1 U20746 (.A1(n14872), .A2(n27206), .ZN(N33618));
    NOR2X1 U20747 (.A1(n27209), .A2(N10152), .ZN(N33619));
    INVX1 U20748 (.I(n20046), .ZN(N33620));
    NANDX1 U20749 (.A1(N8677), .A2(n14202), .ZN(N33621));
    INVX1 U20750 (.I(N10640), .ZN(N33622));
    INVX1 U20751 (.I(N9132), .ZN(N33623));
    INVX1 U20752 (.I(N6880), .ZN(n33624));
    NOR2X1 U20753 (.A1(N7169), .A2(n14431), .ZN(N33625));
    INVX1 U20754 (.I(n25649), .ZN(N33626));
    INVX1 U20755 (.I(N2870), .ZN(N33627));
    NANDX1 U20756 (.A1(N9931), .A2(n25284), .ZN(N33628));
    NANDX1 U20757 (.A1(N446), .A2(n22347), .ZN(N33629));
    NOR2X1 U20758 (.A1(N8365), .A2(N7081), .ZN(N33630));
    NOR2X1 U20759 (.A1(N1609), .A2(N4152), .ZN(N33631));
    INVX1 U20760 (.I(N6156), .ZN(n33632));
    INVX1 U20761 (.I(n27884), .ZN(n33633));
    NANDX1 U20762 (.A1(n26960), .A2(N1018), .ZN(n33634));
    NANDX1 U20763 (.A1(n25040), .A2(n28847), .ZN(N33635));
    NOR2X1 U20764 (.A1(n20481), .A2(n16507), .ZN(n33636));
    NANDX1 U20765 (.A1(N4774), .A2(n15895), .ZN(N33637));
    NOR2X1 U20766 (.A1(N1666), .A2(n18765), .ZN(n33638));
    NANDX1 U20767 (.A1(N11596), .A2(N2472), .ZN(N33639));
    INVX1 U20768 (.I(N12041), .ZN(N33640));
    NANDX1 U20769 (.A1(n24006), .A2(N8967), .ZN(N33641));
    INVX1 U20770 (.I(n21494), .ZN(N33642));
    NOR2X1 U20771 (.A1(n24612), .A2(n17695), .ZN(N33643));
    NANDX1 U20772 (.A1(N7233), .A2(n15441), .ZN(n33644));
    NOR2X1 U20773 (.A1(n22753), .A2(N5019), .ZN(n33645));
    NOR2X1 U20774 (.A1(n17655), .A2(N3729), .ZN(N33646));
    NANDX1 U20775 (.A1(N7998), .A2(N8796), .ZN(N33647));
    INVX1 U20776 (.I(N1332), .ZN(n33648));
    INVX1 U20777 (.I(N2728), .ZN(n33649));
    NOR2X1 U20778 (.A1(n13317), .A2(N4164), .ZN(N33650));
    NOR2X1 U20779 (.A1(n15789), .A2(n16309), .ZN(N33651));
    NOR2X1 U20780 (.A1(n29168), .A2(N10177), .ZN(N33652));
    NANDX1 U20781 (.A1(n19490), .A2(n20232), .ZN(N33653));
    NANDX1 U20782 (.A1(n13964), .A2(N7789), .ZN(N33654));
    NOR2X1 U20783 (.A1(N9757), .A2(n23230), .ZN(N33655));
    INVX1 U20784 (.I(N2372), .ZN(N33656));
    INVX1 U20785 (.I(n29848), .ZN(N33657));
    NOR2X1 U20786 (.A1(n20537), .A2(n28760), .ZN(N33658));
    NOR2X1 U20787 (.A1(n17893), .A2(n22475), .ZN(N33659));
    NOR2X1 U20788 (.A1(N1007), .A2(n13763), .ZN(N33660));
    NANDX1 U20789 (.A1(n14323), .A2(n17926), .ZN(N33661));
    NOR2X1 U20790 (.A1(n18672), .A2(N4098), .ZN(n33662));
    NANDX1 U20791 (.A1(N6263), .A2(N2835), .ZN(N33663));
    INVX1 U20792 (.I(n25753), .ZN(n33664));
    INVX1 U20793 (.I(n22258), .ZN(n33665));
    INVX1 U20794 (.I(N718), .ZN(n33666));
    NANDX1 U20795 (.A1(N7897), .A2(N12508), .ZN(n33667));
    NOR2X1 U20796 (.A1(n28966), .A2(n29316), .ZN(n33668));
    NOR2X1 U20797 (.A1(N7416), .A2(n19716), .ZN(n33669));
    INVX1 U20798 (.I(N12562), .ZN(N33670));
    NANDX1 U20799 (.A1(n25764), .A2(n19039), .ZN(n33671));
    NANDX1 U20800 (.A1(n28088), .A2(n17073), .ZN(N33672));
    INVX1 U20801 (.I(n15876), .ZN(N33673));
    NOR2X1 U20802 (.A1(N7154), .A2(N8534), .ZN(N33674));
    NANDX1 U20803 (.A1(n13417), .A2(N11369), .ZN(N33675));
    NANDX1 U20804 (.A1(n27730), .A2(N4297), .ZN(n33676));
    INVX1 U20805 (.I(n25869), .ZN(N33677));
    NANDX1 U20806 (.A1(n16291), .A2(n22326), .ZN(N33678));
    NOR2X1 U20807 (.A1(N2550), .A2(n21155), .ZN(N33679));
    NOR2X1 U20808 (.A1(n25916), .A2(n17131), .ZN(N33680));
    NOR2X1 U20809 (.A1(n29205), .A2(n29692), .ZN(N33681));
    INVX1 U20810 (.I(n13393), .ZN(n33682));
    NANDX1 U20811 (.A1(N6606), .A2(N11343), .ZN(N33683));
    NOR2X1 U20812 (.A1(n25225), .A2(n15779), .ZN(N33684));
    NANDX1 U20813 (.A1(N2241), .A2(n24313), .ZN(N33685));
    INVX1 U20814 (.I(N4218), .ZN(n33686));
    NANDX1 U20815 (.A1(n20317), .A2(N1810), .ZN(N33687));
    NANDX1 U20816 (.A1(n15903), .A2(n27679), .ZN(n33688));
    NANDX1 U20817 (.A1(N2056), .A2(n19867), .ZN(N33689));
    NANDX1 U20818 (.A1(n23303), .A2(n29582), .ZN(n33690));
    INVX1 U20819 (.I(n19081), .ZN(N33691));
    NANDX1 U20820 (.A1(n16853), .A2(N6710), .ZN(N33692));
    NOR2X1 U20821 (.A1(n14982), .A2(n20102), .ZN(N33693));
    NANDX1 U20822 (.A1(N10148), .A2(n20005), .ZN(N33694));
    INVX1 U20823 (.I(N5235), .ZN(N33695));
    NANDX1 U20824 (.A1(n14102), .A2(n26173), .ZN(n33696));
    NOR2X1 U20825 (.A1(n19514), .A2(N254), .ZN(N33697));
    INVX1 U20826 (.I(n28392), .ZN(n33698));
    NOR2X1 U20827 (.A1(n29722), .A2(n14157), .ZN(n33699));
    NOR2X1 U20828 (.A1(N10258), .A2(N4773), .ZN(N33700));
    INVX1 U20829 (.I(N8314), .ZN(N33701));
    NANDX1 U20830 (.A1(N7476), .A2(N192), .ZN(n33702));
    INVX1 U20831 (.I(n24051), .ZN(N33703));
    NANDX1 U20832 (.A1(N850), .A2(n28742), .ZN(n33704));
    NOR2X1 U20833 (.A1(N9512), .A2(n29147), .ZN(N33705));
    INVX1 U20834 (.I(n29516), .ZN(N33706));
    NOR2X1 U20835 (.A1(N5830), .A2(n23722), .ZN(N33707));
    NANDX1 U20836 (.A1(N1866), .A2(N665), .ZN(N33708));
    NANDX1 U20837 (.A1(N2119), .A2(N1848), .ZN(N33709));
    INVX1 U20838 (.I(N4181), .ZN(N33710));
    NOR2X1 U20839 (.A1(n16651), .A2(n22483), .ZN(N33711));
    NANDX1 U20840 (.A1(N9984), .A2(N377), .ZN(N33712));
    NOR2X1 U20841 (.A1(n15180), .A2(n26550), .ZN(N33713));
    NOR2X1 U20842 (.A1(N9320), .A2(n20464), .ZN(N33714));
    INVX1 U20843 (.I(n28867), .ZN(n33715));
    INVX1 U20844 (.I(N4808), .ZN(n33716));
    NOR2X1 U20845 (.A1(N6638), .A2(N5403), .ZN(n33717));
    INVX1 U20846 (.I(n18839), .ZN(N33718));
    NOR2X1 U20847 (.A1(N8463), .A2(n15004), .ZN(n33719));
    INVX1 U20848 (.I(n27825), .ZN(N33720));
    INVX1 U20849 (.I(N3777), .ZN(N33721));
    INVX1 U20850 (.I(n21738), .ZN(N33722));
    NOR2X1 U20851 (.A1(n19665), .A2(N8251), .ZN(N33723));
    INVX1 U20852 (.I(N8475), .ZN(N33724));
    INVX1 U20853 (.I(N7937), .ZN(N33725));
    NOR2X1 U20854 (.A1(n21975), .A2(N4350), .ZN(N33726));
    NANDX1 U20855 (.A1(n19855), .A2(n13374), .ZN(N33727));
    INVX1 U20856 (.I(n18585), .ZN(n33728));
    NANDX1 U20857 (.A1(N10641), .A2(n15386), .ZN(N33729));
    INVX1 U20858 (.I(N4604), .ZN(N33730));
    NOR2X1 U20859 (.A1(n23599), .A2(N4397), .ZN(N33731));
    NANDX1 U20860 (.A1(N8465), .A2(N6055), .ZN(n33732));
    INVX1 U20861 (.I(n16270), .ZN(N33733));
    INVX1 U20862 (.I(n13069), .ZN(N33734));
    NOR2X1 U20863 (.A1(n25047), .A2(n21294), .ZN(N33735));
    NOR2X1 U20864 (.A1(N2470), .A2(n29769), .ZN(n33736));
    NOR2X1 U20865 (.A1(n29105), .A2(N5230), .ZN(n33737));
    NANDX1 U20866 (.A1(n22015), .A2(n26842), .ZN(N33738));
    NANDX1 U20867 (.A1(N5251), .A2(N2538), .ZN(n33739));
    NOR2X1 U20868 (.A1(n14813), .A2(n13178), .ZN(N33740));
    INVX1 U20869 (.I(N875), .ZN(N33741));
    NANDX1 U20870 (.A1(n22946), .A2(n24473), .ZN(N33742));
    INVX1 U20871 (.I(N8656), .ZN(N33743));
    NANDX1 U20872 (.A1(N5354), .A2(N3492), .ZN(n33744));
    NOR2X1 U20873 (.A1(N3746), .A2(N5122), .ZN(N33745));
    INVX1 U20874 (.I(n17353), .ZN(N33746));
    INVX1 U20875 (.I(N8742), .ZN(N33747));
    INVX1 U20876 (.I(n14607), .ZN(n33748));
    NANDX1 U20877 (.A1(N7350), .A2(N8398), .ZN(N33749));
    NANDX1 U20878 (.A1(n29364), .A2(N5102), .ZN(N33750));
    NOR2X1 U20879 (.A1(n23175), .A2(N7639), .ZN(N33751));
    NOR2X1 U20880 (.A1(n26548), .A2(N9377), .ZN(N33752));
    NOR2X1 U20881 (.A1(n15983), .A2(n15718), .ZN(N33753));
    NOR2X1 U20882 (.A1(n29016), .A2(n15017), .ZN(N33754));
    INVX1 U20883 (.I(n20377), .ZN(N33755));
    NANDX1 U20884 (.A1(N6013), .A2(n16567), .ZN(n33756));
    NOR2X1 U20885 (.A1(n29832), .A2(n20627), .ZN(N33757));
    INVX1 U20886 (.I(n26109), .ZN(N33758));
    INVX1 U20887 (.I(n26972), .ZN(N33759));
    NANDX1 U20888 (.A1(N8009), .A2(N4185), .ZN(n33760));
    NANDX1 U20889 (.A1(N8660), .A2(n22109), .ZN(N33761));
    NOR2X1 U20890 (.A1(N9600), .A2(N3708), .ZN(n33762));
    NOR2X1 U20891 (.A1(n29413), .A2(N118), .ZN(N33763));
    NANDX1 U20892 (.A1(N11771), .A2(n16101), .ZN(N33764));
    NOR2X1 U20893 (.A1(N5636), .A2(n14979), .ZN(N33765));
    NANDX1 U20894 (.A1(N8157), .A2(n23916), .ZN(N33766));
    INVX1 U20895 (.I(N2730), .ZN(N33767));
    NANDX1 U20896 (.A1(n28978), .A2(N2424), .ZN(n33768));
    INVX1 U20897 (.I(n17430), .ZN(N33769));
    NANDX1 U20898 (.A1(N7325), .A2(n14264), .ZN(n33770));
    NOR2X1 U20899 (.A1(N3894), .A2(N7009), .ZN(n33771));
    NANDX1 U20900 (.A1(N1114), .A2(n29118), .ZN(N33772));
    NANDX1 U20901 (.A1(N10713), .A2(N2688), .ZN(N33773));
    INVX1 U20902 (.I(n28686), .ZN(N33774));
    INVX1 U20903 (.I(n29136), .ZN(N33775));
    NANDX1 U20904 (.A1(n18905), .A2(n21490), .ZN(N33776));
    NOR2X1 U20905 (.A1(n22445), .A2(n28860), .ZN(N33777));
    NANDX1 U20906 (.A1(n16223), .A2(n15024), .ZN(N33778));
    NANDX1 U20907 (.A1(n15129), .A2(N2425), .ZN(N33779));
    NOR2X1 U20908 (.A1(N4525), .A2(n19854), .ZN(N33780));
    NANDX1 U20909 (.A1(N410), .A2(N3980), .ZN(n33781));
    NOR2X1 U20910 (.A1(N4303), .A2(N10989), .ZN(N33782));
    INVX1 U20911 (.I(N5416), .ZN(N33783));
    NOR2X1 U20912 (.A1(N8369), .A2(N4689), .ZN(N33784));
    INVX1 U20913 (.I(N594), .ZN(N33785));
    NANDX1 U20914 (.A1(n22719), .A2(n18291), .ZN(N33786));
    INVX1 U20915 (.I(N48), .ZN(N33787));
    INVX1 U20916 (.I(n21149), .ZN(N33788));
    NANDX1 U20917 (.A1(N8365), .A2(N10942), .ZN(N33789));
    INVX1 U20918 (.I(N11949), .ZN(n33790));
    NOR2X1 U20919 (.A1(N828), .A2(n14373), .ZN(n33791));
    NOR2X1 U20920 (.A1(n24050), .A2(n22787), .ZN(N33792));
    NANDX1 U20921 (.A1(n24459), .A2(n15327), .ZN(N33793));
    INVX1 U20922 (.I(n17322), .ZN(N33794));
    NANDX1 U20923 (.A1(N2319), .A2(N11298), .ZN(N33795));
    INVX1 U20924 (.I(N10687), .ZN(N33796));
    INVX1 U20925 (.I(N3182), .ZN(N33797));
    INVX1 U20926 (.I(n26481), .ZN(N33798));
    NOR2X1 U20927 (.A1(n18132), .A2(n24416), .ZN(N33799));
    INVX1 U20928 (.I(n27774), .ZN(N33800));
    NANDX1 U20929 (.A1(n14122), .A2(n24699), .ZN(N33801));
    NOR2X1 U20930 (.A1(N11259), .A2(n25208), .ZN(N33802));
    INVX1 U20931 (.I(N12086), .ZN(N33803));
    INVX1 U20932 (.I(N1183), .ZN(N33804));
    NANDX1 U20933 (.A1(n20790), .A2(n14708), .ZN(N33805));
    NANDX1 U20934 (.A1(N5979), .A2(N10746), .ZN(n33806));
    INVX1 U20935 (.I(N9416), .ZN(N33807));
    INVX1 U20936 (.I(n17498), .ZN(n33808));
    NANDX1 U20937 (.A1(N12312), .A2(n22044), .ZN(N33809));
    NOR2X1 U20938 (.A1(N12153), .A2(N6948), .ZN(n33810));
    NOR2X1 U20939 (.A1(n18845), .A2(N1227), .ZN(N33811));
    NOR2X1 U20940 (.A1(N5042), .A2(n16654), .ZN(N33812));
    INVX1 U20941 (.I(n18301), .ZN(N33813));
    NANDX1 U20942 (.A1(N4457), .A2(n13371), .ZN(N33814));
    NANDX1 U20943 (.A1(N5104), .A2(n30072), .ZN(N33815));
    NANDX1 U20944 (.A1(n29799), .A2(n20724), .ZN(n33816));
    NANDX1 U20945 (.A1(n18679), .A2(n15264), .ZN(n33817));
    NANDX1 U20946 (.A1(n24879), .A2(n13240), .ZN(N33818));
    NANDX1 U20947 (.A1(N801), .A2(n24620), .ZN(n33819));
    NANDX1 U20948 (.A1(n22844), .A2(n27743), .ZN(N33820));
    NOR2X1 U20949 (.A1(n18353), .A2(n15190), .ZN(N33821));
    INVX1 U20950 (.I(n19579), .ZN(N33822));
    NANDX1 U20951 (.A1(N1859), .A2(N6095), .ZN(n33823));
    NANDX1 U20952 (.A1(N8720), .A2(N7540), .ZN(N33824));
    NOR2X1 U20953 (.A1(N10652), .A2(n15940), .ZN(N33825));
    NANDX1 U20954 (.A1(N10586), .A2(n14083), .ZN(N33826));
    INVX1 U20955 (.I(N1173), .ZN(N33827));
    NOR2X1 U20956 (.A1(N3925), .A2(N4997), .ZN(N33828));
    INVX1 U20957 (.I(n17365), .ZN(N33829));
    NOR2X1 U20958 (.A1(n15476), .A2(N6726), .ZN(N33830));
    NANDX1 U20959 (.A1(n22872), .A2(n29569), .ZN(n33831));
    NOR2X1 U20960 (.A1(N844), .A2(N6345), .ZN(N33832));
    INVX1 U20961 (.I(n27797), .ZN(N33833));
    INVX1 U20962 (.I(N8341), .ZN(n33834));
    NOR2X1 U20963 (.A1(n20578), .A2(n25942), .ZN(N33835));
    INVX1 U20964 (.I(n16679), .ZN(N33836));
    INVX1 U20965 (.I(n26148), .ZN(N33837));
    NOR2X1 U20966 (.A1(N3448), .A2(N6596), .ZN(n33838));
    NOR2X1 U20967 (.A1(n18832), .A2(n26466), .ZN(N33839));
    NANDX1 U20968 (.A1(N11317), .A2(n20023), .ZN(n33840));
    NOR2X1 U20969 (.A1(n28681), .A2(n26819), .ZN(N33841));
    NANDX1 U20970 (.A1(N5269), .A2(n28098), .ZN(N33842));
    NOR2X1 U20971 (.A1(n23399), .A2(n26982), .ZN(n33843));
    INVX1 U20972 (.I(n29743), .ZN(N33844));
    NOR2X1 U20973 (.A1(N6145), .A2(n14090), .ZN(n33845));
    NANDX1 U20974 (.A1(n12921), .A2(N4530), .ZN(N33846));
    NANDX1 U20975 (.A1(n28417), .A2(N9769), .ZN(n33847));
    NANDX1 U20976 (.A1(n24427), .A2(N810), .ZN(N33848));
    NOR2X1 U20977 (.A1(n19584), .A2(N5933), .ZN(N33849));
    NOR2X1 U20978 (.A1(n15912), .A2(n26550), .ZN(N33850));
    INVX1 U20979 (.I(n24496), .ZN(N33851));
    INVX1 U20980 (.I(N610), .ZN(N33852));
    INVX1 U20981 (.I(n14932), .ZN(N33853));
    INVX1 U20982 (.I(n19137), .ZN(N33854));
    INVX1 U20983 (.I(n17837), .ZN(n33855));
    NOR2X1 U20984 (.A1(n23799), .A2(N6004), .ZN(N33856));
    NOR2X1 U20985 (.A1(n18504), .A2(N8654), .ZN(n33857));
    NANDX1 U20986 (.A1(N1288), .A2(n13183), .ZN(N33858));
    INVX1 U20987 (.I(n29704), .ZN(N33859));
    INVX1 U20988 (.I(n18250), .ZN(n33860));
    NOR2X1 U20989 (.A1(N12322), .A2(n20305), .ZN(N33861));
    INVX1 U20990 (.I(n18255), .ZN(N33862));
    NANDX1 U20991 (.A1(N6473), .A2(n14667), .ZN(N33863));
    NOR2X1 U20992 (.A1(N831), .A2(n21950), .ZN(N33864));
    NANDX1 U20993 (.A1(N10569), .A2(n25442), .ZN(n33865));
    INVX1 U20994 (.I(n29705), .ZN(N33866));
    INVX1 U20995 (.I(n14564), .ZN(N33867));
    INVX1 U20996 (.I(N11540), .ZN(n33868));
    NANDX1 U20997 (.A1(N871), .A2(n30043), .ZN(N33869));
    INVX1 U20998 (.I(n24148), .ZN(N33870));
    NOR2X1 U20999 (.A1(n19525), .A2(n20912), .ZN(N33871));
    INVX1 U21000 (.I(N900), .ZN(N33872));
    INVX1 U21001 (.I(n20573), .ZN(N33873));
    NOR2X1 U21002 (.A1(n17889), .A2(N11134), .ZN(n33874));
    NANDX1 U21003 (.A1(n28942), .A2(N6167), .ZN(N33875));
    NANDX1 U21004 (.A1(n23362), .A2(N6998), .ZN(N33876));
    NOR2X1 U21005 (.A1(N6953), .A2(N6127), .ZN(N33877));
    INVX1 U21006 (.I(N3680), .ZN(N33878));
    NOR2X1 U21007 (.A1(n28257), .A2(n18243), .ZN(N33879));
    INVX1 U21008 (.I(N9659), .ZN(N33880));
    NOR2X1 U21009 (.A1(N10673), .A2(N9565), .ZN(N33881));
    NOR2X1 U21010 (.A1(n23382), .A2(n29455), .ZN(N33882));
    NOR2X1 U21011 (.A1(N2717), .A2(n18775), .ZN(n33883));
    NOR2X1 U21012 (.A1(N301), .A2(N9210), .ZN(N33884));
    INVX1 U21013 (.I(N6750), .ZN(n33885));
    NOR2X1 U21014 (.A1(n27117), .A2(N5554), .ZN(n33886));
    NOR2X1 U21015 (.A1(N8804), .A2(n17476), .ZN(n33887));
    NANDX1 U21016 (.A1(N12439), .A2(n12989), .ZN(N33888));
    INVX1 U21017 (.I(N11379), .ZN(N33889));
    INVX1 U21018 (.I(n22448), .ZN(N33890));
    NANDX1 U21019 (.A1(N4774), .A2(N2114), .ZN(N33891));
    NANDX1 U21020 (.A1(N2007), .A2(N1347), .ZN(N33892));
    NANDX1 U21021 (.A1(N5581), .A2(n24728), .ZN(n33893));
    NANDX1 U21022 (.A1(N9982), .A2(n16005), .ZN(n33894));
    NANDX1 U21023 (.A1(N3842), .A2(n16305), .ZN(n33895));
    NANDX1 U21024 (.A1(n29621), .A2(N11615), .ZN(N33896));
    NANDX1 U21025 (.A1(n26601), .A2(n17168), .ZN(N33897));
    NANDX1 U21026 (.A1(N5267), .A2(n23205), .ZN(N33898));
    INVX1 U21027 (.I(n17705), .ZN(N33899));
    NANDX1 U21028 (.A1(N12787), .A2(n17645), .ZN(N33900));
    NOR2X1 U21029 (.A1(N5098), .A2(n27143), .ZN(N33901));
    NANDX1 U21030 (.A1(n25909), .A2(n23421), .ZN(n33902));
    NOR2X1 U21031 (.A1(n15816), .A2(n29264), .ZN(N33903));
    NOR2X1 U21032 (.A1(N10407), .A2(n22985), .ZN(N33904));
    INVX1 U21033 (.I(n14972), .ZN(N33905));
    NOR2X1 U21034 (.A1(n14589), .A2(N1140), .ZN(N33906));
    NANDX1 U21035 (.A1(n14072), .A2(N12754), .ZN(N33907));
    NANDX1 U21036 (.A1(n29233), .A2(n18483), .ZN(N33908));
    NOR2X1 U21037 (.A1(n23060), .A2(N11550), .ZN(N33909));
    NANDX1 U21038 (.A1(n29326), .A2(N6166), .ZN(n33910));
    NOR2X1 U21039 (.A1(n16833), .A2(n17450), .ZN(N33911));
    NOR2X1 U21040 (.A1(N2399), .A2(N3370), .ZN(n33912));
    NANDX1 U21041 (.A1(n25819), .A2(n28692), .ZN(n33913));
    INVX1 U21042 (.I(n13506), .ZN(N33914));
    NOR2X1 U21043 (.A1(N10336), .A2(N6353), .ZN(N33915));
    NOR2X1 U21044 (.A1(n25307), .A2(N257), .ZN(N33916));
    NANDX1 U21045 (.A1(n15007), .A2(n15865), .ZN(N33917));
    NOR2X1 U21046 (.A1(n16322), .A2(n20506), .ZN(n33918));
    INVX1 U21047 (.I(N4667), .ZN(N33919));
    INVX1 U21048 (.I(N7867), .ZN(n33920));
    NOR2X1 U21049 (.A1(N3889), .A2(N7055), .ZN(N33921));
    NANDX1 U21050 (.A1(N10012), .A2(N12448), .ZN(N33922));
    INVX1 U21051 (.I(n21233), .ZN(n33923));
    INVX1 U21052 (.I(N8883), .ZN(n33924));
    INVX1 U21053 (.I(n29225), .ZN(N33925));
    INVX1 U21054 (.I(n16714), .ZN(n33926));
    NOR2X1 U21055 (.A1(N6758), .A2(n27049), .ZN(N33927));
    NANDX1 U21056 (.A1(n16824), .A2(n22219), .ZN(N33928));
    NOR2X1 U21057 (.A1(n30040), .A2(n25786), .ZN(N33929));
    NANDX1 U21058 (.A1(n27190), .A2(N11970), .ZN(N33930));
    NANDX1 U21059 (.A1(N11996), .A2(n16636), .ZN(n33931));
    NANDX1 U21060 (.A1(N8423), .A2(N9973), .ZN(n33932));
    INVX1 U21061 (.I(N4038), .ZN(N33933));
    INVX1 U21062 (.I(n22828), .ZN(N33934));
    INVX1 U21063 (.I(n26428), .ZN(N33935));
    NANDX1 U21064 (.A1(n19891), .A2(n23871), .ZN(N33936));
    NANDX1 U21065 (.A1(N7540), .A2(N1171), .ZN(N33937));
    NOR2X1 U21066 (.A1(N8694), .A2(n26626), .ZN(n33938));
    INVX1 U21067 (.I(N4761), .ZN(n33939));
    INVX1 U21068 (.I(n20794), .ZN(N33940));
    NOR2X1 U21069 (.A1(n13215), .A2(n16443), .ZN(n33941));
    NANDX1 U21070 (.A1(n28965), .A2(n28412), .ZN(n33942));
    NOR2X1 U21071 (.A1(n29521), .A2(N3472), .ZN(N33943));
    NOR2X1 U21072 (.A1(N7807), .A2(N2005), .ZN(N33944));
    NOR2X1 U21073 (.A1(N405), .A2(N11480), .ZN(N33945));
    NANDX1 U21074 (.A1(N5451), .A2(n26468), .ZN(N33946));
    NOR2X1 U21075 (.A1(n13902), .A2(n20202), .ZN(N33947));
    NOR2X1 U21076 (.A1(N10002), .A2(N9933), .ZN(N33948));
    NANDX1 U21077 (.A1(n18695), .A2(N6422), .ZN(N33949));
    NOR2X1 U21078 (.A1(N12017), .A2(N8295), .ZN(N33950));
    NOR2X1 U21079 (.A1(N1662), .A2(N10070), .ZN(N33951));
    INVX1 U21080 (.I(N3495), .ZN(N33952));
    NOR2X1 U21081 (.A1(N11869), .A2(n15143), .ZN(N33953));
    NOR2X1 U21082 (.A1(n15340), .A2(n17021), .ZN(n33954));
    NANDX1 U21083 (.A1(n17345), .A2(n20276), .ZN(N33955));
    NOR2X1 U21084 (.A1(n17385), .A2(n27659), .ZN(N33956));
    NOR2X1 U21085 (.A1(n13716), .A2(n26087), .ZN(n33957));
    NANDX1 U21086 (.A1(n22478), .A2(N2206), .ZN(n33958));
    NOR2X1 U21087 (.A1(N2273), .A2(n21565), .ZN(n33959));
    INVX1 U21088 (.I(n27392), .ZN(N33960));
    NANDX1 U21089 (.A1(N661), .A2(n24247), .ZN(N33961));
    NANDX1 U21090 (.A1(n21020), .A2(N4179), .ZN(n33962));
    NOR2X1 U21091 (.A1(n13075), .A2(n24718), .ZN(N33963));
    INVX1 U21092 (.I(N9916), .ZN(n33964));
    NOR2X1 U21093 (.A1(N3662), .A2(n14562), .ZN(N33965));
    NANDX1 U21094 (.A1(n23937), .A2(n26872), .ZN(N33966));
    NOR2X1 U21095 (.A1(N10020), .A2(n25934), .ZN(N33967));
    INVX1 U21096 (.I(N5969), .ZN(N33968));
    NANDX1 U21097 (.A1(n27826), .A2(n26872), .ZN(N33969));
    INVX1 U21098 (.I(n18659), .ZN(N33970));
    NANDX1 U21099 (.A1(N4751), .A2(N4475), .ZN(N33971));
    INVX1 U21100 (.I(n24110), .ZN(N33972));
    INVX1 U21101 (.I(n15476), .ZN(N33973));
    NANDX1 U21102 (.A1(N2763), .A2(n28324), .ZN(N33974));
    NOR2X1 U21103 (.A1(N4398), .A2(n22904), .ZN(N33975));
    INVX1 U21104 (.I(n14313), .ZN(N33976));
    INVX1 U21105 (.I(n18369), .ZN(N33977));
    NOR2X1 U21106 (.A1(N7072), .A2(N730), .ZN(N33978));
    NANDX1 U21107 (.A1(n28842), .A2(N10749), .ZN(N33979));
    NANDX1 U21108 (.A1(n22751), .A2(N5278), .ZN(N33980));
    NOR2X1 U21109 (.A1(n20439), .A2(N2012), .ZN(n33981));
    INVX1 U21110 (.I(n27659), .ZN(n33982));
    NOR2X1 U21111 (.A1(n23964), .A2(N1996), .ZN(N33983));
    NOR2X1 U21112 (.A1(n17936), .A2(N579), .ZN(N33984));
    NOR2X1 U21113 (.A1(N2791), .A2(n22039), .ZN(N33985));
    NOR2X1 U21114 (.A1(n19418), .A2(n26437), .ZN(N33986));
    NOR2X1 U21115 (.A1(N3988), .A2(N10612), .ZN(N33987));
    NOR2X1 U21116 (.A1(N10917), .A2(n16608), .ZN(n33988));
    NOR2X1 U21117 (.A1(N207), .A2(n19339), .ZN(n33989));
    NANDX1 U21118 (.A1(n29653), .A2(n17866), .ZN(N33990));
    NANDX1 U21119 (.A1(N4793), .A2(n20973), .ZN(n33991));
    INVX1 U21120 (.I(n25502), .ZN(N33992));
    NANDX1 U21121 (.A1(N4798), .A2(N4235), .ZN(N33993));
    INVX1 U21122 (.I(N6793), .ZN(N33994));
    NANDX1 U21123 (.A1(n21811), .A2(n26070), .ZN(N33995));
    INVX1 U21124 (.I(n13162), .ZN(N33996));
    NANDX1 U21125 (.A1(n29671), .A2(N2442), .ZN(N33997));
    NOR2X1 U21126 (.A1(N916), .A2(n25127), .ZN(N33998));
    INVX1 U21127 (.I(n23681), .ZN(n33999));
    INVX1 U21128 (.I(n18611), .ZN(N34000));
    NOR2X1 U21129 (.A1(n13372), .A2(N7812), .ZN(N34001));
    NANDX1 U21130 (.A1(n12887), .A2(n25677), .ZN(N34002));
    NOR2X1 U21131 (.A1(N6241), .A2(N5073), .ZN(N34003));
    NOR2X1 U21132 (.A1(N1605), .A2(n15121), .ZN(N34004));
    INVX1 U21133 (.I(n24538), .ZN(N34005));
    NOR2X1 U21134 (.A1(N432), .A2(n23726), .ZN(N34006));
    NANDX1 U21135 (.A1(n26501), .A2(N3205), .ZN(n34007));
    NOR2X1 U21136 (.A1(N2896), .A2(N2739), .ZN(N34008));
    INVX1 U21137 (.I(N5726), .ZN(N34009));
    INVX1 U21138 (.I(n17080), .ZN(N34010));
    NANDX1 U21139 (.A1(N4456), .A2(N11546), .ZN(N34011));
    INVX1 U21140 (.I(N4959), .ZN(n34012));
    NOR2X1 U21141 (.A1(N4014), .A2(n29823), .ZN(n34013));
    NANDX1 U21142 (.A1(n18252), .A2(N4129), .ZN(n34014));
    INVX1 U21143 (.I(N11885), .ZN(n34015));
    NANDX1 U21144 (.A1(n22770), .A2(n27006), .ZN(N34016));
    NOR2X1 U21145 (.A1(n17170), .A2(N4425), .ZN(n34017));
    INVX1 U21146 (.I(n29456), .ZN(n34018));
    NANDX1 U21147 (.A1(n24980), .A2(N2524), .ZN(N34019));
    NANDX1 U21148 (.A1(n16436), .A2(n23960), .ZN(N34020));
    NANDX1 U21149 (.A1(n22162), .A2(N4735), .ZN(N34021));
    NOR2X1 U21150 (.A1(n29890), .A2(N9190), .ZN(n34022));
    NANDX1 U21151 (.A1(n26092), .A2(N2709), .ZN(N34023));
    NOR2X1 U21152 (.A1(n18667), .A2(N2394), .ZN(N34024));
    INVX1 U21153 (.I(N6781), .ZN(N34025));
    INVX1 U21154 (.I(N7217), .ZN(N34026));
    NANDX1 U21155 (.A1(n29629), .A2(n18547), .ZN(n34027));
    NANDX1 U21156 (.A1(n16237), .A2(N5580), .ZN(N34028));
    NOR2X1 U21157 (.A1(n14716), .A2(N4898), .ZN(n34029));
    INVX1 U21158 (.I(n28257), .ZN(n34030));
    NOR2X1 U21159 (.A1(n24034), .A2(n14555), .ZN(N34031));
    INVX1 U21160 (.I(n20591), .ZN(N34032));
    NANDX1 U21161 (.A1(n13236), .A2(N4090), .ZN(N34033));
    INVX1 U21162 (.I(N10987), .ZN(n34034));
    INVX1 U21163 (.I(n20984), .ZN(N34035));
    INVX1 U21164 (.I(n26355), .ZN(N34036));
    NANDX1 U21165 (.A1(N4650), .A2(N967), .ZN(N34037));
    NANDX1 U21166 (.A1(n29869), .A2(n26881), .ZN(n34038));
    INVX1 U21167 (.I(n17921), .ZN(N34039));
    INVX1 U21168 (.I(n16173), .ZN(N34040));
    INVX1 U21169 (.I(N9430), .ZN(n34041));
    NOR2X1 U21170 (.A1(N7297), .A2(N2889), .ZN(N34042));
    NOR2X1 U21171 (.A1(N5416), .A2(n29007), .ZN(N34043));
    INVX1 U21172 (.I(N8532), .ZN(N34044));
    NOR2X1 U21173 (.A1(N5592), .A2(N3671), .ZN(N34045));
    INVX1 U21174 (.I(N9682), .ZN(N34046));
    NOR2X1 U21175 (.A1(N8715), .A2(n27514), .ZN(N34047));
    NOR2X1 U21176 (.A1(N10971), .A2(n23731), .ZN(n34048));
    NANDX1 U21177 (.A1(n15620), .A2(n13258), .ZN(N34049));
    INVX1 U21178 (.I(N3912), .ZN(N34050));
    INVX1 U21179 (.I(n15855), .ZN(n34051));
    INVX1 U21180 (.I(n13851), .ZN(N34052));
    NOR2X1 U21181 (.A1(n14414), .A2(n23281), .ZN(N34053));
    NANDX1 U21182 (.A1(n21710), .A2(n26169), .ZN(N34054));
    NOR2X1 U21183 (.A1(n15687), .A2(n25038), .ZN(N34055));
    NOR2X1 U21184 (.A1(n24218), .A2(N9531), .ZN(n34056));
    NANDX1 U21185 (.A1(n27888), .A2(n18699), .ZN(N34057));
    NANDX1 U21186 (.A1(n26451), .A2(n15974), .ZN(N34058));
    NOR2X1 U21187 (.A1(n15860), .A2(n26944), .ZN(N34059));
    NANDX1 U21188 (.A1(n14781), .A2(N12426), .ZN(N34060));
    INVX1 U21189 (.I(N7117), .ZN(N34061));
    NANDX1 U21190 (.A1(N5126), .A2(n22971), .ZN(N34062));
    NOR2X1 U21191 (.A1(N7538), .A2(N1983), .ZN(N34063));
    INVX1 U21192 (.I(N681), .ZN(n34064));
    INVX1 U21193 (.I(N2579), .ZN(N34065));
    NANDX1 U21194 (.A1(n26447), .A2(N6826), .ZN(N34066));
    INVX1 U21195 (.I(n13513), .ZN(N34067));
    INVX1 U21196 (.I(n19841), .ZN(N34068));
    NOR2X1 U21197 (.A1(n17355), .A2(n27100), .ZN(n34069));
    NANDX1 U21198 (.A1(N2229), .A2(n12936), .ZN(N34070));
    NOR2X1 U21199 (.A1(n18088), .A2(N9743), .ZN(n34071));
    INVX1 U21200 (.I(n21429), .ZN(N34072));
    NANDX1 U21201 (.A1(n22614), .A2(n28546), .ZN(N34073));
    INVX1 U21202 (.I(n16300), .ZN(N34074));
    NANDX1 U21203 (.A1(N12220), .A2(n23837), .ZN(n34075));
    NANDX1 U21204 (.A1(n23226), .A2(n13078), .ZN(N34076));
    INVX1 U21205 (.I(n14366), .ZN(N34077));
    NANDX1 U21206 (.A1(N9735), .A2(N9752), .ZN(n34078));
    NOR2X1 U21207 (.A1(N11809), .A2(N10658), .ZN(n34079));
    NOR2X1 U21208 (.A1(n17979), .A2(n16573), .ZN(n34080));
    NANDX1 U21209 (.A1(n15048), .A2(n18801), .ZN(N34081));
    INVX1 U21210 (.I(n19091), .ZN(N34082));
    INVX1 U21211 (.I(N6563), .ZN(n34083));
    INVX1 U21212 (.I(N5301), .ZN(N34084));
    NOR2X1 U21213 (.A1(n27616), .A2(n22407), .ZN(N34085));
    NOR2X1 U21214 (.A1(N2339), .A2(n20908), .ZN(n34086));
    NOR2X1 U21215 (.A1(n14737), .A2(n21390), .ZN(n34087));
    NOR2X1 U21216 (.A1(n27814), .A2(N4678), .ZN(N34088));
    NOR2X1 U21217 (.A1(n26164), .A2(N2974), .ZN(n34089));
    NANDX1 U21218 (.A1(N4686), .A2(n14782), .ZN(N34090));
    NANDX1 U21219 (.A1(N3048), .A2(N2623), .ZN(n34091));
    NANDX1 U21220 (.A1(n17070), .A2(N6231), .ZN(N34092));
    NOR2X1 U21221 (.A1(n13890), .A2(n25322), .ZN(N34093));
    INVX1 U21222 (.I(N9014), .ZN(n34094));
    NOR2X1 U21223 (.A1(N10212), .A2(n14866), .ZN(N34095));
    NOR2X1 U21224 (.A1(N2482), .A2(N6207), .ZN(N34096));
    NOR2X1 U21225 (.A1(N11950), .A2(n28466), .ZN(N34097));
    NOR2X1 U21226 (.A1(N3202), .A2(n13677), .ZN(N34098));
    NANDX1 U21227 (.A1(N7880), .A2(N1813), .ZN(n34099));
    NOR2X1 U21228 (.A1(N10853), .A2(n29838), .ZN(N34100));
    NOR2X1 U21229 (.A1(n14195), .A2(n15505), .ZN(n34101));
    NOR2X1 U21230 (.A1(n16817), .A2(n29183), .ZN(N34102));
    NANDX1 U21231 (.A1(N11608), .A2(N8646), .ZN(N34103));
    NOR2X1 U21232 (.A1(n25490), .A2(n13557), .ZN(n34104));
    NOR2X1 U21233 (.A1(n14237), .A2(N12330), .ZN(N34105));
    INVX1 U21234 (.I(N462), .ZN(N34106));
    NANDX1 U21235 (.A1(n15842), .A2(N7724), .ZN(N34107));
    INVX1 U21236 (.I(n14170), .ZN(N34108));
    NANDX1 U21237 (.A1(n18522), .A2(n16407), .ZN(N34109));
    INVX1 U21238 (.I(n14962), .ZN(N34110));
    INVX1 U21239 (.I(N7900), .ZN(n34111));
    INVX1 U21240 (.I(N6481), .ZN(N34112));
    NOR2X1 U21241 (.A1(n28569), .A2(n21986), .ZN(n34113));
    NANDX1 U21242 (.A1(N3809), .A2(N9592), .ZN(N34114));
    NOR2X1 U21243 (.A1(n15417), .A2(n18238), .ZN(N34115));
    INVX1 U21244 (.I(n29467), .ZN(N34116));
    NANDX1 U21245 (.A1(N11369), .A2(n13567), .ZN(N34117));
    NANDX1 U21246 (.A1(n21004), .A2(n14028), .ZN(N34118));
    NOR2X1 U21247 (.A1(N6708), .A2(N10312), .ZN(N34119));
    NOR2X1 U21248 (.A1(N9438), .A2(n17155), .ZN(N34120));
    NOR2X1 U21249 (.A1(n25845), .A2(N2095), .ZN(N34121));
    NOR2X1 U21250 (.A1(N2488), .A2(n28693), .ZN(N34122));
    NANDX1 U21251 (.A1(n27666), .A2(n22660), .ZN(N34123));
    NANDX1 U21252 (.A1(N8075), .A2(n24441), .ZN(N34124));
    NOR2X1 U21253 (.A1(n17667), .A2(N2268), .ZN(N34125));
    INVX1 U21254 (.I(n24465), .ZN(n34126));
    INVX1 U21255 (.I(N10188), .ZN(N34127));
    NOR2X1 U21256 (.A1(N7358), .A2(N12315), .ZN(N34128));
    NANDX1 U21257 (.A1(n28361), .A2(n14904), .ZN(N34129));
    INVX1 U21258 (.I(n23629), .ZN(N34130));
    NANDX1 U21259 (.A1(n14247), .A2(n21627), .ZN(N34131));
    NOR2X1 U21260 (.A1(N991), .A2(n17334), .ZN(N34132));
    INVX1 U21261 (.I(n14135), .ZN(N34133));
    NANDX1 U21262 (.A1(n20141), .A2(N78), .ZN(n34134));
    INVX1 U21263 (.I(N12663), .ZN(N34135));
    INVX1 U21264 (.I(n13985), .ZN(N34136));
    NOR2X1 U21265 (.A1(n28730), .A2(n20212), .ZN(N34137));
    INVX1 U21266 (.I(N9451), .ZN(n34138));
    NOR2X1 U21267 (.A1(n23920), .A2(N8199), .ZN(n34139));
    NOR2X1 U21268 (.A1(n19838), .A2(n20514), .ZN(n34140));
    INVX1 U21269 (.I(n18061), .ZN(N34141));
    NANDX1 U21270 (.A1(n28018), .A2(N113), .ZN(N34142));
    INVX1 U21271 (.I(N688), .ZN(N34143));
    INVX1 U21272 (.I(N8409), .ZN(n34144));
    NOR2X1 U21273 (.A1(n27634), .A2(n29994), .ZN(N34145));
    INVX1 U21274 (.I(N5879), .ZN(N34146));
    NANDX1 U21275 (.A1(n23149), .A2(N350), .ZN(N34147));
    INVX1 U21276 (.I(n14860), .ZN(N34148));
    NOR2X1 U21277 (.A1(n28186), .A2(n13452), .ZN(N34149));
    NANDX1 U21278 (.A1(n14541), .A2(N11463), .ZN(N34150));
    NANDX1 U21279 (.A1(N8323), .A2(n19662), .ZN(N34151));
    INVX1 U21280 (.I(n28161), .ZN(n34152));
    INVX1 U21281 (.I(N11463), .ZN(N34153));
    NANDX1 U21282 (.A1(n22576), .A2(N9344), .ZN(n34154));
    NOR2X1 U21283 (.A1(N54), .A2(n28729), .ZN(N34155));
    NOR2X1 U21284 (.A1(N8462), .A2(N270), .ZN(N34156));
    NOR2X1 U21285 (.A1(N8318), .A2(N4643), .ZN(n34157));
    INVX1 U21286 (.I(n28314), .ZN(N34158));
    NOR2X1 U21287 (.A1(n26040), .A2(n19397), .ZN(n34159));
    NOR2X1 U21288 (.A1(N10237), .A2(N6006), .ZN(N34160));
    NANDX1 U21289 (.A1(N3206), .A2(n20546), .ZN(N34161));
    NOR2X1 U21290 (.A1(N10713), .A2(n28868), .ZN(n34162));
    NOR2X1 U21291 (.A1(N5865), .A2(n15452), .ZN(N34163));
    NOR2X1 U21292 (.A1(n17327), .A2(n20097), .ZN(n34164));
    NOR2X1 U21293 (.A1(n15231), .A2(N1976), .ZN(N34165));
    NOR2X1 U21294 (.A1(n13823), .A2(n17033), .ZN(N34166));
    NANDX1 U21295 (.A1(N2653), .A2(N6708), .ZN(n34167));
    NOR2X1 U21296 (.A1(n25993), .A2(N2262), .ZN(n34168));
    NANDX1 U21297 (.A1(N12207), .A2(n28301), .ZN(n34169));
    NOR2X1 U21298 (.A1(n13281), .A2(N8400), .ZN(N34170));
    NANDX1 U21299 (.A1(n16368), .A2(N166), .ZN(N34171));
    NOR2X1 U21300 (.A1(N12219), .A2(N10879), .ZN(n34172));
    INVX1 U21301 (.I(N4853), .ZN(n34173));
    INVX1 U21302 (.I(n24491), .ZN(N34174));
    INVX1 U21303 (.I(n22630), .ZN(n34175));
    NOR2X1 U21304 (.A1(N9892), .A2(n26422), .ZN(n34176));
    INVX1 U21305 (.I(n23752), .ZN(N34177));
    INVX1 U21306 (.I(N10579), .ZN(N34178));
    NANDX1 U21307 (.A1(N1320), .A2(N5847), .ZN(N34179));
    NANDX1 U21308 (.A1(n15873), .A2(N8108), .ZN(N34180));
    INVX1 U21309 (.I(n28079), .ZN(N34181));
    NANDX1 U21310 (.A1(n13395), .A2(n29921), .ZN(n34182));
    NANDX1 U21311 (.A1(n14597), .A2(n16151), .ZN(N34183));
    NANDX1 U21312 (.A1(n24905), .A2(n16930), .ZN(N34184));
    NOR2X1 U21313 (.A1(n22504), .A2(n21782), .ZN(N34185));
    NOR2X1 U21314 (.A1(N5418), .A2(n17866), .ZN(N34186));
    INVX1 U21315 (.I(N8428), .ZN(N34187));
    NANDX1 U21316 (.A1(n15614), .A2(N1974), .ZN(N34188));
    INVX1 U21317 (.I(n14281), .ZN(N34189));
    NOR2X1 U21318 (.A1(N2991), .A2(N4161), .ZN(n34190));
    NOR2X1 U21319 (.A1(n15250), .A2(n20033), .ZN(n34191));
    INVX1 U21320 (.I(n14749), .ZN(n34192));
    NANDX1 U21321 (.A1(n21338), .A2(n16704), .ZN(N34193));
    NOR2X1 U21322 (.A1(n13131), .A2(n19861), .ZN(n34194));
    NOR2X1 U21323 (.A1(n16528), .A2(n14628), .ZN(N34195));
    INVX1 U21324 (.I(n19364), .ZN(N34196));
    INVX1 U21325 (.I(n26862), .ZN(N34197));
    NANDX1 U21326 (.A1(N973), .A2(N3151), .ZN(N34198));
    NANDX1 U21327 (.A1(n28098), .A2(n19468), .ZN(N34199));
    NOR2X1 U21328 (.A1(n30072), .A2(n17960), .ZN(n34200));
    INVX1 U21329 (.I(n19745), .ZN(N34201));
    INVX1 U21330 (.I(n27872), .ZN(N34202));
    NOR2X1 U21331 (.A1(N6062), .A2(N6328), .ZN(n34203));
    NANDX1 U21332 (.A1(N9371), .A2(N1424), .ZN(n34204));
    INVX1 U21333 (.I(n26074), .ZN(N34205));
    NANDX1 U21334 (.A1(N11784), .A2(n15797), .ZN(N34206));
    INVX1 U21335 (.I(n28311), .ZN(n34207));
    NOR2X1 U21336 (.A1(N973), .A2(N6098), .ZN(n34208));
    INVX1 U21337 (.I(n16395), .ZN(N34209));
    INVX1 U21338 (.I(n15512), .ZN(N34210));
    NANDX1 U21339 (.A1(n27417), .A2(n13472), .ZN(n34211));
    INVX1 U21340 (.I(N6710), .ZN(N34212));
    NOR2X1 U21341 (.A1(n15396), .A2(N283), .ZN(n34213));
    INVX1 U21342 (.I(n24906), .ZN(N34214));
    NOR2X1 U21343 (.A1(n25537), .A2(n19529), .ZN(n34215));
    INVX1 U21344 (.I(n14292), .ZN(n34216));
    NOR2X1 U21345 (.A1(n13027), .A2(n12946), .ZN(N34217));
    INVX1 U21346 (.I(N9330), .ZN(N34218));
    NOR2X1 U21347 (.A1(n17754), .A2(n23920), .ZN(n34219));
    NANDX1 U21348 (.A1(N6602), .A2(n13454), .ZN(n34220));
    INVX1 U21349 (.I(N9702), .ZN(N34221));
    NOR2X1 U21350 (.A1(N9585), .A2(n25213), .ZN(n34222));
    NANDX1 U21351 (.A1(n25562), .A2(n27245), .ZN(N34223));
    NOR2X1 U21352 (.A1(n20832), .A2(n17773), .ZN(n34224));
    NANDX1 U21353 (.A1(n21114), .A2(n28045), .ZN(N34225));
    NANDX1 U21354 (.A1(n26390), .A2(N12005), .ZN(n34226));
    NOR2X1 U21355 (.A1(N7856), .A2(n14858), .ZN(n34227));
    NANDX1 U21356 (.A1(n20882), .A2(n27803), .ZN(N34228));
    NANDX1 U21357 (.A1(N74), .A2(N10955), .ZN(N34229));
    NOR2X1 U21358 (.A1(N12555), .A2(n22418), .ZN(n34230));
    NANDX1 U21359 (.A1(n26008), .A2(N9842), .ZN(N34231));
    NANDX1 U21360 (.A1(n14279), .A2(N7987), .ZN(N34232));
    INVX1 U21361 (.I(n22095), .ZN(N34233));
    NOR2X1 U21362 (.A1(N4705), .A2(N4469), .ZN(n34234));
    INVX1 U21363 (.I(N11038), .ZN(N34235));
    INVX1 U21364 (.I(n22477), .ZN(N34236));
    NOR2X1 U21365 (.A1(n13472), .A2(n18729), .ZN(N34237));
    NOR2X1 U21366 (.A1(n14098), .A2(n26584), .ZN(n34238));
    INVX1 U21367 (.I(N2047), .ZN(N34239));
    NANDX1 U21368 (.A1(N10594), .A2(N3391), .ZN(N34240));
    INVX1 U21369 (.I(n21548), .ZN(n34241));
    NOR2X1 U21370 (.A1(n18517), .A2(N2390), .ZN(N34242));
    NANDX1 U21371 (.A1(N2948), .A2(N792), .ZN(N34243));
    NOR2X1 U21372 (.A1(n17227), .A2(N8778), .ZN(N34244));
    INVX1 U21373 (.I(n27882), .ZN(N34245));
    NOR2X1 U21374 (.A1(N12738), .A2(N2213), .ZN(N34246));
    INVX1 U21375 (.I(n23775), .ZN(N34247));
    NOR2X1 U21376 (.A1(n24588), .A2(N9842), .ZN(N34248));
    NOR2X1 U21377 (.A1(n13180), .A2(n19352), .ZN(n34249));
    NANDX1 U21378 (.A1(N9626), .A2(N2143), .ZN(N34250));
    INVX1 U21379 (.I(n15515), .ZN(N34251));
    NOR2X1 U21380 (.A1(N3138), .A2(N10039), .ZN(N34252));
    NOR2X1 U21381 (.A1(n25627), .A2(n28555), .ZN(N34253));
    INVX1 U21382 (.I(N2101), .ZN(n34254));
    NOR2X1 U21383 (.A1(n14585), .A2(N2537), .ZN(n34255));
    NOR2X1 U21384 (.A1(N11923), .A2(N10569), .ZN(n34256));
    INVX1 U21385 (.I(N1232), .ZN(N34257));
    NOR2X1 U21386 (.A1(n25808), .A2(N3343), .ZN(n34258));
    NANDX1 U21387 (.A1(n18818), .A2(n16492), .ZN(N34259));
    NOR2X1 U21388 (.A1(n13860), .A2(n29671), .ZN(N34260));
    INVX1 U21389 (.I(N11561), .ZN(N34261));
    NOR2X1 U21390 (.A1(N2522), .A2(N11308), .ZN(n34262));
    NOR2X1 U21391 (.A1(N3818), .A2(n14446), .ZN(N34263));
    NOR2X1 U21392 (.A1(n15222), .A2(n28633), .ZN(n34264));
    NOR2X1 U21393 (.A1(n17577), .A2(n19294), .ZN(N34265));
    NOR2X1 U21394 (.A1(n20722), .A2(n21830), .ZN(N34266));
    NOR2X1 U21395 (.A1(N2508), .A2(n20960), .ZN(N34267));
    INVX1 U21396 (.I(n22437), .ZN(n34268));
    INVX1 U21397 (.I(n15155), .ZN(n34269));
    NANDX1 U21398 (.A1(n15452), .A2(N3835), .ZN(N34270));
    NOR2X1 U21399 (.A1(n19358), .A2(N6255), .ZN(N34271));
    NANDX1 U21400 (.A1(N1039), .A2(n17816), .ZN(n34272));
    NANDX1 U21401 (.A1(n22258), .A2(n17684), .ZN(n34273));
    INVX1 U21402 (.I(n26075), .ZN(N34274));
    INVX1 U21403 (.I(N136), .ZN(n34275));
    NANDX1 U21404 (.A1(n19185), .A2(n29085), .ZN(N34276));
    NANDX1 U21405 (.A1(N8342), .A2(n17822), .ZN(N34277));
    NANDX1 U21406 (.A1(n18732), .A2(N2273), .ZN(N34278));
    NANDX1 U21407 (.A1(n28252), .A2(n21757), .ZN(N34279));
    INVX1 U21408 (.I(n19502), .ZN(n34280));
    NOR2X1 U21409 (.A1(N12848), .A2(N4816), .ZN(N34281));
    NANDX1 U21410 (.A1(n13542), .A2(n24174), .ZN(N34282));
    INVX1 U21411 (.I(n13769), .ZN(n34283));
    INVX1 U21412 (.I(N11799), .ZN(N34284));
    NANDX1 U21413 (.A1(N5894), .A2(n18044), .ZN(N34285));
    NOR2X1 U21414 (.A1(n20529), .A2(N8596), .ZN(n34286));
    NOR2X1 U21415 (.A1(N8810), .A2(n16342), .ZN(N34287));
    INVX1 U21416 (.I(n14667), .ZN(n34288));
    INVX1 U21417 (.I(n20001), .ZN(N34289));
    NOR2X1 U21418 (.A1(N1838), .A2(n22273), .ZN(N34290));
    NANDX1 U21419 (.A1(n18651), .A2(n13892), .ZN(n34291));
    NANDX1 U21420 (.A1(N8015), .A2(n20665), .ZN(N34292));
    INVX1 U21421 (.I(N12830), .ZN(N34293));
    NOR2X1 U21422 (.A1(N635), .A2(n25564), .ZN(N34294));
    INVX1 U21423 (.I(N2964), .ZN(N34295));
    NOR2X1 U21424 (.A1(n14176), .A2(n21938), .ZN(N34296));
    NOR2X1 U21425 (.A1(N2082), .A2(n17775), .ZN(n34297));
    NOR2X1 U21426 (.A1(N10677), .A2(n13747), .ZN(N34298));
    NOR2X1 U21427 (.A1(n27018), .A2(n15926), .ZN(N34299));
    NOR2X1 U21428 (.A1(N10124), .A2(N5789), .ZN(N34300));
    NANDX1 U21429 (.A1(N523), .A2(n28061), .ZN(N34301));
    INVX1 U21430 (.I(n19173), .ZN(N34302));
    INVX1 U21431 (.I(n23270), .ZN(N34303));
    INVX1 U21432 (.I(n21040), .ZN(n34304));
    NANDX1 U21433 (.A1(n28577), .A2(n29433), .ZN(N34305));
    INVX1 U21434 (.I(N12565), .ZN(N34306));
    NOR2X1 U21435 (.A1(n13962), .A2(N10325), .ZN(N34307));
    NANDX1 U21436 (.A1(n24460), .A2(N2539), .ZN(n34308));
    NANDX1 U21437 (.A1(N12097), .A2(n15281), .ZN(N34309));
    NANDX1 U21438 (.A1(n14404), .A2(n25394), .ZN(N34310));
    NANDX1 U21439 (.A1(N192), .A2(n27296), .ZN(n34311));
    NOR2X1 U21440 (.A1(n24678), .A2(N10168), .ZN(N34312));
    NOR2X1 U21441 (.A1(n22601), .A2(n17615), .ZN(N34313));
    NANDX1 U21442 (.A1(n22976), .A2(n29446), .ZN(N34314));
    NOR2X1 U21443 (.A1(n13878), .A2(N9672), .ZN(n34315));
    NANDX1 U21444 (.A1(N1734), .A2(N9230), .ZN(N34316));
    NANDX1 U21445 (.A1(n14845), .A2(N11752), .ZN(n34317));
    INVX1 U21446 (.I(N554), .ZN(N34318));
    INVX1 U21447 (.I(n19022), .ZN(N34319));
    NOR2X1 U21448 (.A1(n18170), .A2(n22864), .ZN(n34320));
    INVX1 U21449 (.I(n21135), .ZN(N34321));
    INVX1 U21450 (.I(N857), .ZN(N34322));
    INVX1 U21451 (.I(N3839), .ZN(N34323));
    NANDX1 U21452 (.A1(n15867), .A2(N2568), .ZN(N34324));
    INVX1 U21453 (.I(n27028), .ZN(N34325));
    INVX1 U21454 (.I(n17687), .ZN(n34326));
    INVX1 U21455 (.I(N8051), .ZN(n34327));
    NANDX1 U21456 (.A1(n22305), .A2(N6283), .ZN(n34328));
    NANDX1 U21457 (.A1(n24039), .A2(N4074), .ZN(n34329));
    NOR2X1 U21458 (.A1(n27444), .A2(n15825), .ZN(N34330));
    NANDX1 U21459 (.A1(n27997), .A2(n21899), .ZN(N34331));
    INVX1 U21460 (.I(N4902), .ZN(n34332));
    INVX1 U21461 (.I(N10692), .ZN(n34333));
    NOR2X1 U21462 (.A1(n19626), .A2(n17373), .ZN(N34334));
    NOR2X1 U21463 (.A1(n29513), .A2(N9772), .ZN(n34335));
    NANDX1 U21464 (.A1(N3803), .A2(N12339), .ZN(N34336));
    NOR2X1 U21465 (.A1(N693), .A2(n21082), .ZN(N34337));
    NOR2X1 U21466 (.A1(N9120), .A2(n17693), .ZN(N34338));
    NANDX1 U21467 (.A1(N1288), .A2(n23976), .ZN(n34339));
    INVX1 U21468 (.I(n13887), .ZN(n34340));
    INVX1 U21469 (.I(n29544), .ZN(N34341));
    NOR2X1 U21470 (.A1(N2297), .A2(n28488), .ZN(n34342));
    NANDX1 U21471 (.A1(n24195), .A2(n16317), .ZN(N34343));
    NANDX1 U21472 (.A1(N11248), .A2(n15569), .ZN(N34344));
    NANDX1 U21473 (.A1(n19434), .A2(n21502), .ZN(N34345));
    NANDX1 U21474 (.A1(n18809), .A2(n19835), .ZN(N34346));
    INVX1 U21475 (.I(n22611), .ZN(N34347));
    NOR2X1 U21476 (.A1(N6147), .A2(n23304), .ZN(n34348));
    NOR2X1 U21477 (.A1(N11071), .A2(N2286), .ZN(n34349));
    NANDX1 U21478 (.A1(n21579), .A2(n22271), .ZN(N34350));
    NOR2X1 U21479 (.A1(n27086), .A2(n24718), .ZN(N34351));
    INVX1 U21480 (.I(n26493), .ZN(N34352));
    NANDX1 U21481 (.A1(N538), .A2(n24843), .ZN(n34353));
    NANDX1 U21482 (.A1(n13294), .A2(n29720), .ZN(n34354));
    INVX1 U21483 (.I(n13102), .ZN(N34355));
    NANDX1 U21484 (.A1(n14644), .A2(N2398), .ZN(N34356));
    NANDX1 U21485 (.A1(n15958), .A2(n21207), .ZN(n34357));
    NOR2X1 U21486 (.A1(N11988), .A2(N2241), .ZN(N34358));
    INVX1 U21487 (.I(N6695), .ZN(N34359));
    NOR2X1 U21488 (.A1(n17185), .A2(n17765), .ZN(n34360));
    NOR2X1 U21489 (.A1(N4979), .A2(n27905), .ZN(N34361));
    INVX1 U21490 (.I(n16748), .ZN(n34362));
    INVX1 U21491 (.I(n21803), .ZN(N34363));
    NANDX1 U21492 (.A1(n21208), .A2(N4697), .ZN(N34364));
    NANDX1 U21493 (.A1(N4475), .A2(n15341), .ZN(N34365));
    NANDX1 U21494 (.A1(N4057), .A2(n17060), .ZN(n34366));
    NANDX1 U21495 (.A1(N7769), .A2(n20265), .ZN(n34367));
    NOR2X1 U21496 (.A1(n21544), .A2(N6085), .ZN(n34368));
    NOR2X1 U21497 (.A1(n25015), .A2(N6633), .ZN(N34369));
    INVX1 U21498 (.I(N385), .ZN(n34370));
    NANDX1 U21499 (.A1(n17415), .A2(N6131), .ZN(N34371));
    NOR2X1 U21500 (.A1(n22366), .A2(N11109), .ZN(N34372));
    NANDX1 U21501 (.A1(n19451), .A2(n16418), .ZN(N34373));
    INVX1 U21502 (.I(n29814), .ZN(N34374));
    NOR2X1 U21503 (.A1(N10464), .A2(N4373), .ZN(N34375));
    NANDX1 U21504 (.A1(n14938), .A2(N8275), .ZN(N34376));
    NOR2X1 U21505 (.A1(N7556), .A2(n13895), .ZN(n34377));
    NANDX1 U21506 (.A1(N3885), .A2(N4022), .ZN(N34378));
    NANDX1 U21507 (.A1(n25428), .A2(n28804), .ZN(N34379));
    NANDX1 U21508 (.A1(n20306), .A2(N5299), .ZN(N34380));
    NANDX1 U21509 (.A1(N9251), .A2(n18625), .ZN(n34381));
    NOR2X1 U21510 (.A1(n15381), .A2(n26838), .ZN(n34382));
    INVX1 U21511 (.I(n15051), .ZN(n34383));
    INVX1 U21512 (.I(n16617), .ZN(N34384));
    NANDX1 U21513 (.A1(n14814), .A2(N4854), .ZN(n34385));
    INVX1 U21514 (.I(n13839), .ZN(N34386));
    NANDX1 U21515 (.A1(n29732), .A2(n28776), .ZN(n34387));
    NOR2X1 U21516 (.A1(n25409), .A2(N6194), .ZN(N34388));
    INVX1 U21517 (.I(N9992), .ZN(N34389));
    NANDX1 U21518 (.A1(N12539), .A2(N4575), .ZN(N34390));
    NANDX1 U21519 (.A1(N11205), .A2(N227), .ZN(n34391));
    NOR2X1 U21520 (.A1(N5065), .A2(n29327), .ZN(N34392));
    INVX1 U21521 (.I(n23689), .ZN(N34393));
    INVX1 U21522 (.I(n15988), .ZN(n34394));
    NANDX1 U21523 (.A1(N1294), .A2(n19599), .ZN(n34395));
    INVX1 U21524 (.I(N6472), .ZN(N34396));
    INVX1 U21525 (.I(n26443), .ZN(N34397));
    NOR2X1 U21526 (.A1(n26607), .A2(N10144), .ZN(n34398));
    INVX1 U21527 (.I(n14762), .ZN(N34399));
    NOR2X1 U21528 (.A1(N10993), .A2(N10033), .ZN(N34400));
    NANDX1 U21529 (.A1(n19510), .A2(N8585), .ZN(N34401));
    NOR2X1 U21530 (.A1(N1911), .A2(n13159), .ZN(n34402));
    NOR2X1 U21531 (.A1(N1676), .A2(n13386), .ZN(N34403));
    NANDX1 U21532 (.A1(N6740), .A2(N12575), .ZN(n34404));
    NOR2X1 U21533 (.A1(n18990), .A2(N5263), .ZN(N34405));
    NOR2X1 U21534 (.A1(n27939), .A2(n25254), .ZN(N34406));
    NANDX1 U21535 (.A1(N9431), .A2(N1588), .ZN(n34407));
    INVX1 U21536 (.I(n24435), .ZN(n34408));
    NOR2X1 U21537 (.A1(n13995), .A2(N4441), .ZN(N34409));
    INVX1 U21538 (.I(n28756), .ZN(N34410));
    NOR2X1 U21539 (.A1(n17398), .A2(n27349), .ZN(N34411));
    NANDX1 U21540 (.A1(N6770), .A2(n24495), .ZN(N34412));
    INVX1 U21541 (.I(n27378), .ZN(N34413));
    INVX1 U21542 (.I(N6680), .ZN(N34414));
    INVX1 U21543 (.I(n20901), .ZN(n34415));
    NOR2X1 U21544 (.A1(n24354), .A2(n22036), .ZN(N34416));
    NANDX1 U21545 (.A1(N1767), .A2(n15859), .ZN(N34417));
    INVX1 U21546 (.I(n18266), .ZN(N34418));
    NOR2X1 U21547 (.A1(N8820), .A2(n27697), .ZN(N34419));
    INVX1 U21548 (.I(n26345), .ZN(N34420));
    NANDX1 U21549 (.A1(n21295), .A2(N10202), .ZN(N34421));
    NANDX1 U21550 (.A1(n27700), .A2(n27518), .ZN(N34422));
    NANDX1 U21551 (.A1(n14960), .A2(n13290), .ZN(n34423));
    NOR2X1 U21552 (.A1(n21729), .A2(N7647), .ZN(N34424));
    INVX1 U21553 (.I(n18969), .ZN(N34425));
    NANDX1 U21554 (.A1(N5036), .A2(N6445), .ZN(N34426));
    NANDX1 U21555 (.A1(N6436), .A2(N661), .ZN(N34427));
    NOR2X1 U21556 (.A1(N3163), .A2(n21125), .ZN(n34428));
    NOR2X1 U21557 (.A1(N11206), .A2(N9254), .ZN(n34429));
    NANDX1 U21558 (.A1(N8586), .A2(n25511), .ZN(N34430));
    INVX1 U21559 (.I(N4793), .ZN(n34431));
    NOR2X1 U21560 (.A1(n24198), .A2(n14994), .ZN(N34432));
    INVX1 U21561 (.I(n21760), .ZN(N34433));
    INVX1 U21562 (.I(n14822), .ZN(n34434));
    INVX1 U21563 (.I(n14224), .ZN(N34435));
    NANDX1 U21564 (.A1(n28310), .A2(N10432), .ZN(N34436));
    INVX1 U21565 (.I(N5702), .ZN(N34437));
    INVX1 U21566 (.I(N5994), .ZN(n34438));
    INVX1 U21567 (.I(N8641), .ZN(N34439));
    NOR2X1 U21568 (.A1(N1368), .A2(n13724), .ZN(N34440));
    NANDX1 U21569 (.A1(n22493), .A2(N4529), .ZN(n34441));
    INVX1 U21570 (.I(n20307), .ZN(N34442));
    INVX1 U21571 (.I(N12503), .ZN(n34443));
    NOR2X1 U21572 (.A1(n27909), .A2(n17295), .ZN(n34444));
    NANDX1 U21573 (.A1(N10531), .A2(n20849), .ZN(N34445));
    NANDX1 U21574 (.A1(N2153), .A2(n21783), .ZN(N34446));
    NANDX1 U21575 (.A1(n27433), .A2(n24568), .ZN(N34447));
    INVX1 U21576 (.I(n14166), .ZN(N34448));
    NOR2X1 U21577 (.A1(N7895), .A2(n19868), .ZN(N34449));
    INVX1 U21578 (.I(N2449), .ZN(N34450));
    NOR2X1 U21579 (.A1(n27656), .A2(N3438), .ZN(N34451));
    INVX1 U21580 (.I(n29941), .ZN(n34452));
    NOR2X1 U21581 (.A1(n14297), .A2(n23030), .ZN(n34453));
    NOR2X1 U21582 (.A1(N4466), .A2(n17898), .ZN(N34454));
    NOR2X1 U21583 (.A1(N8706), .A2(N4231), .ZN(N34455));
    NOR2X1 U21584 (.A1(N175), .A2(n14761), .ZN(N34456));
    NANDX1 U21585 (.A1(N1127), .A2(N5474), .ZN(N34457));
    INVX1 U21586 (.I(n16900), .ZN(N34458));
    NOR2X1 U21587 (.A1(n13911), .A2(n23836), .ZN(N34459));
    NANDX1 U21588 (.A1(N7333), .A2(N1594), .ZN(N34460));
    INVX1 U21589 (.I(n26348), .ZN(N34461));
    INVX1 U21590 (.I(n27239), .ZN(N34462));
    NANDX1 U21591 (.A1(n26178), .A2(N7604), .ZN(N34463));
    NANDX1 U21592 (.A1(n22328), .A2(n21901), .ZN(n34464));
    NOR2X1 U21593 (.A1(N10956), .A2(n14927), .ZN(n34465));
    NANDX1 U21594 (.A1(n23526), .A2(N12194), .ZN(N34466));
    NANDX1 U21595 (.A1(N376), .A2(N929), .ZN(N34467));
    NANDX1 U21596 (.A1(N9513), .A2(N2055), .ZN(N34468));
    NOR2X1 U21597 (.A1(n17554), .A2(N7515), .ZN(N34469));
    NANDX1 U21598 (.A1(N1328), .A2(n19912), .ZN(N34470));
    NOR2X1 U21599 (.A1(N8660), .A2(N10066), .ZN(N34471));
    INVX1 U21600 (.I(n23569), .ZN(n34472));
    INVX1 U21601 (.I(n13756), .ZN(N34473));
    NANDX1 U21602 (.A1(n28845), .A2(n21360), .ZN(n34474));
    NOR2X1 U21603 (.A1(N9596), .A2(N1684), .ZN(n34475));
    NANDX1 U21604 (.A1(n20552), .A2(N5171), .ZN(n34476));
    NOR2X1 U21605 (.A1(n13940), .A2(n17364), .ZN(n34477));
    NOR2X1 U21606 (.A1(N2876), .A2(n18293), .ZN(N34478));
    INVX1 U21607 (.I(N949), .ZN(n34479));
    NANDX1 U21608 (.A1(N2826), .A2(n18503), .ZN(N34480));
    NANDX1 U21609 (.A1(N7322), .A2(N8391), .ZN(N34481));
    NOR2X1 U21610 (.A1(N10053), .A2(n17050), .ZN(n34482));
    NANDX1 U21611 (.A1(n26708), .A2(n29179), .ZN(n34483));
    NANDX1 U21612 (.A1(N10326), .A2(n23598), .ZN(N34484));
    NANDX1 U21613 (.A1(N1548), .A2(n18808), .ZN(n34485));
    INVX1 U21614 (.I(n21929), .ZN(n34486));
    NOR2X1 U21615 (.A1(n24905), .A2(n27100), .ZN(N34487));
    INVX1 U21616 (.I(n27406), .ZN(N34488));
    NANDX1 U21617 (.A1(n16099), .A2(N144), .ZN(n34489));
    NOR2X1 U21618 (.A1(n24456), .A2(N1093), .ZN(N34490));
    NOR2X1 U21619 (.A1(n15843), .A2(n19595), .ZN(n34491));
    INVX1 U21620 (.I(n23164), .ZN(n34492));
    INVX1 U21621 (.I(N6949), .ZN(N34493));
    NOR2X1 U21622 (.A1(N3458), .A2(N11771), .ZN(N34494));
    NOR2X1 U21623 (.A1(n21198), .A2(N7821), .ZN(N34495));
    NOR2X1 U21624 (.A1(n14658), .A2(N2579), .ZN(N34496));
    NANDX1 U21625 (.A1(n22027), .A2(n25631), .ZN(N34497));
    NOR2X1 U21626 (.A1(n18288), .A2(n20398), .ZN(N34498));
    INVX1 U21627 (.I(n22282), .ZN(N34499));
    NOR2X1 U21628 (.A1(n29119), .A2(n26941), .ZN(N34500));
    NANDX1 U21629 (.A1(N8722), .A2(N9821), .ZN(N34501));
    INVX1 U21630 (.I(n27369), .ZN(N34502));
    NOR2X1 U21631 (.A1(N4179), .A2(N9423), .ZN(N34503));
    NOR2X1 U21632 (.A1(n20724), .A2(n16371), .ZN(n34504));
    NOR2X1 U21633 (.A1(n24181), .A2(n16702), .ZN(N34505));
    NOR2X1 U21634 (.A1(N3802), .A2(n24522), .ZN(n34506));
    NOR2X1 U21635 (.A1(N7021), .A2(n15662), .ZN(n34507));
    INVX1 U21636 (.I(n29047), .ZN(N34508));
    NOR2X1 U21637 (.A1(n18065), .A2(N5758), .ZN(n34509));
    INVX1 U21638 (.I(n14160), .ZN(n34510));
    NANDX1 U21639 (.A1(n26340), .A2(N1703), .ZN(n34511));
    NANDX1 U21640 (.A1(n21271), .A2(n29122), .ZN(N34512));
    NOR2X1 U21641 (.A1(n17294), .A2(n14914), .ZN(n34513));
    NANDX1 U21642 (.A1(n21472), .A2(n24336), .ZN(N34514));
    NANDX1 U21643 (.A1(N12058), .A2(N10569), .ZN(n34515));
    NANDX1 U21644 (.A1(n24799), .A2(n27270), .ZN(n34516));
    NANDX1 U21645 (.A1(n17162), .A2(N10215), .ZN(N34517));
    INVX1 U21646 (.I(n24182), .ZN(n34518));
    NANDX1 U21647 (.A1(N12369), .A2(n23091), .ZN(N34519));
    INVX1 U21648 (.I(N297), .ZN(n34520));
    INVX1 U21649 (.I(N4128), .ZN(N34521));
    INVX1 U21650 (.I(n15311), .ZN(N34522));
    INVX1 U21651 (.I(n23417), .ZN(N34523));
    NANDX1 U21652 (.A1(N10161), .A2(N10962), .ZN(n34524));
    NANDX1 U21653 (.A1(n27454), .A2(n25875), .ZN(N34525));
    NANDX1 U21654 (.A1(N7349), .A2(n20073), .ZN(N34526));
    NOR2X1 U21655 (.A1(N7967), .A2(n19202), .ZN(N34527));
    NANDX1 U21656 (.A1(n21326), .A2(N4895), .ZN(N34528));
    INVX1 U21657 (.I(N8350), .ZN(n34529));
    NOR2X1 U21658 (.A1(n28220), .A2(N2394), .ZN(n34530));
    INVX1 U21659 (.I(N10452), .ZN(N34531));
    INVX1 U21660 (.I(N2122), .ZN(N34532));
    INVX1 U21661 (.I(N12756), .ZN(N34533));
    NANDX1 U21662 (.A1(N2325), .A2(n28066), .ZN(N34534));
    NANDX1 U21663 (.A1(n14303), .A2(n15204), .ZN(N34535));
    INVX1 U21664 (.I(n25264), .ZN(N34536));
    INVX1 U21665 (.I(n21313), .ZN(N34537));
    NOR2X1 U21666 (.A1(N1661), .A2(n17222), .ZN(n34538));
    INVX1 U21667 (.I(n15192), .ZN(N34539));
    NANDX1 U21668 (.A1(N7261), .A2(N595), .ZN(N34540));
    NANDX1 U21669 (.A1(N12155), .A2(n16679), .ZN(N34541));
    NOR2X1 U21670 (.A1(n15825), .A2(n14762), .ZN(N34542));
    INVX1 U21671 (.I(n22493), .ZN(n34543));
    INVX1 U21672 (.I(N11027), .ZN(N34544));
    NANDX1 U21673 (.A1(n13082), .A2(N12343), .ZN(N34545));
    NOR2X1 U21674 (.A1(N3967), .A2(n28969), .ZN(N34546));
    NANDX1 U21675 (.A1(N6830), .A2(n14036), .ZN(N34547));
    NOR2X1 U21676 (.A1(N1957), .A2(n16723), .ZN(N34548));
    NANDX1 U21677 (.A1(N11519), .A2(n18383), .ZN(N34549));
    NANDX1 U21678 (.A1(N11016), .A2(n22135), .ZN(n34550));
    NOR2X1 U21679 (.A1(N6837), .A2(n22729), .ZN(n34551));
    NANDX1 U21680 (.A1(N7553), .A2(N9271), .ZN(N34552));
    INVX1 U21681 (.I(N11938), .ZN(n34553));
    INVX1 U21682 (.I(n15631), .ZN(N34554));
    NANDX1 U21683 (.A1(n14927), .A2(n15218), .ZN(N34555));
    NOR2X1 U21684 (.A1(n16569), .A2(n27560), .ZN(N34556));
    NANDX1 U21685 (.A1(n20535), .A2(n26391), .ZN(N34557));
    INVX1 U21686 (.I(n27365), .ZN(N34558));
    NOR2X1 U21687 (.A1(N11033), .A2(n17882), .ZN(n34559));
    NOR2X1 U21688 (.A1(n29325), .A2(n29400), .ZN(N34560));
    INVX1 U21689 (.I(N4564), .ZN(N34561));
    INVX1 U21690 (.I(n25952), .ZN(n34562));
    NANDX1 U21691 (.A1(N5676), .A2(N7104), .ZN(N34563));
    NANDX1 U21692 (.A1(N1789), .A2(N4935), .ZN(N34564));
    NOR2X1 U21693 (.A1(n13726), .A2(n17527), .ZN(N34565));
    NANDX1 U21694 (.A1(n18019), .A2(n21014), .ZN(N34566));
    NANDX1 U21695 (.A1(n16787), .A2(N7445), .ZN(N34567));
    NOR2X1 U21696 (.A1(N4841), .A2(n27980), .ZN(N34568));
    INVX1 U21697 (.I(N7454), .ZN(N34569));
    NOR2X1 U21698 (.A1(n18056), .A2(N7048), .ZN(N34570));
    INVX1 U21699 (.I(n22189), .ZN(N34571));
    INVX1 U21700 (.I(n19472), .ZN(N34572));
    NANDX1 U21701 (.A1(N10799), .A2(N6871), .ZN(n34573));
    NOR2X1 U21702 (.A1(N4349), .A2(N1107), .ZN(N34574));
    INVX1 U21703 (.I(N3262), .ZN(n34575));
    INVX1 U21704 (.I(N10979), .ZN(N34576));
    INVX1 U21705 (.I(N5182), .ZN(N34577));
    NANDX1 U21706 (.A1(N12439), .A2(n23200), .ZN(N34578));
    NANDX1 U21707 (.A1(n19272), .A2(n28547), .ZN(N34579));
    NANDX1 U21708 (.A1(N12087), .A2(n21948), .ZN(N34580));
    NOR2X1 U21709 (.A1(N1156), .A2(n17963), .ZN(N34581));
    NOR2X1 U21710 (.A1(N7773), .A2(n25010), .ZN(n34582));
    NOR2X1 U21711 (.A1(n18522), .A2(n19805), .ZN(N34583));
    NANDX1 U21712 (.A1(N2950), .A2(N466), .ZN(n34584));
    NANDX1 U21713 (.A1(N1891), .A2(n23513), .ZN(N34585));
    NANDX1 U21714 (.A1(n26633), .A2(n15335), .ZN(N34586));
    NOR2X1 U21715 (.A1(n26172), .A2(N6021), .ZN(N34587));
    NANDX1 U21716 (.A1(N1662), .A2(N7021), .ZN(n34588));
    INVX1 U21717 (.I(n28303), .ZN(N34589));
    NANDX1 U21718 (.A1(n24265), .A2(n13553), .ZN(N34590));
    NOR2X1 U21719 (.A1(n16075), .A2(N3904), .ZN(N34591));
    NOR2X1 U21720 (.A1(n22598), .A2(n26720), .ZN(n34592));
    NOR2X1 U21721 (.A1(N6031), .A2(n20910), .ZN(N34593));
    NOR2X1 U21722 (.A1(n25836), .A2(N11693), .ZN(N34594));
    INVX1 U21723 (.I(n26301), .ZN(N34595));
    INVX1 U21724 (.I(n24910), .ZN(N34596));
    INVX1 U21725 (.I(n26804), .ZN(N34597));
    NOR2X1 U21726 (.A1(n23572), .A2(n17020), .ZN(N34598));
    NOR2X1 U21727 (.A1(n29592), .A2(N977), .ZN(N34599));
    NOR2X1 U21728 (.A1(n25173), .A2(N8134), .ZN(N34600));
    NOR2X1 U21729 (.A1(N9888), .A2(N2261), .ZN(n34601));
    NANDX1 U21730 (.A1(n25388), .A2(N6896), .ZN(N34602));
    INVX1 U21731 (.I(N467), .ZN(n34603));
    NOR2X1 U21732 (.A1(n15684), .A2(n13455), .ZN(N34604));
    INVX1 U21733 (.I(n25154), .ZN(N34605));
    INVX1 U21734 (.I(n19783), .ZN(N34606));
    NANDX1 U21735 (.A1(N7709), .A2(n15947), .ZN(n34607));
    INVX1 U21736 (.I(n21180), .ZN(N34608));
    INVX1 U21737 (.I(N1282), .ZN(n34609));
    NOR2X1 U21738 (.A1(n17617), .A2(N6862), .ZN(n34610));
    NANDX1 U21739 (.A1(N5633), .A2(N7839), .ZN(n34611));
    NANDX1 U21740 (.A1(n19366), .A2(n15972), .ZN(N34612));
    NANDX1 U21741 (.A1(n17815), .A2(N6793), .ZN(N34613));
    INVX1 U21742 (.I(N1626), .ZN(N34614));
    INVX1 U21743 (.I(N9040), .ZN(n34615));
    NANDX1 U21744 (.A1(n20303), .A2(n13285), .ZN(N34616));
    NOR2X1 U21745 (.A1(n14251), .A2(N8301), .ZN(n34617));
    INVX1 U21746 (.I(N3896), .ZN(N34618));
    NOR2X1 U21747 (.A1(n15202), .A2(N8403), .ZN(N34619));
    INVX1 U21748 (.I(n24942), .ZN(n34620));
    NANDX1 U21749 (.A1(n28165), .A2(n14511), .ZN(n34621));
    NANDX1 U21750 (.A1(N4890), .A2(n28777), .ZN(N34622));
    INVX1 U21751 (.I(N1289), .ZN(N34623));
    NOR2X1 U21752 (.A1(N10746), .A2(N5821), .ZN(N34624));
    NANDX1 U21753 (.A1(n17121), .A2(N12613), .ZN(N34625));
    NOR2X1 U21754 (.A1(n18746), .A2(N3422), .ZN(N34626));
    INVX1 U21755 (.I(N9398), .ZN(N34627));
    INVX1 U21756 (.I(N10648), .ZN(N34628));
    NANDX1 U21757 (.A1(n26536), .A2(N7510), .ZN(N34629));
    NANDX1 U21758 (.A1(N294), .A2(N11080), .ZN(N34630));
    NANDX1 U21759 (.A1(N8697), .A2(N7826), .ZN(N34631));
    NANDX1 U21760 (.A1(n18404), .A2(n24551), .ZN(n34632));
    NANDX1 U21761 (.A1(n15590), .A2(n18001), .ZN(N34633));
    NOR2X1 U21762 (.A1(N6970), .A2(n19289), .ZN(n34634));
    NOR2X1 U21763 (.A1(N6276), .A2(n25109), .ZN(n34635));
    NANDX1 U21764 (.A1(N11957), .A2(n26282), .ZN(N34636));
    INVX1 U21765 (.I(N565), .ZN(N34637));
    NOR2X1 U21766 (.A1(n25915), .A2(N9962), .ZN(N34638));
    INVX1 U21767 (.I(n25124), .ZN(n34639));
    NOR2X1 U21768 (.A1(N8250), .A2(N2496), .ZN(N34640));
    NANDX1 U21769 (.A1(n27241), .A2(n13575), .ZN(N34641));
    NOR2X1 U21770 (.A1(n24498), .A2(N9961), .ZN(N34642));
    NANDX1 U21771 (.A1(N12764), .A2(N4374), .ZN(N34643));
    NOR2X1 U21772 (.A1(n28354), .A2(n22375), .ZN(N34644));
    NOR2X1 U21773 (.A1(n23884), .A2(N87), .ZN(n34645));
    NANDX1 U21774 (.A1(n18720), .A2(n25196), .ZN(N34646));
    INVX1 U21775 (.I(N539), .ZN(N34647));
    NOR2X1 U21776 (.A1(n28170), .A2(n19801), .ZN(N34648));
    NOR2X1 U21777 (.A1(N12508), .A2(n29762), .ZN(N34649));
    NOR2X1 U21778 (.A1(N7494), .A2(N11650), .ZN(N34650));
    NOR2X1 U21779 (.A1(N9989), .A2(N3095), .ZN(n34651));
    INVX1 U21780 (.I(N12124), .ZN(n34652));
    INVX1 U21781 (.I(n28290), .ZN(N34653));
    NOR2X1 U21782 (.A1(N10410), .A2(n29615), .ZN(n34654));
    NOR2X1 U21783 (.A1(N1277), .A2(n16392), .ZN(N34655));
    NOR2X1 U21784 (.A1(n24857), .A2(N10138), .ZN(n34656));
    INVX1 U21785 (.I(n25824), .ZN(N34657));
    NOR2X1 U21786 (.A1(N9659), .A2(n25442), .ZN(n34658));
    INVX1 U21787 (.I(n19560), .ZN(N34659));
    NANDX1 U21788 (.A1(N7619), .A2(N6148), .ZN(N34660));
    NANDX1 U21789 (.A1(n25941), .A2(N4588), .ZN(n34661));
    NANDX1 U21790 (.A1(n26151), .A2(N11276), .ZN(N34662));
    INVX1 U21791 (.I(n29245), .ZN(N34663));
    NANDX1 U21792 (.A1(n19831), .A2(N11146), .ZN(n34664));
    NANDX1 U21793 (.A1(N11778), .A2(N10116), .ZN(N34665));
    NANDX1 U21794 (.A1(n15357), .A2(N11393), .ZN(n34666));
    NANDX1 U21795 (.A1(N11173), .A2(n24810), .ZN(N34667));
    INVX1 U21796 (.I(n25773), .ZN(n34668));
    NOR2X1 U21797 (.A1(n22326), .A2(n23993), .ZN(n34669));
    INVX1 U21798 (.I(n28842), .ZN(N34670));
    NANDX1 U21799 (.A1(N4958), .A2(N6323), .ZN(N34671));
    NOR2X1 U21800 (.A1(n18061), .A2(N2126), .ZN(N34672));
    INVX1 U21801 (.I(n27218), .ZN(N34673));
    NANDX1 U21802 (.A1(N12547), .A2(n16227), .ZN(N34674));
    INVX1 U21803 (.I(n16175), .ZN(N34675));
    INVX1 U21804 (.I(n15650), .ZN(n34676));
    NOR2X1 U21805 (.A1(N6259), .A2(n25766), .ZN(N34677));
    NANDX1 U21806 (.A1(N10176), .A2(n25719), .ZN(N34678));
    NOR2X1 U21807 (.A1(N9909), .A2(n20391), .ZN(N34679));
    INVX1 U21808 (.I(N5544), .ZN(N34680));
    NANDX1 U21809 (.A1(N2721), .A2(n29536), .ZN(N34681));
    NOR2X1 U21810 (.A1(N1425), .A2(N1374), .ZN(N34682));
    INVX1 U21811 (.I(N7747), .ZN(N34683));
    NANDX1 U21812 (.A1(n15251), .A2(n28570), .ZN(n34684));
    NOR2X1 U21813 (.A1(N12331), .A2(n15269), .ZN(N34685));
    NANDX1 U21814 (.A1(n17119), .A2(N1075), .ZN(N34686));
    INVX1 U21815 (.I(N11600), .ZN(N34687));
    NOR2X1 U21816 (.A1(N11687), .A2(N6419), .ZN(N34688));
    INVX1 U21817 (.I(n15282), .ZN(N34689));
    NOR2X1 U21818 (.A1(n26632), .A2(N2208), .ZN(n34690));
    NANDX1 U21819 (.A1(N5446), .A2(n24180), .ZN(n34691));
    INVX1 U21820 (.I(N4757), .ZN(n34692));
    NOR2X1 U21821 (.A1(N8566), .A2(n27127), .ZN(N34693));
    NOR2X1 U21822 (.A1(n28637), .A2(n24317), .ZN(n34694));
    INVX1 U21823 (.I(n26694), .ZN(n34695));
    INVX1 U21824 (.I(N11626), .ZN(n34696));
    NOR2X1 U21825 (.A1(N10321), .A2(n26894), .ZN(N34697));
    NANDX1 U21826 (.A1(n16000), .A2(n16530), .ZN(N34698));
    NANDX1 U21827 (.A1(n27599), .A2(n21815), .ZN(N34699));
    NOR2X1 U21828 (.A1(N3880), .A2(n22728), .ZN(n34700));
    NOR2X1 U21829 (.A1(N9034), .A2(N7783), .ZN(N34701));
    NANDX1 U21830 (.A1(n24096), .A2(N1789), .ZN(n34702));
    NOR2X1 U21831 (.A1(n14565), .A2(n25243), .ZN(N34703));
    NOR2X1 U21832 (.A1(N11691), .A2(N10793), .ZN(N34704));
    NOR2X1 U21833 (.A1(N10190), .A2(n23670), .ZN(N34705));
    NOR2X1 U21834 (.A1(n25445), .A2(n21660), .ZN(n34706));
    INVX1 U21835 (.I(n21329), .ZN(N34707));
    INVX1 U21836 (.I(n18352), .ZN(N34708));
    INVX1 U21837 (.I(N6404), .ZN(n34709));
    INVX1 U21838 (.I(n27496), .ZN(n34710));
    NANDX1 U21839 (.A1(n15119), .A2(n14714), .ZN(N34711));
    NANDX1 U21840 (.A1(n26407), .A2(n17213), .ZN(N34712));
    NANDX1 U21841 (.A1(n22750), .A2(N10480), .ZN(N34713));
    NOR2X1 U21842 (.A1(n24538), .A2(n16488), .ZN(n34714));
    NOR2X1 U21843 (.A1(N8205), .A2(n19258), .ZN(n34715));
    NANDX1 U21844 (.A1(n18997), .A2(n27474), .ZN(n34716));
    INVX1 U21845 (.I(N12530), .ZN(n34717));
    NANDX1 U21846 (.A1(n15430), .A2(n22750), .ZN(n34718));
    INVX1 U21847 (.I(N6621), .ZN(N34719));
    NOR2X1 U21848 (.A1(n28554), .A2(n17008), .ZN(N34720));
    INVX1 U21849 (.I(n21858), .ZN(n34721));
    NOR2X1 U21850 (.A1(n19243), .A2(N6839), .ZN(N34722));
    NANDX1 U21851 (.A1(N4109), .A2(N3108), .ZN(n34723));
    INVX1 U21852 (.I(n16707), .ZN(N34724));
    INVX1 U21853 (.I(N3756), .ZN(N34725));
    INVX1 U21854 (.I(N8818), .ZN(N34726));
    NOR2X1 U21855 (.A1(n14247), .A2(n17022), .ZN(N34727));
    INVX1 U21856 (.I(N5482), .ZN(N34728));
    INVX1 U21857 (.I(n13958), .ZN(N34729));
    NOR2X1 U21858 (.A1(N6972), .A2(n21263), .ZN(N34730));
    NOR2X1 U21859 (.A1(n18282), .A2(N1328), .ZN(N34731));
    NOR2X1 U21860 (.A1(N1299), .A2(n29881), .ZN(N34732));
    NANDX1 U21861 (.A1(n28115), .A2(N10162), .ZN(n34733));
    NOR2X1 U21862 (.A1(n17220), .A2(n17000), .ZN(n34734));
    INVX1 U21863 (.I(n21328), .ZN(N34735));
    NOR2X1 U21864 (.A1(n14048), .A2(n26596), .ZN(n34736));
    NOR2X1 U21865 (.A1(N6364), .A2(n19722), .ZN(n34737));
    INVX1 U21866 (.I(n15167), .ZN(N34738));
    NANDX1 U21867 (.A1(n18787), .A2(N1651), .ZN(n34739));
    INVX1 U21868 (.I(n13229), .ZN(n34740));
    NOR2X1 U21869 (.A1(n23476), .A2(N8761), .ZN(N34741));
    NANDX1 U21870 (.A1(n22932), .A2(n27043), .ZN(N34742));
    NOR2X1 U21871 (.A1(n29008), .A2(n16902), .ZN(N34743));
    INVX1 U21872 (.I(N10516), .ZN(N34744));
    NANDX1 U21873 (.A1(n25225), .A2(n25087), .ZN(N34745));
    NOR2X1 U21874 (.A1(N12087), .A2(n15721), .ZN(N34746));
    NANDX1 U21875 (.A1(n20755), .A2(n18329), .ZN(n34747));
    INVX1 U21876 (.I(n13702), .ZN(N34748));
    NOR2X1 U21877 (.A1(n16589), .A2(n15467), .ZN(N34749));
    NANDX1 U21878 (.A1(N8981), .A2(n22815), .ZN(N34750));
    INVX1 U21879 (.I(N6853), .ZN(N34751));
    NOR2X1 U21880 (.A1(n15539), .A2(n18890), .ZN(N34752));
    NANDX1 U21881 (.A1(N10833), .A2(N245), .ZN(N34753));
    NANDX1 U21882 (.A1(N7454), .A2(n29253), .ZN(N34754));
    NOR2X1 U21883 (.A1(N11077), .A2(n28329), .ZN(n34755));
    INVX1 U21884 (.I(N6164), .ZN(N34756));
    NOR2X1 U21885 (.A1(N6814), .A2(n18251), .ZN(n34757));
    NANDX1 U21886 (.A1(N7223), .A2(n27566), .ZN(N34758));
    INVX1 U21887 (.I(n22789), .ZN(n34759));
    NOR2X1 U21888 (.A1(n17564), .A2(N9240), .ZN(n34760));
    NANDX1 U21889 (.A1(n15846), .A2(n18220), .ZN(n34761));
    NANDX1 U21890 (.A1(n15777), .A2(n25073), .ZN(n34762));
    NANDX1 U21891 (.A1(n19877), .A2(N2386), .ZN(N34763));
    NOR2X1 U21892 (.A1(n19270), .A2(N2630), .ZN(N34764));
    INVX1 U21893 (.I(n15284), .ZN(n34765));
    NOR2X1 U21894 (.A1(N2894), .A2(n26360), .ZN(N34766));
    INVX1 U21895 (.I(n19186), .ZN(N34767));
    NOR2X1 U21896 (.A1(N335), .A2(n25999), .ZN(n34768));
    INVX1 U21897 (.I(N5016), .ZN(N34769));
    NANDX1 U21898 (.A1(N6626), .A2(N9327), .ZN(n34770));
    NANDX1 U21899 (.A1(N6316), .A2(n26890), .ZN(N34771));
    INVX1 U21900 (.I(n21473), .ZN(N34772));
    NANDX1 U21901 (.A1(N317), .A2(n17868), .ZN(N34773));
    NOR2X1 U21902 (.A1(n13950), .A2(n27428), .ZN(N34774));
    NOR2X1 U21903 (.A1(n16335), .A2(N10077), .ZN(N34775));
    NOR2X1 U21904 (.A1(n18964), .A2(n18816), .ZN(n34776));
    NANDX1 U21905 (.A1(n27968), .A2(n21709), .ZN(N34777));
    NOR2X1 U21906 (.A1(n16464), .A2(n29456), .ZN(N34778));
    NANDX1 U21907 (.A1(N5360), .A2(n25317), .ZN(n34779));
    NOR2X1 U21908 (.A1(N10375), .A2(N5523), .ZN(N34780));
    INVX1 U21909 (.I(N8262), .ZN(N34781));
    NOR2X1 U21910 (.A1(n20397), .A2(N5014), .ZN(n34782));
    NANDX1 U21911 (.A1(N293), .A2(N6173), .ZN(n34783));
    NOR2X1 U21912 (.A1(N6722), .A2(n23108), .ZN(n34784));
    NANDX1 U21913 (.A1(N4012), .A2(n18343), .ZN(n34785));
    INVX1 U21914 (.I(n14088), .ZN(n34786));
    NANDX1 U21915 (.A1(n17298), .A2(n21464), .ZN(N34787));
    INVX1 U21916 (.I(n15128), .ZN(N34788));
    INVX1 U21917 (.I(N9671), .ZN(N34789));
    NOR2X1 U21918 (.A1(N915), .A2(N7930), .ZN(n34790));
    NANDX1 U21919 (.A1(n14792), .A2(n15385), .ZN(n34791));
    INVX1 U21920 (.I(n20315), .ZN(n34792));
    NANDX1 U21921 (.A1(N2571), .A2(n28831), .ZN(n34793));
    NOR2X1 U21922 (.A1(n26282), .A2(n19444), .ZN(N34794));
    INVX1 U21923 (.I(N2317), .ZN(N34795));
    NANDX1 U21924 (.A1(n15299), .A2(n25424), .ZN(N34796));
    INVX1 U21925 (.I(n19310), .ZN(N34797));
    INVX1 U21926 (.I(n13585), .ZN(n34798));
    NANDX1 U21927 (.A1(n16338), .A2(n19444), .ZN(N34799));
    NOR2X1 U21928 (.A1(n30136), .A2(N4434), .ZN(N34800));
    NOR2X1 U21929 (.A1(n28368), .A2(n24586), .ZN(n34801));
    INVX1 U21930 (.I(N6160), .ZN(n34802));
    INVX1 U21931 (.I(n19148), .ZN(n34803));
    NANDX1 U21932 (.A1(n21528), .A2(n28023), .ZN(N34804));
    NOR2X1 U21933 (.A1(N12659), .A2(n26716), .ZN(n34805));
    NOR2X1 U21934 (.A1(N8804), .A2(n16023), .ZN(N34806));
    INVX1 U21935 (.I(N11120), .ZN(N34807));
    NOR2X1 U21936 (.A1(N11457), .A2(n25105), .ZN(N34808));
    INVX1 U21937 (.I(n19328), .ZN(N34809));
    INVX1 U21938 (.I(n20913), .ZN(N34810));
    NOR2X1 U21939 (.A1(N2056), .A2(N10219), .ZN(N34811));
    NANDX1 U21940 (.A1(n20752), .A2(N3214), .ZN(n34812));
    NANDX1 U21941 (.A1(n18982), .A2(n16360), .ZN(n34813));
    NOR2X1 U21942 (.A1(n25141), .A2(n24881), .ZN(N34814));
    NANDX1 U21943 (.A1(n16548), .A2(N4832), .ZN(N34815));
    NOR2X1 U21944 (.A1(n25980), .A2(n17491), .ZN(n34816));
    INVX1 U21945 (.I(n25000), .ZN(n34817));
    INVX1 U21946 (.I(N4668), .ZN(N34818));
    INVX1 U21947 (.I(n25974), .ZN(n34819));
    NANDX1 U21948 (.A1(n21175), .A2(N9502), .ZN(n34820));
    NANDX1 U21949 (.A1(N10365), .A2(n25357), .ZN(N34821));
    NANDX1 U21950 (.A1(n28772), .A2(n27412), .ZN(N34822));
    INVX1 U21951 (.I(N190), .ZN(N34823));
    INVX1 U21952 (.I(N8280), .ZN(n34824));
    NOR2X1 U21953 (.A1(n25569), .A2(n24640), .ZN(n34825));
    NOR2X1 U21954 (.A1(n20572), .A2(N7944), .ZN(N34826));
    NOR2X1 U21955 (.A1(n25680), .A2(N1336), .ZN(N34827));
    NANDX1 U21956 (.A1(N10084), .A2(n18826), .ZN(n34828));
    NANDX1 U21957 (.A1(n23644), .A2(N3543), .ZN(N34829));
    INVX1 U21958 (.I(N3225), .ZN(N34830));
    INVX1 U21959 (.I(n20979), .ZN(N34831));
    NANDX1 U21960 (.A1(n16140), .A2(N6353), .ZN(N34832));
    NANDX1 U21961 (.A1(N11359), .A2(N12640), .ZN(N34833));
    NOR2X1 U21962 (.A1(n27331), .A2(N6268), .ZN(n34834));
    INVX1 U21963 (.I(n15220), .ZN(n34835));
    INVX1 U21964 (.I(n23153), .ZN(N34836));
    NANDX1 U21965 (.A1(n27747), .A2(N3373), .ZN(N34837));
    INVX1 U21966 (.I(N5553), .ZN(n34838));
    NOR2X1 U21967 (.A1(N3887), .A2(N6889), .ZN(N34839));
    INVX1 U21968 (.I(N2531), .ZN(N34840));
    NANDX1 U21969 (.A1(n16823), .A2(n26174), .ZN(N34841));
    NANDX1 U21970 (.A1(n18178), .A2(n29398), .ZN(N34842));
    NOR2X1 U21971 (.A1(N9019), .A2(N12220), .ZN(n34843));
    NOR2X1 U21972 (.A1(N3933), .A2(N5407), .ZN(N34844));
    NOR2X1 U21973 (.A1(N5133), .A2(n15927), .ZN(N34845));
    INVX1 U21974 (.I(N11400), .ZN(n34846));
    NOR2X1 U21975 (.A1(N11351), .A2(n25947), .ZN(N34847));
    NANDX1 U21976 (.A1(N10562), .A2(N12117), .ZN(N34848));
    NANDX1 U21977 (.A1(n18906), .A2(n17670), .ZN(n34849));
    NANDX1 U21978 (.A1(N11353), .A2(n13119), .ZN(N34850));
    NOR2X1 U21979 (.A1(n13883), .A2(n15954), .ZN(N34851));
    INVX1 U21980 (.I(n28617), .ZN(n34852));
    NOR2X1 U21981 (.A1(N10173), .A2(n16438), .ZN(N34853));
    NOR2X1 U21982 (.A1(N7752), .A2(n17218), .ZN(N34854));
    INVX1 U21983 (.I(N11684), .ZN(N34855));
    NOR2X1 U21984 (.A1(n26046), .A2(N5378), .ZN(N34856));
    NOR2X1 U21985 (.A1(N3479), .A2(n16777), .ZN(N34857));
    NOR2X1 U21986 (.A1(n14830), .A2(N1147), .ZN(n34858));
    INVX1 U21987 (.I(n13952), .ZN(n34859));
    INVX1 U21988 (.I(n20525), .ZN(n34860));
    NOR2X1 U21989 (.A1(n19494), .A2(N9881), .ZN(N34861));
    NANDX1 U21990 (.A1(N2475), .A2(n15191), .ZN(n34862));
    INVX1 U21991 (.I(n18428), .ZN(N34863));
    NANDX1 U21992 (.A1(n22253), .A2(N10623), .ZN(n34864));
    NANDX1 U21993 (.A1(N8553), .A2(n15833), .ZN(N34865));
    NOR2X1 U21994 (.A1(n14332), .A2(N1364), .ZN(n34866));
    INVX1 U21995 (.I(N6819), .ZN(N34867));
    NANDX1 U21996 (.A1(n19291), .A2(n22491), .ZN(N34868));
    NOR2X1 U21997 (.A1(n24629), .A2(N4523), .ZN(N34869));
    NOR2X1 U21998 (.A1(n25775), .A2(n24904), .ZN(N34870));
    NOR2X1 U21999 (.A1(N8901), .A2(N3852), .ZN(N34871));
    NOR2X1 U22000 (.A1(n16955), .A2(N2294), .ZN(n34872));
    NANDX1 U22001 (.A1(N7990), .A2(n17484), .ZN(n34873));
    NOR2X1 U22002 (.A1(n26418), .A2(n13229), .ZN(N34874));
    NANDX1 U22003 (.A1(n25601), .A2(n19147), .ZN(n34875));
    INVX1 U22004 (.I(n29994), .ZN(n34876));
    NOR2X1 U22005 (.A1(n16461), .A2(N1221), .ZN(N34877));
    INVX1 U22006 (.I(N11840), .ZN(N34878));
    NOR2X1 U22007 (.A1(N1566), .A2(N4193), .ZN(N34879));
    NANDX1 U22008 (.A1(n26194), .A2(N8715), .ZN(n34880));
    NANDX1 U22009 (.A1(N10392), .A2(n22179), .ZN(N34881));
    NANDX1 U22010 (.A1(N7854), .A2(n26031), .ZN(N34882));
    INVX1 U22011 (.I(n24808), .ZN(N34883));
    NANDX1 U22012 (.A1(n23051), .A2(N2661), .ZN(n34884));
    NOR2X1 U22013 (.A1(N5814), .A2(n17639), .ZN(N34885));
    INVX1 U22014 (.I(N10830), .ZN(N34886));
    NOR2X1 U22015 (.A1(n25166), .A2(n12959), .ZN(n34887));
    NOR2X1 U22016 (.A1(N4966), .A2(n17980), .ZN(n34888));
    NOR2X1 U22017 (.A1(n17378), .A2(n29819), .ZN(N34889));
    NOR2X1 U22018 (.A1(n18943), .A2(N3874), .ZN(n34890));
    NANDX1 U22019 (.A1(n14999), .A2(N1149), .ZN(N34891));
    INVX1 U22020 (.I(n13951), .ZN(n34892));
    NOR2X1 U22021 (.A1(n20046), .A2(n21804), .ZN(N34893));
    INVX1 U22022 (.I(N12394), .ZN(n34894));
    INVX1 U22023 (.I(n24666), .ZN(N34895));
    NANDX1 U22024 (.A1(N7696), .A2(n17457), .ZN(N34896));
    NANDX1 U22025 (.A1(n25334), .A2(n23476), .ZN(N34897));
    NANDX1 U22026 (.A1(n15557), .A2(N7066), .ZN(N34898));
    NOR2X1 U22027 (.A1(n17075), .A2(N12031), .ZN(N34899));
    INVX1 U22028 (.I(N8375), .ZN(N34900));
    NOR2X1 U22029 (.A1(N6812), .A2(n16864), .ZN(N34901));
    NOR2X1 U22030 (.A1(N10685), .A2(N1716), .ZN(n34902));
    NANDX1 U22031 (.A1(N11833), .A2(n15907), .ZN(N34903));
    NOR2X1 U22032 (.A1(n23721), .A2(n24513), .ZN(N34904));
    INVX1 U22033 (.I(n20063), .ZN(n34905));
    NANDX1 U22034 (.A1(n20985), .A2(N3152), .ZN(N34906));
    NANDX1 U22035 (.A1(n28680), .A2(n20608), .ZN(N34907));
    NOR2X1 U22036 (.A1(N12437), .A2(n13947), .ZN(N34908));
    NANDX1 U22037 (.A1(n27993), .A2(N9573), .ZN(N34909));
    INVX1 U22038 (.I(N3492), .ZN(N34910));
    INVX1 U22039 (.I(N2929), .ZN(N34911));
    INVX1 U22040 (.I(n28133), .ZN(N34912));
    NOR2X1 U22041 (.A1(n28729), .A2(N4769), .ZN(N34913));
    INVX1 U22042 (.I(n19005), .ZN(N34914));
    NOR2X1 U22043 (.A1(N9378), .A2(N4775), .ZN(N34915));
    NOR2X1 U22044 (.A1(n21660), .A2(n29287), .ZN(n34916));
    INVX1 U22045 (.I(N146), .ZN(N34917));
    INVX1 U22046 (.I(n23304), .ZN(N34918));
    NANDX1 U22047 (.A1(n13814), .A2(N10407), .ZN(N34919));
    INVX1 U22048 (.I(n21390), .ZN(N34920));
    INVX1 U22049 (.I(n26412), .ZN(N34921));
    NANDX1 U22050 (.A1(N9260), .A2(N5847), .ZN(N34922));
    NOR2X1 U22051 (.A1(N12751), .A2(n16011), .ZN(N34923));
    INVX1 U22052 (.I(n13177), .ZN(n34924));
    NOR2X1 U22053 (.A1(n20883), .A2(N11768), .ZN(N34925));
    INVX1 U22054 (.I(n18428), .ZN(N34926));
    NANDX1 U22055 (.A1(N10997), .A2(n16366), .ZN(n34927));
    NOR2X1 U22056 (.A1(N8805), .A2(n26586), .ZN(N34928));
    INVX1 U22057 (.I(N11124), .ZN(N34929));
    INVX1 U22058 (.I(N6297), .ZN(n34930));
    INVX1 U22059 (.I(n30029), .ZN(n34931));
    NOR2X1 U22060 (.A1(N3257), .A2(N12357), .ZN(N34932));
    NOR2X1 U22061 (.A1(n14661), .A2(N8632), .ZN(N34933));
    NANDX1 U22062 (.A1(N12482), .A2(N3039), .ZN(N34934));
    INVX1 U22063 (.I(n13793), .ZN(n34935));
    NOR2X1 U22064 (.A1(n17180), .A2(n26970), .ZN(n34936));
    NOR2X1 U22065 (.A1(n26623), .A2(n27298), .ZN(N34937));
    INVX1 U22066 (.I(n14913), .ZN(N34938));
    NANDX1 U22067 (.A1(n28507), .A2(n19840), .ZN(N34939));
    INVX1 U22068 (.I(N7175), .ZN(N34940));
    INVX1 U22069 (.I(N10843), .ZN(n34941));
    NANDX1 U22070 (.A1(N1443), .A2(N5700), .ZN(n34942));
    NANDX1 U22071 (.A1(N1334), .A2(n14371), .ZN(n34943));
    NANDX1 U22072 (.A1(N2252), .A2(n14293), .ZN(N34944));
    NANDX1 U22073 (.A1(N10883), .A2(N7935), .ZN(N34945));
    NANDX1 U22074 (.A1(N2482), .A2(n13971), .ZN(N34946));
    INVX1 U22075 (.I(N10092), .ZN(n34947));
    NOR2X1 U22076 (.A1(n17853), .A2(n20267), .ZN(N34948));
    INVX1 U22077 (.I(n15014), .ZN(n34949));
    INVX1 U22078 (.I(n19671), .ZN(n34950));
    NOR2X1 U22079 (.A1(n24708), .A2(N9373), .ZN(N34951));
    NANDX1 U22080 (.A1(n20443), .A2(n14221), .ZN(n34952));
    INVX1 U22081 (.I(n15862), .ZN(N34953));
    INVX1 U22082 (.I(N5497), .ZN(N34954));
    NOR2X1 U22083 (.A1(N5558), .A2(n19867), .ZN(n34955));
    INVX1 U22084 (.I(N7809), .ZN(N34956));
    NOR2X1 U22085 (.A1(N1842), .A2(N7252), .ZN(N34957));
    NANDX1 U22086 (.A1(N9070), .A2(N9734), .ZN(N34958));
    NANDX1 U22087 (.A1(n18652), .A2(N8386), .ZN(N34959));
    INVX1 U22088 (.I(N6367), .ZN(N34960));
    NOR2X1 U22089 (.A1(N8820), .A2(N9941), .ZN(N34961));
    INVX1 U22090 (.I(n28490), .ZN(N34962));
    NOR2X1 U22091 (.A1(n26682), .A2(n26423), .ZN(N34963));
    INVX1 U22092 (.I(N5548), .ZN(n34964));
    INVX1 U22093 (.I(N63), .ZN(N34965));
    INVX1 U22094 (.I(n14730), .ZN(n34966));
    NOR2X1 U22095 (.A1(n25539), .A2(n20288), .ZN(N34967));
    NOR2X1 U22096 (.A1(N2496), .A2(n28096), .ZN(N34968));
    NANDX1 U22097 (.A1(n23036), .A2(n23909), .ZN(n34969));
    INVX1 U22098 (.I(n20666), .ZN(N34970));
    NOR2X1 U22099 (.A1(n28833), .A2(N9180), .ZN(n34971));
    NOR2X1 U22100 (.A1(N10017), .A2(N4108), .ZN(n34972));
    NANDX1 U22101 (.A1(n18836), .A2(n14048), .ZN(n34973));
    NOR2X1 U22102 (.A1(N5749), .A2(n13919), .ZN(n34974));
    NOR2X1 U22103 (.A1(n20732), .A2(N2745), .ZN(n34975));
    NANDX1 U22104 (.A1(N1100), .A2(n21505), .ZN(n34976));
    NOR2X1 U22105 (.A1(N4391), .A2(n15625), .ZN(N34977));
    NOR2X1 U22106 (.A1(n24678), .A2(n29611), .ZN(N34978));
    NANDX1 U22107 (.A1(N11197), .A2(n24741), .ZN(N34979));
    NOR2X1 U22108 (.A1(N4968), .A2(n20388), .ZN(n34980));
    NOR2X1 U22109 (.A1(n27170), .A2(N7644), .ZN(n34981));
    NANDX1 U22110 (.A1(n27620), .A2(n17660), .ZN(N34982));
    NANDX1 U22111 (.A1(N3707), .A2(n25056), .ZN(N34983));
    NANDX1 U22112 (.A1(N11904), .A2(n19365), .ZN(N34984));
    NOR2X1 U22113 (.A1(n16646), .A2(N9959), .ZN(N34985));
    INVX1 U22114 (.I(n15495), .ZN(N34986));
    NOR2X1 U22115 (.A1(n28586), .A2(N5616), .ZN(N34987));
    NOR2X1 U22116 (.A1(n14073), .A2(N9835), .ZN(N34988));
    NANDX1 U22117 (.A1(N2107), .A2(n16550), .ZN(n34989));
    NANDX1 U22118 (.A1(n15408), .A2(N4724), .ZN(N34990));
    NOR2X1 U22119 (.A1(n24356), .A2(n13564), .ZN(n34991));
    INVX1 U22120 (.I(N1862), .ZN(N34992));
    NANDX1 U22121 (.A1(N5049), .A2(n19522), .ZN(N34993));
    NOR2X1 U22122 (.A1(N8755), .A2(n14440), .ZN(N34994));
    NANDX1 U22123 (.A1(n20658), .A2(N3668), .ZN(N34995));
    NANDX1 U22124 (.A1(n25864), .A2(n13626), .ZN(N34996));
    NOR2X1 U22125 (.A1(N11222), .A2(N1806), .ZN(n34997));
    NANDX1 U22126 (.A1(N5398), .A2(N5815), .ZN(n34998));
    INVX1 U22127 (.I(n15232), .ZN(N34999));
    INVX1 U22128 (.I(N9895), .ZN(N35000));
    NANDX1 U22129 (.A1(n21369), .A2(n13863), .ZN(N35001));
    NANDX1 U22130 (.A1(n24643), .A2(N8081), .ZN(N35002));
    NANDX1 U22131 (.A1(N2071), .A2(N9942), .ZN(n35003));
    INVX1 U22132 (.I(N7119), .ZN(n35004));
    INVX1 U22133 (.I(n25148), .ZN(N35005));
    NANDX1 U22134 (.A1(N2327), .A2(N9000), .ZN(N35006));
    NOR2X1 U22135 (.A1(n24692), .A2(n27324), .ZN(N35007));
    NANDX1 U22136 (.A1(N8180), .A2(N3894), .ZN(n35008));
    INVX1 U22137 (.I(N9986), .ZN(N35009));
    NOR2X1 U22138 (.A1(n25997), .A2(N4361), .ZN(n35010));
    NOR2X1 U22139 (.A1(N11092), .A2(n27423), .ZN(n35011));
    NANDX1 U22140 (.A1(N1297), .A2(n18654), .ZN(n35012));
    INVX1 U22141 (.I(n14923), .ZN(N35013));
    NANDX1 U22142 (.A1(N7097), .A2(N11976), .ZN(n35014));
    NOR2X1 U22143 (.A1(N5600), .A2(n17732), .ZN(N35015));
    NANDX1 U22144 (.A1(n23623), .A2(N12743), .ZN(n35016));
    NOR2X1 U22145 (.A1(n25949), .A2(N10303), .ZN(N35017));
    NOR2X1 U22146 (.A1(n20503), .A2(N7489), .ZN(N35018));
    NOR2X1 U22147 (.A1(n17244), .A2(n30081), .ZN(N35019));
    NOR2X1 U22148 (.A1(n15790), .A2(N8992), .ZN(N35020));
    INVX1 U22149 (.I(n20150), .ZN(N35021));
    INVX1 U22150 (.I(N5649), .ZN(N35022));
    INVX1 U22151 (.I(n29681), .ZN(n35023));
    NANDX1 U22152 (.A1(n24649), .A2(n28698), .ZN(N35024));
    NANDX1 U22153 (.A1(n26368), .A2(n24355), .ZN(N35025));
    NANDX1 U22154 (.A1(N21), .A2(n18515), .ZN(N35026));
    NANDX1 U22155 (.A1(N10929), .A2(N12001), .ZN(N35027));
    NOR2X1 U22156 (.A1(n26270), .A2(n26510), .ZN(N35028));
    NOR2X1 U22157 (.A1(n25127), .A2(N5437), .ZN(N35029));
    NANDX1 U22158 (.A1(n14664), .A2(N11241), .ZN(N35030));
    NOR2X1 U22159 (.A1(n24800), .A2(n27030), .ZN(n35031));
    NANDX1 U22160 (.A1(n19357), .A2(N5603), .ZN(N35032));
    NANDX1 U22161 (.A1(n25005), .A2(N11599), .ZN(N35033));
    INVX1 U22162 (.I(n20510), .ZN(N35034));
    NANDX1 U22163 (.A1(n27640), .A2(N801), .ZN(N35035));
    INVX1 U22164 (.I(N10419), .ZN(N35036));
    NOR2X1 U22165 (.A1(n21059), .A2(n28933), .ZN(n35037));
    INVX1 U22166 (.I(n20548), .ZN(n35038));
    NANDX1 U22167 (.A1(N2924), .A2(n16680), .ZN(N35039));
    NOR2X1 U22168 (.A1(n13087), .A2(N11669), .ZN(n35040));
    NANDX1 U22169 (.A1(N602), .A2(n14893), .ZN(n35041));
    INVX1 U22170 (.I(N6757), .ZN(N35042));
    NOR2X1 U22171 (.A1(n27996), .A2(n21904), .ZN(N35043));
    NOR2X1 U22172 (.A1(n22159), .A2(n21303), .ZN(n35044));
    INVX1 U22173 (.I(n22318), .ZN(N35045));
    NANDX1 U22174 (.A1(n21411), .A2(n16989), .ZN(N35046));
    NOR2X1 U22175 (.A1(n22211), .A2(N7890), .ZN(n35047));
    NANDX1 U22176 (.A1(n15277), .A2(n17509), .ZN(N35048));
    NOR2X1 U22177 (.A1(N6900), .A2(N7919), .ZN(N35049));
    NANDX1 U22178 (.A1(N9824), .A2(n13159), .ZN(N35050));
    INVX1 U22179 (.I(n22910), .ZN(n35051));
    NOR2X1 U22180 (.A1(N334), .A2(N12072), .ZN(N35052));
    NOR2X1 U22181 (.A1(N1300), .A2(N7390), .ZN(N35053));
    NOR2X1 U22182 (.A1(n29295), .A2(n29293), .ZN(N35054));
    NOR2X1 U22183 (.A1(N9878), .A2(n20459), .ZN(N35055));
    INVX1 U22184 (.I(N2058), .ZN(N35056));
    NANDX1 U22185 (.A1(n24605), .A2(N7607), .ZN(N35057));
    INVX1 U22186 (.I(N5240), .ZN(N35058));
    INVX1 U22187 (.I(N3465), .ZN(N35059));
    NOR2X1 U22188 (.A1(N10126), .A2(N7548), .ZN(N35060));
    NOR2X1 U22189 (.A1(N6605), .A2(n22426), .ZN(n35061));
    NANDX1 U22190 (.A1(n19764), .A2(N2897), .ZN(N35062));
    NANDX1 U22191 (.A1(N3015), .A2(n21928), .ZN(N35063));
    INVX1 U22192 (.I(n19856), .ZN(N35064));
    INVX1 U22193 (.I(N3715), .ZN(N35065));
    NOR2X1 U22194 (.A1(N10946), .A2(N2871), .ZN(N35066));
    NOR2X1 U22195 (.A1(N9384), .A2(N11890), .ZN(N35067));
    NOR2X1 U22196 (.A1(N11442), .A2(N11017), .ZN(n35068));
    NANDX1 U22197 (.A1(N7609), .A2(n16452), .ZN(N35069));
    INVX1 U22198 (.I(N11666), .ZN(N35070));
    NOR2X1 U22199 (.A1(n18946), .A2(N10352), .ZN(N35071));
    NOR2X1 U22200 (.A1(n23483), .A2(n16957), .ZN(n35072));
    NOR2X1 U22201 (.A1(N7705), .A2(N6583), .ZN(N35073));
    NOR2X1 U22202 (.A1(n22096), .A2(n28295), .ZN(N35074));
    NANDX1 U22203 (.A1(n18422), .A2(n18013), .ZN(n35075));
    NOR2X1 U22204 (.A1(n22136), .A2(n22689), .ZN(n35076));
    NANDX1 U22205 (.A1(n13567), .A2(N10960), .ZN(N35077));
    INVX1 U22206 (.I(n14017), .ZN(N35078));
    INVX1 U22207 (.I(N12240), .ZN(n35079));
    NANDX1 U22208 (.A1(n25754), .A2(N8410), .ZN(n35080));
    INVX1 U22209 (.I(N5486), .ZN(n35081));
    INVX1 U22210 (.I(n27083), .ZN(N35082));
    INVX1 U22211 (.I(N289), .ZN(N35083));
    NANDX1 U22212 (.A1(N6338), .A2(n17245), .ZN(n35084));
    INVX1 U22213 (.I(N2603), .ZN(N35085));
    NANDX1 U22214 (.A1(N5432), .A2(n13260), .ZN(N35086));
    NANDX1 U22215 (.A1(n15689), .A2(N1544), .ZN(N35087));
    INVX1 U22216 (.I(N7598), .ZN(N35088));
    NOR2X1 U22217 (.A1(n28368), .A2(n29150), .ZN(N35089));
    NANDX1 U22218 (.A1(N9191), .A2(N11250), .ZN(n35090));
    NANDX1 U22219 (.A1(N176), .A2(N12051), .ZN(N35091));
    INVX1 U22220 (.I(n25929), .ZN(N35092));
    NANDX1 U22221 (.A1(N11749), .A2(n19976), .ZN(N35093));
    NOR2X1 U22222 (.A1(n27392), .A2(n21529), .ZN(n35094));
    NOR2X1 U22223 (.A1(n28922), .A2(n27866), .ZN(N35095));
    NOR2X1 U22224 (.A1(n15886), .A2(n19029), .ZN(N35096));
    INVX1 U22225 (.I(n21317), .ZN(N35097));
    NOR2X1 U22226 (.A1(N5106), .A2(n25567), .ZN(N35098));
    NANDX1 U22227 (.A1(N10785), .A2(N3027), .ZN(N35099));
    NOR2X1 U22228 (.A1(N9015), .A2(n20737), .ZN(N35100));
    NANDX1 U22229 (.A1(N6766), .A2(N1849), .ZN(N35101));
    NOR2X1 U22230 (.A1(n25640), .A2(N2460), .ZN(n35102));
    NOR2X1 U22231 (.A1(n21431), .A2(n22919), .ZN(N35103));
    NANDX1 U22232 (.A1(n29967), .A2(N10437), .ZN(N35104));
    NANDX1 U22233 (.A1(n21358), .A2(n28381), .ZN(n35105));
    NANDX1 U22234 (.A1(N7647), .A2(n21993), .ZN(n35106));
    NANDX1 U22235 (.A1(n15237), .A2(n16553), .ZN(N35107));
    INVX1 U22236 (.I(n17387), .ZN(N35108));
    NANDX1 U22237 (.A1(N9092), .A2(N9642), .ZN(N35109));
    NOR2X1 U22238 (.A1(N679), .A2(n14136), .ZN(N35110));
    NOR2X1 U22239 (.A1(n21415), .A2(n14299), .ZN(N35111));
    INVX1 U22240 (.I(N11825), .ZN(n35112));
    NOR2X1 U22241 (.A1(n20846), .A2(n14284), .ZN(N35113));
    INVX1 U22242 (.I(N701), .ZN(n35114));
    NOR2X1 U22243 (.A1(N7559), .A2(N530), .ZN(N35115));
    NANDX1 U22244 (.A1(N8113), .A2(N10449), .ZN(n35116));
    INVX1 U22245 (.I(n26150), .ZN(N35117));
    INVX1 U22246 (.I(n14859), .ZN(N35118));
    INVX1 U22247 (.I(n21892), .ZN(N35119));
    NOR2X1 U22248 (.A1(n13460), .A2(N9142), .ZN(N35120));
    NANDX1 U22249 (.A1(N11113), .A2(N7344), .ZN(n35121));
    NANDX1 U22250 (.A1(N11791), .A2(n21479), .ZN(n35122));
    NANDX1 U22251 (.A1(N3069), .A2(n24338), .ZN(N35123));
    NANDX1 U22252 (.A1(n14893), .A2(N6908), .ZN(n35124));
    NANDX1 U22253 (.A1(n29176), .A2(N11167), .ZN(N35125));
    INVX1 U22254 (.I(n13363), .ZN(N35126));
    NOR2X1 U22255 (.A1(n26779), .A2(n19426), .ZN(n35127));
    NOR2X1 U22256 (.A1(N7090), .A2(N12292), .ZN(N35128));
    NANDX1 U22257 (.A1(N2307), .A2(n27151), .ZN(N35129));
    NOR2X1 U22258 (.A1(n24198), .A2(n16986), .ZN(n35130));
    NANDX1 U22259 (.A1(N3202), .A2(n28478), .ZN(N35131));
    NANDX1 U22260 (.A1(N10545), .A2(N699), .ZN(N35132));
    NOR2X1 U22261 (.A1(n20584), .A2(N10196), .ZN(N35133));
    INVX1 U22262 (.I(n14784), .ZN(N35134));
    NANDX1 U22263 (.A1(N1076), .A2(N10253), .ZN(N35135));
    INVX1 U22264 (.I(n18813), .ZN(N35136));
    INVX1 U22265 (.I(n17863), .ZN(n35137));
    NOR2X1 U22266 (.A1(n28705), .A2(n14504), .ZN(n35138));
    NOR2X1 U22267 (.A1(N2528), .A2(N10155), .ZN(N35139));
    NOR2X1 U22268 (.A1(N2499), .A2(N12461), .ZN(N35140));
    NANDX1 U22269 (.A1(n20966), .A2(N6521), .ZN(n35141));
    NOR2X1 U22270 (.A1(n22755), .A2(n28421), .ZN(n35142));
    NANDX1 U22271 (.A1(n24217), .A2(n27526), .ZN(N35143));
    INVX1 U22272 (.I(N7332), .ZN(N35144));
    NOR2X1 U22273 (.A1(n29929), .A2(n23653), .ZN(N35145));
    NANDX1 U22274 (.A1(n26130), .A2(n13289), .ZN(N35146));
    NANDX1 U22275 (.A1(N6304), .A2(n20662), .ZN(N35147));
    INVX1 U22276 (.I(n24166), .ZN(N35148));
    NANDX1 U22277 (.A1(n28677), .A2(n27231), .ZN(N35149));
    INVX1 U22278 (.I(n19765), .ZN(N35150));
    INVX1 U22279 (.I(n20721), .ZN(N35151));
    NANDX1 U22280 (.A1(N8269), .A2(n17171), .ZN(N35152));
    NOR2X1 U22281 (.A1(N3350), .A2(N469), .ZN(N35153));
    NOR2X1 U22282 (.A1(N1633), .A2(N806), .ZN(N35154));
    INVX1 U22283 (.I(n17720), .ZN(N35155));
    NANDX1 U22284 (.A1(n25817), .A2(n24253), .ZN(N35156));
    NANDX1 U22285 (.A1(N7893), .A2(n15432), .ZN(n35157));
    NANDX1 U22286 (.A1(n21182), .A2(N5425), .ZN(n35158));
    INVX1 U22287 (.I(N267), .ZN(N35159));
    NANDX1 U22288 (.A1(n23914), .A2(N11527), .ZN(N35160));
    INVX1 U22289 (.I(n21007), .ZN(N35161));
    NANDX1 U22290 (.A1(N12262), .A2(n16815), .ZN(n35162));
    NANDX1 U22291 (.A1(N4388), .A2(n25083), .ZN(N35163));
    NANDX1 U22292 (.A1(n17479), .A2(n16993), .ZN(n35164));
    NANDX1 U22293 (.A1(N11748), .A2(N7187), .ZN(n35165));
    NOR2X1 U22294 (.A1(n18794), .A2(n24906), .ZN(N35166));
    INVX1 U22295 (.I(n14473), .ZN(N35167));
    NOR2X1 U22296 (.A1(N6813), .A2(N10927), .ZN(N35168));
    INVX1 U22297 (.I(N11696), .ZN(N35169));
    NANDX1 U22298 (.A1(n28437), .A2(N11443), .ZN(n35170));
    INVX1 U22299 (.I(n22394), .ZN(N35171));
    NANDX1 U22300 (.A1(N2325), .A2(n14891), .ZN(N35172));
    NOR2X1 U22301 (.A1(n23696), .A2(n27152), .ZN(N35173));
    NOR2X1 U22302 (.A1(n24211), .A2(N1402), .ZN(N35174));
    NANDX1 U22303 (.A1(N11760), .A2(N7441), .ZN(N35175));
    INVX1 U22304 (.I(n29915), .ZN(N35176));
    NOR2X1 U22305 (.A1(N9148), .A2(n25996), .ZN(N35177));
    INVX1 U22306 (.I(N3916), .ZN(N35178));
    NOR2X1 U22307 (.A1(N10877), .A2(n22936), .ZN(N35179));
    NOR2X1 U22308 (.A1(n21803), .A2(n15811), .ZN(N35180));
    INVX1 U22309 (.I(N12334), .ZN(N35181));
    NOR2X1 U22310 (.A1(N12291), .A2(N3132), .ZN(n35182));
    NANDX1 U22311 (.A1(N6071), .A2(n24154), .ZN(n35183));
    NANDX1 U22312 (.A1(n20856), .A2(n17712), .ZN(n35184));
    NOR2X1 U22313 (.A1(n22319), .A2(N11785), .ZN(N35185));
    INVX1 U22314 (.I(N7287), .ZN(N35186));
    INVX1 U22315 (.I(N4234), .ZN(N35187));
    NANDX1 U22316 (.A1(N11883), .A2(N11982), .ZN(N35188));
    NOR2X1 U22317 (.A1(n26439), .A2(n19825), .ZN(N35189));
    INVX1 U22318 (.I(N8780), .ZN(N35190));
    NANDX1 U22319 (.A1(N3669), .A2(n28070), .ZN(N35191));
    NANDX1 U22320 (.A1(N8041), .A2(n17479), .ZN(N35192));
    NANDX1 U22321 (.A1(N10712), .A2(n18331), .ZN(N35193));
    NANDX1 U22322 (.A1(n24337), .A2(n24401), .ZN(n35194));
    NANDX1 U22323 (.A1(N4018), .A2(n15119), .ZN(n35195));
    NOR2X1 U22324 (.A1(n29547), .A2(n25998), .ZN(N35196));
    NANDX1 U22325 (.A1(n26341), .A2(N3148), .ZN(N35197));
    NOR2X1 U22326 (.A1(N437), .A2(N12395), .ZN(N35198));
    NANDX1 U22327 (.A1(N12419), .A2(n19351), .ZN(N35199));
    NANDX1 U22328 (.A1(n20804), .A2(N84), .ZN(N35200));
    INVX1 U22329 (.I(n28627), .ZN(n35201));
    NANDX1 U22330 (.A1(N8271), .A2(n28116), .ZN(n35202));
    NOR2X1 U22331 (.A1(n14310), .A2(n17060), .ZN(N35203));
    NANDX1 U22332 (.A1(N2503), .A2(N9135), .ZN(N35204));
    INVX1 U22333 (.I(n15464), .ZN(n35205));
    NOR2X1 U22334 (.A1(n27979), .A2(n19144), .ZN(N35206));
    NOR2X1 U22335 (.A1(n15950), .A2(n15004), .ZN(N35207));
    NANDX1 U22336 (.A1(N12153), .A2(n18151), .ZN(N35208));
    NANDX1 U22337 (.A1(N1150), .A2(n19107), .ZN(N35209));
    INVX1 U22338 (.I(n13568), .ZN(N35210));
    NOR2X1 U22339 (.A1(N3364), .A2(n22933), .ZN(N35211));
    NANDX1 U22340 (.A1(n13702), .A2(n21422), .ZN(N35212));
    INVX1 U22341 (.I(N10533), .ZN(n35213));
    NANDX1 U22342 (.A1(N1069), .A2(n24842), .ZN(n35214));
    NANDX1 U22343 (.A1(N694), .A2(n15906), .ZN(N35215));
    INVX1 U22344 (.I(n24656), .ZN(n35216));
    NANDX1 U22345 (.A1(n17940), .A2(N11058), .ZN(N35217));
    NOR2X1 U22346 (.A1(n24226), .A2(n15568), .ZN(N35218));
    INVX1 U22347 (.I(N4523), .ZN(n35219));
    INVX1 U22348 (.I(N514), .ZN(N35220));
    INVX1 U22349 (.I(n28870), .ZN(N35221));
    NOR2X1 U22350 (.A1(N10136), .A2(N861), .ZN(N35222));
    NANDX1 U22351 (.A1(n13500), .A2(n23793), .ZN(n35223));
    NANDX1 U22352 (.A1(n27201), .A2(N3639), .ZN(N35224));
    NOR2X1 U22353 (.A1(n26294), .A2(N160), .ZN(N35225));
    INVX1 U22354 (.I(n20998), .ZN(n35226));
    INVX1 U22355 (.I(N11761), .ZN(N35227));
    NANDX1 U22356 (.A1(n17757), .A2(n24977), .ZN(N35228));
    NANDX1 U22357 (.A1(n24258), .A2(N5898), .ZN(n35229));
    INVX1 U22358 (.I(N6907), .ZN(N35230));
    INVX1 U22359 (.I(N6555), .ZN(n35231));
    INVX1 U22360 (.I(N7609), .ZN(N35232));
    INVX1 U22361 (.I(n19759), .ZN(n35233));
    NOR2X1 U22362 (.A1(N3810), .A2(n18456), .ZN(N35234));
    INVX1 U22363 (.I(N8871), .ZN(n35235));
    NANDX1 U22364 (.A1(N8116), .A2(N10895), .ZN(N35236));
    INVX1 U22365 (.I(N315), .ZN(N35237));
    INVX1 U22366 (.I(n13735), .ZN(n35238));
    NANDX1 U22367 (.A1(N6003), .A2(n23293), .ZN(N35239));
    NOR2X1 U22368 (.A1(n17764), .A2(n18620), .ZN(N35240));
    NANDX1 U22369 (.A1(N12603), .A2(N3739), .ZN(N35241));
    INVX1 U22370 (.I(N7061), .ZN(N35242));
    NOR2X1 U22371 (.A1(N10119), .A2(n17087), .ZN(n35243));
    NOR2X1 U22372 (.A1(N10109), .A2(n13256), .ZN(N35244));
    NOR2X1 U22373 (.A1(n18428), .A2(N8157), .ZN(n35245));
    NANDX1 U22374 (.A1(N6746), .A2(n22616), .ZN(N35246));
    NANDX1 U22375 (.A1(N8563), .A2(N594), .ZN(N35247));
    NOR2X1 U22376 (.A1(n14702), .A2(n19606), .ZN(N35248));
    INVX1 U22377 (.I(n28436), .ZN(N35249));
    NOR2X1 U22378 (.A1(N8869), .A2(n21592), .ZN(n35250));
    NOR2X1 U22379 (.A1(n15193), .A2(n28772), .ZN(n35251));
    INVX1 U22380 (.I(n16357), .ZN(N35252));
    NANDX1 U22381 (.A1(n16460), .A2(N11978), .ZN(N35253));
    NANDX1 U22382 (.A1(n26579), .A2(n17625), .ZN(N35254));
    INVX1 U22383 (.I(n25248), .ZN(n35255));
    INVX1 U22384 (.I(n19006), .ZN(N35256));
    NOR2X1 U22385 (.A1(N8899), .A2(n30051), .ZN(N35257));
    NANDX1 U22386 (.A1(n20076), .A2(n19828), .ZN(N35258));
    NOR2X1 U22387 (.A1(n20669), .A2(n20500), .ZN(N35259));
    INVX1 U22388 (.I(n28836), .ZN(N35260));
    NOR2X1 U22389 (.A1(n18968), .A2(n18778), .ZN(N35261));
    NANDX1 U22390 (.A1(n29120), .A2(N11494), .ZN(N35262));
    NOR2X1 U22391 (.A1(n27754), .A2(n13303), .ZN(N35263));
    NOR2X1 U22392 (.A1(n30126), .A2(n29762), .ZN(N35264));
    INVX1 U22393 (.I(N7413), .ZN(N35265));
    INVX1 U22394 (.I(N10233), .ZN(N35266));
    NOR2X1 U22395 (.A1(n28572), .A2(n29673), .ZN(N35267));
    INVX1 U22396 (.I(N11973), .ZN(N35268));
    INVX1 U22397 (.I(n26663), .ZN(N35269));
    NANDX1 U22398 (.A1(n17071), .A2(N4914), .ZN(n35270));
    NANDX1 U22399 (.A1(n26300), .A2(n13974), .ZN(n35271));
    NANDX1 U22400 (.A1(n24998), .A2(N7202), .ZN(n35272));
    INVX1 U22401 (.I(N2199), .ZN(n35273));
    INVX1 U22402 (.I(n23827), .ZN(n35274));
    NANDX1 U22403 (.A1(N10969), .A2(N10005), .ZN(N35275));
    NANDX1 U22404 (.A1(n21736), .A2(n28691), .ZN(n35276));
    NOR2X1 U22405 (.A1(N2904), .A2(N5966), .ZN(n35277));
    INVX1 U22406 (.I(N1697), .ZN(N35278));
    NANDX1 U22407 (.A1(N5500), .A2(N1233), .ZN(N35279));
    NANDX1 U22408 (.A1(n17472), .A2(n16926), .ZN(N35280));
    NOR2X1 U22409 (.A1(n26849), .A2(N3859), .ZN(N35281));
    NOR2X1 U22410 (.A1(N12057), .A2(N21), .ZN(N35282));
    NANDX1 U22411 (.A1(n17933), .A2(n25019), .ZN(N35283));
    NANDX1 U22412 (.A1(N12640), .A2(n27217), .ZN(N35284));
    NOR2X1 U22413 (.A1(n25028), .A2(n29470), .ZN(n35285));
    NANDX1 U22414 (.A1(n23593), .A2(N3449), .ZN(N35286));
    INVX1 U22415 (.I(n22146), .ZN(n35287));
    NANDX1 U22416 (.A1(n27904), .A2(n16673), .ZN(N35288));
    NOR2X1 U22417 (.A1(n18161), .A2(n18943), .ZN(N35289));
    INVX1 U22418 (.I(N7954), .ZN(N35290));
    INVX1 U22419 (.I(n25787), .ZN(N35291));
    NOR2X1 U22420 (.A1(n20491), .A2(N11059), .ZN(n35292));
    NOR2X1 U22421 (.A1(n28070), .A2(n23115), .ZN(n35293));
    NANDX1 U22422 (.A1(n19486), .A2(N10911), .ZN(n35294));
    NOR2X1 U22423 (.A1(N6665), .A2(N12111), .ZN(N35295));
    NANDX1 U22424 (.A1(N10400), .A2(n25699), .ZN(N35296));
    NANDX1 U22425 (.A1(n13665), .A2(n19154), .ZN(n35297));
    INVX1 U22426 (.I(N8527), .ZN(N35298));
    NANDX1 U22427 (.A1(n15069), .A2(n24991), .ZN(N35299));
    NOR2X1 U22428 (.A1(n29323), .A2(N1576), .ZN(N35300));
    NOR2X1 U22429 (.A1(N7501), .A2(N9529), .ZN(N35301));
    INVX1 U22430 (.I(n21848), .ZN(N35302));
    NANDX1 U22431 (.A1(N1939), .A2(N2769), .ZN(n35303));
    NANDX1 U22432 (.A1(n18569), .A2(n14445), .ZN(N35304));
    INVX1 U22433 (.I(n26616), .ZN(N35305));
    NANDX1 U22434 (.A1(N9509), .A2(N3143), .ZN(n35306));
    NOR2X1 U22435 (.A1(N7349), .A2(N2103), .ZN(n35307));
    NOR2X1 U22436 (.A1(n23219), .A2(n15767), .ZN(N35308));
    INVX1 U22437 (.I(N961), .ZN(N35309));
    NOR2X1 U22438 (.A1(n29025), .A2(n16030), .ZN(N35310));
    NOR2X1 U22439 (.A1(n15283), .A2(N3776), .ZN(N35311));
    NANDX1 U22440 (.A1(n20483), .A2(n29974), .ZN(n35312));
    INVX1 U22441 (.I(N1931), .ZN(N35313));
    NOR2X1 U22442 (.A1(n18902), .A2(n22567), .ZN(N35314));
    NOR2X1 U22443 (.A1(n29030), .A2(N10999), .ZN(N35315));
    NOR2X1 U22444 (.A1(n14901), .A2(N7477), .ZN(n35316));
    INVX1 U22445 (.I(n24409), .ZN(n35317));
    NOR2X1 U22446 (.A1(N7124), .A2(n20318), .ZN(N35318));
    NOR2X1 U22447 (.A1(n17272), .A2(N1960), .ZN(N35319));
    NOR2X1 U22448 (.A1(N4998), .A2(N2921), .ZN(n35320));
    NANDX1 U22449 (.A1(N3885), .A2(n18950), .ZN(N35321));
    NANDX1 U22450 (.A1(n19168), .A2(N11286), .ZN(N35322));
    NANDX1 U22451 (.A1(n28211), .A2(N11123), .ZN(N35323));
    NOR2X1 U22452 (.A1(N5), .A2(N2669), .ZN(N35324));
    NANDX1 U22453 (.A1(n22571), .A2(n15682), .ZN(n35325));
    NOR2X1 U22454 (.A1(n22130), .A2(n13002), .ZN(N35326));
    NANDX1 U22455 (.A1(n18167), .A2(n24237), .ZN(N35327));
    NANDX1 U22456 (.A1(N5907), .A2(n19922), .ZN(N35328));
    NANDX1 U22457 (.A1(n25887), .A2(n25754), .ZN(n35329));
    INVX1 U22458 (.I(N8618), .ZN(N35330));
    NOR2X1 U22459 (.A1(n14915), .A2(N4203), .ZN(N35331));
    INVX1 U22460 (.I(n22425), .ZN(N35332));
    INVX1 U22461 (.I(N788), .ZN(N35333));
    NOR2X1 U22462 (.A1(n27329), .A2(n28998), .ZN(N35334));
    INVX1 U22463 (.I(n24398), .ZN(n35335));
    NOR2X1 U22464 (.A1(N5925), .A2(N10231), .ZN(n35336));
    NOR2X1 U22465 (.A1(n21606), .A2(N2216), .ZN(N35337));
    NOR2X1 U22466 (.A1(n23169), .A2(n20539), .ZN(N35338));
    NANDX1 U22467 (.A1(n17268), .A2(n21695), .ZN(n35339));
    NANDX1 U22468 (.A1(n25750), .A2(n13032), .ZN(N35340));
    NANDX1 U22469 (.A1(n21367), .A2(n25026), .ZN(n35341));
    NOR2X1 U22470 (.A1(N10541), .A2(n28501), .ZN(N35342));
    NANDX1 U22471 (.A1(N3600), .A2(n20788), .ZN(N35343));
    INVX1 U22472 (.I(n23085), .ZN(N35344));
    INVX1 U22473 (.I(N4999), .ZN(N35345));
    INVX1 U22474 (.I(n27616), .ZN(N35346));
    NANDX1 U22475 (.A1(n28069), .A2(N3403), .ZN(n35347));
    NANDX1 U22476 (.A1(N7928), .A2(n25008), .ZN(n35348));
    NANDX1 U22477 (.A1(n28615), .A2(n18039), .ZN(N35349));
    NANDX1 U22478 (.A1(N7194), .A2(n23868), .ZN(N35350));
    INVX1 U22479 (.I(n21816), .ZN(N35351));
    NANDX1 U22480 (.A1(N2515), .A2(n20749), .ZN(N35352));
    NOR2X1 U22481 (.A1(n16101), .A2(n28298), .ZN(N35353));
    INVX1 U22482 (.I(n14464), .ZN(N35354));
    NANDX1 U22483 (.A1(N1971), .A2(n23812), .ZN(N35355));
    NANDX1 U22484 (.A1(n13617), .A2(n18035), .ZN(N35356));
    INVX1 U22485 (.I(n24123), .ZN(N35357));
    INVX1 U22486 (.I(n29236), .ZN(N35358));
    NOR2X1 U22487 (.A1(N7476), .A2(n15848), .ZN(N35359));
    INVX1 U22488 (.I(n21044), .ZN(n35360));
    NANDX1 U22489 (.A1(n17020), .A2(n27644), .ZN(n35361));
    NOR2X1 U22490 (.A1(N12774), .A2(n21374), .ZN(N35362));
    INVX1 U22491 (.I(n23150), .ZN(N35363));
    NANDX1 U22492 (.A1(N6037), .A2(N2322), .ZN(n35364));
    NANDX1 U22493 (.A1(n22138), .A2(n19181), .ZN(n35365));
    NOR2X1 U22494 (.A1(n25162), .A2(n17654), .ZN(N35366));
    NANDX1 U22495 (.A1(n18837), .A2(n23934), .ZN(n35367));
    NOR2X1 U22496 (.A1(n25432), .A2(n23773), .ZN(N35368));
    NANDX1 U22497 (.A1(n29505), .A2(N11433), .ZN(n35369));
    NOR2X1 U22498 (.A1(N6843), .A2(n27280), .ZN(N35370));
    NOR2X1 U22499 (.A1(n16447), .A2(N1816), .ZN(N35371));
    NOR2X1 U22500 (.A1(n13953), .A2(N4416), .ZN(n35372));
    NOR2X1 U22501 (.A1(n23887), .A2(N7938), .ZN(N35373));
    NOR2X1 U22502 (.A1(N11725), .A2(n13974), .ZN(N35374));
    NOR2X1 U22503 (.A1(N10271), .A2(n24672), .ZN(N35375));
    NANDX1 U22504 (.A1(n25886), .A2(n19697), .ZN(N35376));
    NANDX1 U22505 (.A1(N1895), .A2(N8396), .ZN(N35377));
    INVX1 U22506 (.I(n21658), .ZN(N35378));
    NOR2X1 U22507 (.A1(N9143), .A2(N5268), .ZN(N35379));
    NOR2X1 U22508 (.A1(N9136), .A2(N10932), .ZN(N35380));
    INVX1 U22509 (.I(N6278), .ZN(N35381));
    NOR2X1 U22510 (.A1(N3467), .A2(n26792), .ZN(n35382));
    NOR2X1 U22511 (.A1(N5981), .A2(N1070), .ZN(N35383));
    NANDX1 U22512 (.A1(n29867), .A2(n27705), .ZN(N35384));
    NOR2X1 U22513 (.A1(N11454), .A2(N11541), .ZN(N35385));
    NANDX1 U22514 (.A1(N10285), .A2(n24774), .ZN(N35386));
    NOR2X1 U22515 (.A1(n24731), .A2(n14333), .ZN(N35387));
    NANDX1 U22516 (.A1(n26626), .A2(N11289), .ZN(N35388));
    NOR2X1 U22517 (.A1(N6707), .A2(N3539), .ZN(N35389));
    NOR2X1 U22518 (.A1(N11974), .A2(n25293), .ZN(n35390));
    INVX1 U22519 (.I(n22906), .ZN(N35391));
    INVX1 U22520 (.I(N8762), .ZN(N35392));
    NOR2X1 U22521 (.A1(N4340), .A2(N5416), .ZN(n35393));
    INVX1 U22522 (.I(n29018), .ZN(N35394));
    NANDX1 U22523 (.A1(n26749), .A2(n17309), .ZN(N35395));
    INVX1 U22524 (.I(n26377), .ZN(N35396));
    NANDX1 U22525 (.A1(n22852), .A2(n22322), .ZN(n35397));
    NANDX1 U22526 (.A1(n17488), .A2(n22325), .ZN(N35398));
    NANDX1 U22527 (.A1(N1683), .A2(n13902), .ZN(N35399));
    INVX1 U22528 (.I(N1532), .ZN(N35400));
    INVX1 U22529 (.I(N2517), .ZN(N35401));
    INVX1 U22530 (.I(n14335), .ZN(N35402));
    NANDX1 U22531 (.A1(N225), .A2(n28258), .ZN(N35403));
    NANDX1 U22532 (.A1(N1098), .A2(N6882), .ZN(n35404));
    NANDX1 U22533 (.A1(n24135), .A2(N859), .ZN(n35405));
    NANDX1 U22534 (.A1(N11577), .A2(n26041), .ZN(N35406));
    NANDX1 U22535 (.A1(n28885), .A2(N7215), .ZN(N35407));
    INVX1 U22536 (.I(n16070), .ZN(N35408));
    NANDX1 U22537 (.A1(n18438), .A2(N2101), .ZN(N35409));
    NANDX1 U22538 (.A1(n29323), .A2(N12863), .ZN(n35410));
    NANDX1 U22539 (.A1(N1649), .A2(N8673), .ZN(N35411));
    NANDX1 U22540 (.A1(N11195), .A2(n29888), .ZN(n35412));
    NANDX1 U22541 (.A1(n25529), .A2(n14241), .ZN(N35413));
    NANDX1 U22542 (.A1(n23649), .A2(N10060), .ZN(N35414));
    NANDX1 U22543 (.A1(n19092), .A2(n22345), .ZN(N35415));
    NOR2X1 U22544 (.A1(n19950), .A2(N6912), .ZN(N35416));
    NOR2X1 U22545 (.A1(N4414), .A2(N6788), .ZN(N35417));
    INVX1 U22546 (.I(N11628), .ZN(N35418));
    NANDX1 U22547 (.A1(N1653), .A2(N117), .ZN(N35419));
    NOR2X1 U22548 (.A1(N3753), .A2(n17532), .ZN(n35420));
    INVX1 U22549 (.I(N5176), .ZN(n35421));
    NANDX1 U22550 (.A1(n29433), .A2(N2410), .ZN(N35422));
    INVX1 U22551 (.I(N10490), .ZN(N35423));
    NANDX1 U22552 (.A1(n14320), .A2(N5882), .ZN(N35424));
    INVX1 U22553 (.I(N5924), .ZN(N35425));
    NOR2X1 U22554 (.A1(N3581), .A2(n28762), .ZN(n35426));
    INVX1 U22555 (.I(n25925), .ZN(N35427));
    INVX1 U22556 (.I(N4116), .ZN(N35428));
    NOR2X1 U22557 (.A1(n28253), .A2(N8530), .ZN(N35429));
    INVX1 U22558 (.I(n13836), .ZN(n35430));
    NANDX1 U22559 (.A1(N8209), .A2(N4049), .ZN(N35431));
    INVX1 U22560 (.I(N6670), .ZN(n35432));
    NANDX1 U22561 (.A1(n14927), .A2(N4317), .ZN(N35433));
    NANDX1 U22562 (.A1(n28678), .A2(n22310), .ZN(n35434));
    INVX1 U22563 (.I(n28739), .ZN(N35435));
    NOR2X1 U22564 (.A1(n24804), .A2(n12922), .ZN(N35436));
    NANDX1 U22565 (.A1(n18325), .A2(n18845), .ZN(n35437));
    NANDX1 U22566 (.A1(n21905), .A2(N6031), .ZN(N35438));
    NOR2X1 U22567 (.A1(n17692), .A2(n17311), .ZN(N35439));
    NANDX1 U22568 (.A1(N8952), .A2(n15426), .ZN(N35440));
    INVX1 U22569 (.I(n25696), .ZN(N35441));
    NANDX1 U22570 (.A1(n27983), .A2(n22465), .ZN(N35442));
    NANDX1 U22571 (.A1(n25378), .A2(n29135), .ZN(N35443));
    INVX1 U22572 (.I(N10167), .ZN(N35444));
    NANDX1 U22573 (.A1(N8330), .A2(n27405), .ZN(N35445));
    NANDX1 U22574 (.A1(N837), .A2(n26007), .ZN(N35446));
    NANDX1 U22575 (.A1(n14201), .A2(n27489), .ZN(n35447));
    NOR2X1 U22576 (.A1(N2388), .A2(N4757), .ZN(N35448));
    INVX1 U22577 (.I(n24292), .ZN(N35449));
    INVX1 U22578 (.I(N8707), .ZN(n35450));
    NANDX1 U22579 (.A1(n16658), .A2(n19443), .ZN(n35451));
    NANDX1 U22580 (.A1(N1947), .A2(N8570), .ZN(n35452));
    INVX1 U22581 (.I(N1070), .ZN(N35453));
    INVX1 U22582 (.I(n15942), .ZN(n35454));
    INVX1 U22583 (.I(n20353), .ZN(n35455));
    NOR2X1 U22584 (.A1(n18293), .A2(n19081), .ZN(N35456));
    NOR2X1 U22585 (.A1(n26622), .A2(N4909), .ZN(N35457));
    NANDX1 U22586 (.A1(n16019), .A2(n19476), .ZN(N35458));
    NOR2X1 U22587 (.A1(N82), .A2(n16827), .ZN(N35459));
    NANDX1 U22588 (.A1(n21167), .A2(N10145), .ZN(N35460));
    NOR2X1 U22589 (.A1(n15321), .A2(n20931), .ZN(n35461));
    INVX1 U22590 (.I(n15727), .ZN(n35462));
    INVX1 U22591 (.I(n20654), .ZN(N35463));
    INVX1 U22592 (.I(n28096), .ZN(N35464));
    NANDX1 U22593 (.A1(N7123), .A2(n17726), .ZN(n35465));
    NOR2X1 U22594 (.A1(N11625), .A2(n29226), .ZN(n35466));
    INVX1 U22595 (.I(n15125), .ZN(N35467));
    NOR2X1 U22596 (.A1(n29314), .A2(N10499), .ZN(N35468));
    INVX1 U22597 (.I(N4086), .ZN(N35469));
    NOR2X1 U22598 (.A1(n18444), .A2(N12122), .ZN(N35470));
    NANDX1 U22599 (.A1(N7086), .A2(n28949), .ZN(N35471));
    INVX1 U22600 (.I(n28252), .ZN(N35472));
    NANDX1 U22601 (.A1(n13764), .A2(N1996), .ZN(n35473));
    INVX1 U22602 (.I(N3536), .ZN(N35474));
    NOR2X1 U22603 (.A1(n14459), .A2(n24189), .ZN(n35475));
    INVX1 U22604 (.I(N12417), .ZN(N35476));
    NOR2X1 U22605 (.A1(n27051), .A2(N6), .ZN(N35477));
    NOR2X1 U22606 (.A1(n27236), .A2(n17792), .ZN(n35478));
    INVX1 U22607 (.I(N12223), .ZN(N35479));
    NOR2X1 U22608 (.A1(N11127), .A2(N11282), .ZN(n35480));
    NOR2X1 U22609 (.A1(N3773), .A2(n19899), .ZN(N35481));
    NANDX1 U22610 (.A1(n15894), .A2(N9164), .ZN(N35482));
    INVX1 U22611 (.I(N3266), .ZN(n35483));
    NOR2X1 U22612 (.A1(N8227), .A2(N12221), .ZN(n35484));
    NOR2X1 U22613 (.A1(N10222), .A2(n19229), .ZN(N35485));
    INVX1 U22614 (.I(n16505), .ZN(N35486));
    NOR2X1 U22615 (.A1(n18896), .A2(N6296), .ZN(n35487));
    NOR2X1 U22616 (.A1(n19292), .A2(n21907), .ZN(N35488));
    INVX1 U22617 (.I(n21008), .ZN(n35489));
    NOR2X1 U22618 (.A1(n29583), .A2(n14259), .ZN(N35490));
    INVX1 U22619 (.I(n23179), .ZN(n35491));
    INVX1 U22620 (.I(N934), .ZN(N35492));
    INVX1 U22621 (.I(n17718), .ZN(n35493));
    NANDX1 U22622 (.A1(N3529), .A2(N3475), .ZN(n35494));
    NANDX1 U22623 (.A1(n13640), .A2(N6740), .ZN(N35495));
    INVX1 U22624 (.I(N10427), .ZN(N35496));
    NOR2X1 U22625 (.A1(n28711), .A2(n20649), .ZN(N35497));
    INVX1 U22626 (.I(n23418), .ZN(N35498));
    INVX1 U22627 (.I(N7421), .ZN(N35499));
    INVX1 U22628 (.I(n13312), .ZN(N35500));
    NOR2X1 U22629 (.A1(n20028), .A2(N5081), .ZN(N35501));
    NOR2X1 U22630 (.A1(N10898), .A2(N12647), .ZN(N35502));
    INVX1 U22631 (.I(n13717), .ZN(N35503));
    NOR2X1 U22632 (.A1(N12046), .A2(n27663), .ZN(N35504));
    NOR2X1 U22633 (.A1(N1109), .A2(n15243), .ZN(n35505));
    INVX1 U22634 (.I(n23335), .ZN(n35506));
    NANDX1 U22635 (.A1(N1043), .A2(n25536), .ZN(N35507));
    NOR2X1 U22636 (.A1(N8446), .A2(n24523), .ZN(N35508));
    NANDX1 U22637 (.A1(n25717), .A2(n15034), .ZN(n35509));
    NANDX1 U22638 (.A1(N7558), .A2(N10611), .ZN(n35510));
    INVX1 U22639 (.I(N8294), .ZN(N35511));
    NANDX1 U22640 (.A1(n21900), .A2(n16882), .ZN(N35512));
    INVX1 U22641 (.I(n22760), .ZN(N35513));
    NOR2X1 U22642 (.A1(n18771), .A2(N11627), .ZN(N35514));
    NANDX1 U22643 (.A1(n21069), .A2(N12234), .ZN(n35515));
    NOR2X1 U22644 (.A1(n24300), .A2(N1903), .ZN(N35516));
    NOR2X1 U22645 (.A1(N6786), .A2(n13799), .ZN(N35517));
    NANDX1 U22646 (.A1(N7829), .A2(n27895), .ZN(n35518));
    INVX1 U22647 (.I(N4835), .ZN(N35519));
    NANDX1 U22648 (.A1(N2505), .A2(N414), .ZN(n35520));
    NOR2X1 U22649 (.A1(N9216), .A2(N7972), .ZN(N35521));
    INVX1 U22650 (.I(N11908), .ZN(N35522));
    INVX1 U22651 (.I(n18830), .ZN(n35523));
    NOR2X1 U22652 (.A1(n21708), .A2(n24953), .ZN(N35524));
    NANDX1 U22653 (.A1(N7910), .A2(n13586), .ZN(N35525));
    NANDX1 U22654 (.A1(n26527), .A2(n23215), .ZN(N35526));
    INVX1 U22655 (.I(N12532), .ZN(N35527));
    NANDX1 U22656 (.A1(n29314), .A2(N2341), .ZN(n35528));
    NANDX1 U22657 (.A1(N1536), .A2(n29564), .ZN(N35529));
    INVX1 U22658 (.I(n29430), .ZN(N35530));
    INVX1 U22659 (.I(n25386), .ZN(N35531));
    INVX1 U22660 (.I(n13034), .ZN(N35532));
    NOR2X1 U22661 (.A1(n17309), .A2(N10810), .ZN(N35533));
    NOR2X1 U22662 (.A1(N12217), .A2(n22717), .ZN(N35534));
    INVX1 U22663 (.I(N909), .ZN(n35535));
    NANDX1 U22664 (.A1(N7288), .A2(n14423), .ZN(N35536));
    NOR2X1 U22665 (.A1(n15197), .A2(n16569), .ZN(n35537));
    NANDX1 U22666 (.A1(N11587), .A2(N9647), .ZN(N35538));
    INVX1 U22667 (.I(n24118), .ZN(n35539));
    NOR2X1 U22668 (.A1(N11428), .A2(n15019), .ZN(n35540));
    INVX1 U22669 (.I(n12963), .ZN(n35541));
    NOR2X1 U22670 (.A1(N23), .A2(N816), .ZN(N35542));
    INVX1 U22671 (.I(n25408), .ZN(n35543));
    INVX1 U22672 (.I(n26568), .ZN(N35544));
    INVX1 U22673 (.I(n28257), .ZN(N35545));
    NOR2X1 U22674 (.A1(N1824), .A2(N10336), .ZN(n35546));
    NOR2X1 U22675 (.A1(n17541), .A2(N11245), .ZN(N35547));
    NANDX1 U22676 (.A1(n24828), .A2(n14228), .ZN(N35548));
    INVX1 U22677 (.I(n28586), .ZN(N35549));
    NANDX1 U22678 (.A1(n29544), .A2(N10035), .ZN(N35550));
    NOR2X1 U22679 (.A1(N11658), .A2(n22713), .ZN(N35551));
    NOR2X1 U22680 (.A1(N11646), .A2(n26293), .ZN(n35552));
    NOR2X1 U22681 (.A1(n13169), .A2(n29298), .ZN(N35553));
    NOR2X1 U22682 (.A1(n13984), .A2(N12696), .ZN(N35554));
    NANDX1 U22683 (.A1(N6234), .A2(n27824), .ZN(N35555));
    NANDX1 U22684 (.A1(N4353), .A2(n23625), .ZN(n35556));
    NANDX1 U22685 (.A1(N3249), .A2(N12005), .ZN(N35557));
    NOR2X1 U22686 (.A1(n14493), .A2(n15332), .ZN(N35558));
    NOR2X1 U22687 (.A1(n17281), .A2(n18459), .ZN(n35559));
    NOR2X1 U22688 (.A1(n17940), .A2(N6426), .ZN(N35560));
    NOR2X1 U22689 (.A1(n16805), .A2(n18084), .ZN(N35561));
    NANDX1 U22690 (.A1(n19815), .A2(n18290), .ZN(n35562));
    INVX1 U22691 (.I(N2297), .ZN(N35563));
    NOR2X1 U22692 (.A1(N12351), .A2(n14938), .ZN(N35564));
    NOR2X1 U22693 (.A1(n25046), .A2(n22849), .ZN(N35565));
    NANDX1 U22694 (.A1(n22732), .A2(N10254), .ZN(n35566));
    NANDX1 U22695 (.A1(n16219), .A2(n18180), .ZN(N35567));
    INVX1 U22696 (.I(n16784), .ZN(n35568));
    NANDX1 U22697 (.A1(N9314), .A2(N1978), .ZN(N35569));
    INVX1 U22698 (.I(n26595), .ZN(N35570));
    NOR2X1 U22699 (.A1(n17954), .A2(N2958), .ZN(N35571));
    NANDX1 U22700 (.A1(n23715), .A2(N8323), .ZN(n35572));
    INVX1 U22701 (.I(N10613), .ZN(N35573));
    NOR2X1 U22702 (.A1(N10219), .A2(n23802), .ZN(N35574));
    NOR2X1 U22703 (.A1(N101), .A2(n24713), .ZN(N35575));
    NANDX1 U22704 (.A1(N3967), .A2(n19621), .ZN(N35576));
    NANDX1 U22705 (.A1(n14065), .A2(N777), .ZN(N35577));
    NANDX1 U22706 (.A1(n17077), .A2(N5556), .ZN(N35578));
    INVX1 U22707 (.I(N11898), .ZN(N35579));
    INVX1 U22708 (.I(n15569), .ZN(n35580));
    NOR2X1 U22709 (.A1(n12878), .A2(n26356), .ZN(n35581));
    INVX1 U22710 (.I(n21875), .ZN(N35582));
    INVX1 U22711 (.I(n20625), .ZN(N35583));
    NOR2X1 U22712 (.A1(n15009), .A2(n17509), .ZN(N35584));
    NOR2X1 U22713 (.A1(n14182), .A2(n15509), .ZN(N35585));
    NANDX1 U22714 (.A1(n26545), .A2(n15805), .ZN(N35586));
    INVX1 U22715 (.I(n21120), .ZN(N35587));
    INVX1 U22716 (.I(N1935), .ZN(N35588));
    INVX1 U22717 (.I(n16104), .ZN(N35589));
    INVX1 U22718 (.I(n30078), .ZN(n35590));
    NANDX1 U22719 (.A1(N10197), .A2(n24194), .ZN(N35591));
    NANDX1 U22720 (.A1(n22094), .A2(n16396), .ZN(N35592));
    NANDX1 U22721 (.A1(N1729), .A2(n29274), .ZN(N35593));
    NOR2X1 U22722 (.A1(N7957), .A2(n21011), .ZN(N35594));
    NOR2X1 U22723 (.A1(n17143), .A2(n16731), .ZN(N35595));
    NOR2X1 U22724 (.A1(N4514), .A2(N4380), .ZN(N35596));
    NANDX1 U22725 (.A1(n20022), .A2(N2247), .ZN(n35597));
    INVX1 U22726 (.I(n24387), .ZN(N35598));
    INVX1 U22727 (.I(N10265), .ZN(n35599));
    NANDX1 U22728 (.A1(N9408), .A2(N9429), .ZN(N35600));
    INVX1 U22729 (.I(N2529), .ZN(N35601));
    NOR2X1 U22730 (.A1(N11237), .A2(N12725), .ZN(n35602));
    NANDX1 U22731 (.A1(N6022), .A2(n23380), .ZN(N35603));
    NOR2X1 U22732 (.A1(n16374), .A2(n25108), .ZN(N35604));
    INVX1 U22733 (.I(N11506), .ZN(N35605));
    NANDX1 U22734 (.A1(n17089), .A2(n28069), .ZN(N35606));
    NANDX1 U22735 (.A1(N3682), .A2(n29504), .ZN(n35607));
    NOR2X1 U22736 (.A1(N8061), .A2(N3544), .ZN(N35608));
    NANDX1 U22737 (.A1(n29006), .A2(n22826), .ZN(N35609));
    INVX1 U22738 (.I(N6342), .ZN(n35610));
    NOR2X1 U22739 (.A1(n29821), .A2(n15750), .ZN(N35611));
    NANDX1 U22740 (.A1(n18196), .A2(N6839), .ZN(N35612));
    INVX1 U22741 (.I(n29432), .ZN(N35613));
    NOR2X1 U22742 (.A1(N9556), .A2(N5316), .ZN(n35614));
    INVX1 U22743 (.I(N6499), .ZN(N35615));
    NOR2X1 U22744 (.A1(n26473), .A2(N2577), .ZN(n35616));
    NOR2X1 U22745 (.A1(n17961), .A2(n19666), .ZN(n35617));
    NOR2X1 U22746 (.A1(n26590), .A2(N11908), .ZN(N35618));
    NOR2X1 U22747 (.A1(N9596), .A2(N8530), .ZN(N35619));
    INVX1 U22748 (.I(N12622), .ZN(N35620));
    INVX1 U22749 (.I(n22544), .ZN(N35621));
    NANDX1 U22750 (.A1(N2300), .A2(n25496), .ZN(n35622));
    INVX1 U22751 (.I(N6610), .ZN(N35623));
    INVX1 U22752 (.I(N4898), .ZN(N35624));
    INVX1 U22753 (.I(n13871), .ZN(N35625));
    NANDX1 U22754 (.A1(n21572), .A2(n23426), .ZN(N35626));
    NOR2X1 U22755 (.A1(n22937), .A2(n29924), .ZN(N35627));
    NOR2X1 U22756 (.A1(n19273), .A2(n21062), .ZN(n35628));
    INVX1 U22757 (.I(n25794), .ZN(N35629));
    NOR2X1 U22758 (.A1(N8186), .A2(n22246), .ZN(N35630));
    NOR2X1 U22759 (.A1(N4361), .A2(N1704), .ZN(N35631));
    NANDX1 U22760 (.A1(N4079), .A2(N2887), .ZN(N35632));
    NANDX1 U22761 (.A1(n26622), .A2(n20043), .ZN(N35633));
    NOR2X1 U22762 (.A1(n21980), .A2(N6745), .ZN(n35634));
    INVX1 U22763 (.I(N6842), .ZN(N35635));
    NOR2X1 U22764 (.A1(n22283), .A2(N9273), .ZN(n35636));
    NANDX1 U22765 (.A1(n13717), .A2(N2561), .ZN(N35637));
    NANDX1 U22766 (.A1(n25214), .A2(n21046), .ZN(n35638));
    NANDX1 U22767 (.A1(n14349), .A2(N11970), .ZN(n35639));
    NOR2X1 U22768 (.A1(n28703), .A2(N11120), .ZN(n35640));
    NANDX1 U22769 (.A1(n20812), .A2(N10738), .ZN(n35641));
    INVX1 U22770 (.I(n22515), .ZN(N35642));
    NANDX1 U22771 (.A1(N285), .A2(n13962), .ZN(N35643));
    INVX1 U22772 (.I(n15467), .ZN(n35644));
    NANDX1 U22773 (.A1(n25216), .A2(N7309), .ZN(N35645));
    INVX1 U22774 (.I(N3914), .ZN(n35646));
    NOR2X1 U22775 (.A1(n18074), .A2(n26196), .ZN(N35647));
    INVX1 U22776 (.I(n29728), .ZN(n35648));
    NANDX1 U22777 (.A1(N3105), .A2(n28011), .ZN(N35649));
    NANDX1 U22778 (.A1(n24150), .A2(n23174), .ZN(N35650));
    INVX1 U22779 (.I(n24680), .ZN(n35651));
    INVX1 U22780 (.I(N6326), .ZN(N35652));
    NOR2X1 U22781 (.A1(n17379), .A2(n15698), .ZN(N35653));
    NOR2X1 U22782 (.A1(n13585), .A2(N8076), .ZN(n35654));
    NANDX1 U22783 (.A1(N2430), .A2(N10598), .ZN(N35655));
    INVX1 U22784 (.I(n17896), .ZN(n35656));
    NANDX1 U22785 (.A1(N7597), .A2(n13766), .ZN(n35657));
    NANDX1 U22786 (.A1(N71), .A2(N5037), .ZN(n35658));
    NOR2X1 U22787 (.A1(n26266), .A2(n17020), .ZN(N35659));
    INVX1 U22788 (.I(n24601), .ZN(n35660));
    INVX1 U22789 (.I(n17734), .ZN(N35661));
    INVX1 U22790 (.I(N2697), .ZN(n35662));
    NANDX1 U22791 (.A1(n14334), .A2(n15937), .ZN(N35663));
    NANDX1 U22792 (.A1(N9220), .A2(N10159), .ZN(n35664));
    NANDX1 U22793 (.A1(n24918), .A2(n15118), .ZN(N35665));
    NANDX1 U22794 (.A1(n21554), .A2(n27524), .ZN(N35666));
    INVX1 U22795 (.I(N2014), .ZN(n35667));
    INVX1 U22796 (.I(N4439), .ZN(N35668));
    NANDX1 U22797 (.A1(n24760), .A2(N6765), .ZN(N35669));
    NOR2X1 U22798 (.A1(n24831), .A2(N11802), .ZN(N35670));
    NOR2X1 U22799 (.A1(n20959), .A2(n28821), .ZN(n35671));
    NOR2X1 U22800 (.A1(n15423), .A2(N7368), .ZN(N35672));
    NOR2X1 U22801 (.A1(N3298), .A2(n28762), .ZN(n35673));
    NANDX1 U22802 (.A1(N6192), .A2(N3122), .ZN(N35674));
    INVX1 U22803 (.I(n15411), .ZN(N35675));
    INVX1 U22804 (.I(N3729), .ZN(N35676));
    INVX1 U22805 (.I(n28397), .ZN(N35677));
    NOR2X1 U22806 (.A1(N1607), .A2(n14344), .ZN(N35678));
    NOR2X1 U22807 (.A1(N3621), .A2(N12809), .ZN(n35679));
    NOR2X1 U22808 (.A1(N8659), .A2(N7432), .ZN(N35680));
    INVX1 U22809 (.I(n15895), .ZN(N35681));
    NANDX1 U22810 (.A1(N8829), .A2(n13263), .ZN(N35682));
    NOR2X1 U22811 (.A1(n26210), .A2(n19053), .ZN(n35683));
    NANDX1 U22812 (.A1(n22138), .A2(N12439), .ZN(N35684));
    NOR2X1 U22813 (.A1(N9323), .A2(n16595), .ZN(n35685));
    INVX1 U22814 (.I(N12444), .ZN(n35686));
    NANDX1 U22815 (.A1(n29087), .A2(n25723), .ZN(N35687));
    NANDX1 U22816 (.A1(N9140), .A2(N12543), .ZN(n35688));
    INVX1 U22817 (.I(N10747), .ZN(n35689));
    NANDX1 U22818 (.A1(N4311), .A2(N2928), .ZN(N35690));
    NOR2X1 U22819 (.A1(n13271), .A2(N147), .ZN(N35691));
    NOR2X1 U22820 (.A1(N10298), .A2(N4602), .ZN(N35692));
    NANDX1 U22821 (.A1(N7687), .A2(N6426), .ZN(n35693));
    NANDX1 U22822 (.A1(n22457), .A2(n25478), .ZN(N35694));
    NOR2X1 U22823 (.A1(N3018), .A2(N7779), .ZN(N35695));
    INVX1 U22824 (.I(N12340), .ZN(n35696));
    NOR2X1 U22825 (.A1(n21787), .A2(n13344), .ZN(N35697));
    INVX1 U22826 (.I(n20736), .ZN(N35698));
    INVX1 U22827 (.I(N6039), .ZN(n35699));
    NOR2X1 U22828 (.A1(n28731), .A2(n13086), .ZN(N35700));
    INVX1 U22829 (.I(n14041), .ZN(N35701));
    NANDX1 U22830 (.A1(n20671), .A2(n19418), .ZN(N35702));
    NOR2X1 U22831 (.A1(n20817), .A2(N2090), .ZN(N35703));
    INVX1 U22832 (.I(n13980), .ZN(N35704));
    INVX1 U22833 (.I(n14334), .ZN(N35705));
    NANDX1 U22834 (.A1(N9281), .A2(N6653), .ZN(n35706));
    INVX1 U22835 (.I(N9908), .ZN(N35707));
    INVX1 U22836 (.I(N12084), .ZN(n35708));
    INVX1 U22837 (.I(N10571), .ZN(n35709));
    NANDX1 U22838 (.A1(n16927), .A2(N12476), .ZN(N35710));
    NOR2X1 U22839 (.A1(N7526), .A2(N9965), .ZN(N35711));
    NOR2X1 U22840 (.A1(n25962), .A2(n27256), .ZN(n35712));
    NOR2X1 U22841 (.A1(n13568), .A2(N11159), .ZN(n35713));
    NANDX1 U22842 (.A1(n22799), .A2(n19138), .ZN(n35714));
    INVX1 U22843 (.I(n13478), .ZN(N35715));
    NANDX1 U22844 (.A1(N2530), .A2(n16018), .ZN(N35716));
    NOR2X1 U22845 (.A1(n16863), .A2(N6285), .ZN(n35717));
    NOR2X1 U22846 (.A1(n23516), .A2(N10590), .ZN(N35718));
    NOR2X1 U22847 (.A1(n21747), .A2(n22673), .ZN(n35719));
    NOR2X1 U22848 (.A1(n20878), .A2(N6113), .ZN(N35720));
    NANDX1 U22849 (.A1(N3216), .A2(n17963), .ZN(N35721));
    INVX1 U22850 (.I(N1742), .ZN(N35722));
    NOR2X1 U22851 (.A1(n15656), .A2(n28997), .ZN(N35723));
    NOR2X1 U22852 (.A1(n29223), .A2(n28717), .ZN(N35724));
    INVX1 U22853 (.I(n21884), .ZN(N35725));
    NANDX1 U22854 (.A1(n16485), .A2(n23923), .ZN(N35726));
    INVX1 U22855 (.I(n19015), .ZN(n35727));
    INVX1 U22856 (.I(N12736), .ZN(N35728));
    NOR2X1 U22857 (.A1(N4649), .A2(N7249), .ZN(n35729));
    NOR2X1 U22858 (.A1(n15238), .A2(n18928), .ZN(n35730));
    INVX1 U22859 (.I(n26472), .ZN(N35731));
    NANDX1 U22860 (.A1(n18864), .A2(N2447), .ZN(N35732));
    INVX1 U22861 (.I(N10640), .ZN(n35733));
    NOR2X1 U22862 (.A1(n13230), .A2(N942), .ZN(N35734));
    NOR2X1 U22863 (.A1(n28886), .A2(n18500), .ZN(N35735));
    NOR2X1 U22864 (.A1(n16532), .A2(n17079), .ZN(n35736));
    INVX1 U22865 (.I(n26977), .ZN(N35737));
    NANDX1 U22866 (.A1(n16743), .A2(n20762), .ZN(n35738));
    NANDX1 U22867 (.A1(N5620), .A2(n19125), .ZN(N35739));
    NANDX1 U22868 (.A1(N11359), .A2(n23773), .ZN(N35740));
    NANDX1 U22869 (.A1(n29175), .A2(N8874), .ZN(n35741));
    NOR2X1 U22870 (.A1(n27160), .A2(N5208), .ZN(n35742));
    NANDX1 U22871 (.A1(N4447), .A2(n26352), .ZN(N35743));
    NOR2X1 U22872 (.A1(N3648), .A2(N5185), .ZN(n35744));
    NOR2X1 U22873 (.A1(N4589), .A2(N8428), .ZN(N35745));
    INVX1 U22874 (.I(N11649), .ZN(n35746));
    NANDX1 U22875 (.A1(N1257), .A2(n28727), .ZN(N35747));
    INVX1 U22876 (.I(n28233), .ZN(n35748));
    NOR2X1 U22877 (.A1(n23782), .A2(N7418), .ZN(N35749));
    NANDX1 U22878 (.A1(n29401), .A2(n15103), .ZN(n35750));
    INVX1 U22879 (.I(n29320), .ZN(N35751));
    INVX1 U22880 (.I(n29496), .ZN(N35752));
    NANDX1 U22881 (.A1(N6173), .A2(N5976), .ZN(n35753));
    NANDX1 U22882 (.A1(n30078), .A2(N8203), .ZN(N35754));
    INVX1 U22883 (.I(n26292), .ZN(N35755));
    NANDX1 U22884 (.A1(n29293), .A2(n20037), .ZN(N35756));
    NOR2X1 U22885 (.A1(N3745), .A2(n28465), .ZN(N35757));
    NOR2X1 U22886 (.A1(N3954), .A2(N5109), .ZN(N35758));
    INVX1 U22887 (.I(n21242), .ZN(N35759));
    NOR2X1 U22888 (.A1(n29974), .A2(N1610), .ZN(N35760));
    NANDX1 U22889 (.A1(n25952), .A2(n21398), .ZN(n35761));
    INVX1 U22890 (.I(N10918), .ZN(N35762));
    NOR2X1 U22891 (.A1(n22936), .A2(N8217), .ZN(n35763));
    NANDX1 U22892 (.A1(N9716), .A2(n14389), .ZN(N35764));
    NOR2X1 U22893 (.A1(N12217), .A2(N2890), .ZN(n35765));
    NOR2X1 U22894 (.A1(n19165), .A2(n17742), .ZN(N35766));
    INVX1 U22895 (.I(n18320), .ZN(N35767));
    NANDX1 U22896 (.A1(n13175), .A2(N10625), .ZN(N35768));
    NOR2X1 U22897 (.A1(N6402), .A2(n14579), .ZN(N35769));
    NANDX1 U22898 (.A1(N8143), .A2(N5683), .ZN(N35770));
    NOR2X1 U22899 (.A1(N7980), .A2(n25990), .ZN(N35771));
    INVX1 U22900 (.I(N3794), .ZN(n35772));
    NOR2X1 U22901 (.A1(n18452), .A2(n14711), .ZN(n35773));
    NOR2X1 U22902 (.A1(N11250), .A2(N11488), .ZN(n35774));
    INVX1 U22903 (.I(N9526), .ZN(n35775));
    NANDX1 U22904 (.A1(N3668), .A2(n21743), .ZN(N35776));
    INVX1 U22905 (.I(n27391), .ZN(N35777));
    NOR2X1 U22906 (.A1(N4931), .A2(N1926), .ZN(n35778));
    NOR2X1 U22907 (.A1(N12572), .A2(N3662), .ZN(N35779));
    NANDX1 U22908 (.A1(N7101), .A2(N10063), .ZN(n35780));
    NOR2X1 U22909 (.A1(n25436), .A2(n18205), .ZN(N35781));
    INVX1 U22910 (.I(n25782), .ZN(N35782));
    NOR2X1 U22911 (.A1(n28768), .A2(n20481), .ZN(n35783));
    NANDX1 U22912 (.A1(N4442), .A2(N8795), .ZN(n35784));
    NANDX1 U22913 (.A1(N1741), .A2(n20044), .ZN(N35785));
    NANDX1 U22914 (.A1(n20025), .A2(n29569), .ZN(N35786));
    INVX1 U22915 (.I(N12253), .ZN(n35787));
    NANDX1 U22916 (.A1(N4786), .A2(n28204), .ZN(n35788));
    INVX1 U22917 (.I(N9716), .ZN(n35789));
    NOR2X1 U22918 (.A1(n15276), .A2(N10848), .ZN(n35790));
    NANDX1 U22919 (.A1(n20672), .A2(N6509), .ZN(N35791));
    INVX1 U22920 (.I(n29207), .ZN(n35792));
    INVX1 U22921 (.I(N9042), .ZN(N35793));
    NANDX1 U22922 (.A1(n27589), .A2(n23786), .ZN(n35794));
    NOR2X1 U22923 (.A1(n17932), .A2(N748), .ZN(N35795));
    NOR2X1 U22924 (.A1(n15287), .A2(N11119), .ZN(N35796));
    INVX1 U22925 (.I(N5193), .ZN(N35797));
    NOR2X1 U22926 (.A1(n22504), .A2(n23322), .ZN(N35798));
    INVX1 U22927 (.I(N4619), .ZN(N35799));
    NOR2X1 U22928 (.A1(n13782), .A2(N2685), .ZN(N35800));
    INVX1 U22929 (.I(N12058), .ZN(N35801));
    NOR2X1 U22930 (.A1(n15820), .A2(n22905), .ZN(N35802));
    NOR2X1 U22931 (.A1(n25052), .A2(n29413), .ZN(N35803));
    INVX1 U22932 (.I(N12682), .ZN(N35804));
    NANDX1 U22933 (.A1(N2026), .A2(N3090), .ZN(N35805));
    INVX1 U22934 (.I(n14373), .ZN(N35806));
    NOR2X1 U22935 (.A1(n23724), .A2(N3681), .ZN(N35807));
    NANDX1 U22936 (.A1(N8873), .A2(N3360), .ZN(N35808));
    NOR2X1 U22937 (.A1(N2626), .A2(n24897), .ZN(n35809));
    INVX1 U22938 (.I(n14508), .ZN(n35810));
    NOR2X1 U22939 (.A1(n15208), .A2(N5988), .ZN(N35811));
    NOR2X1 U22940 (.A1(N6453), .A2(N6533), .ZN(n35812));
    NANDX1 U22941 (.A1(n16388), .A2(N10913), .ZN(n35813));
    NOR2X1 U22942 (.A1(n18536), .A2(N5828), .ZN(N35814));
    INVX1 U22943 (.I(N11520), .ZN(N35815));
    NANDX1 U22944 (.A1(N7102), .A2(N2107), .ZN(N35816));
    NANDX1 U22945 (.A1(N1455), .A2(N5040), .ZN(n35817));
    INVX1 U22946 (.I(n25178), .ZN(N35818));
    NANDX1 U22947 (.A1(N6593), .A2(n22611), .ZN(n35819));
    NANDX1 U22948 (.A1(n24817), .A2(n13797), .ZN(N35820));
    NOR2X1 U22949 (.A1(N5269), .A2(n16865), .ZN(N35821));
    NANDX1 U22950 (.A1(N9038), .A2(n22853), .ZN(N35822));
    NANDX1 U22951 (.A1(N4051), .A2(n29385), .ZN(N35823));
    INVX1 U22952 (.I(n20438), .ZN(n35824));
    NANDX1 U22953 (.A1(N17), .A2(n27534), .ZN(n35825));
    NOR2X1 U22954 (.A1(n17475), .A2(n27615), .ZN(n35826));
    NANDX1 U22955 (.A1(n13137), .A2(n18282), .ZN(n35827));
    NOR2X1 U22956 (.A1(n14591), .A2(n23321), .ZN(N35828));
    INVX1 U22957 (.I(n28329), .ZN(n35829));
    NANDX1 U22958 (.A1(N7778), .A2(N9363), .ZN(n35830));
    NOR2X1 U22959 (.A1(n21155), .A2(N11720), .ZN(N35831));
    NOR2X1 U22960 (.A1(n14985), .A2(n28585), .ZN(N35832));
    NANDX1 U22961 (.A1(N12583), .A2(n21300), .ZN(N35833));
    INVX1 U22962 (.I(n16633), .ZN(n35834));
    NANDX1 U22963 (.A1(N10143), .A2(n25632), .ZN(N35835));
    NOR2X1 U22964 (.A1(N10160), .A2(N11589), .ZN(N35836));
    NOR2X1 U22965 (.A1(n16195), .A2(N9066), .ZN(N35837));
    NANDX1 U22966 (.A1(n29332), .A2(n27347), .ZN(N35838));
    INVX1 U22967 (.I(N2346), .ZN(n35839));
    NANDX1 U22968 (.A1(n19896), .A2(N538), .ZN(N35840));
    INVX1 U22969 (.I(n16234), .ZN(N35841));
    NOR2X1 U22970 (.A1(N9356), .A2(N7252), .ZN(N35842));
    NOR2X1 U22971 (.A1(n14557), .A2(N10797), .ZN(N35843));
    NANDX1 U22972 (.A1(n18914), .A2(n23379), .ZN(N35844));
    NOR2X1 U22973 (.A1(n17085), .A2(N9874), .ZN(N35845));
    INVX1 U22974 (.I(n15789), .ZN(N35846));
    INVX1 U22975 (.I(N5285), .ZN(N35847));
    INVX1 U22976 (.I(N5518), .ZN(N35848));
    NOR2X1 U22977 (.A1(N566), .A2(N3144), .ZN(N35849));
    INVX1 U22978 (.I(n18458), .ZN(n35850));
    INVX1 U22979 (.I(N3167), .ZN(N35851));
    NANDX1 U22980 (.A1(n28142), .A2(n23062), .ZN(N35852));
    NOR2X1 U22981 (.A1(n16257), .A2(n27857), .ZN(N35853));
    NOR2X1 U22982 (.A1(n25613), .A2(n23669), .ZN(n35854));
    NANDX1 U22983 (.A1(N10032), .A2(N4328), .ZN(N35855));
    INVX1 U22984 (.I(n17506), .ZN(N35856));
    NANDX1 U22985 (.A1(n22778), .A2(n23152), .ZN(n35857));
    NANDX1 U22986 (.A1(n20235), .A2(N8803), .ZN(N35858));
    NOR2X1 U22987 (.A1(n14081), .A2(n23311), .ZN(n35859));
    NANDX1 U22988 (.A1(N8862), .A2(N12437), .ZN(N35860));
    NOR2X1 U22989 (.A1(N12017), .A2(n19456), .ZN(N35861));
    NOR2X1 U22990 (.A1(N3744), .A2(n28820), .ZN(N35862));
    NANDX1 U22991 (.A1(n15367), .A2(N8584), .ZN(N35863));
    NANDX1 U22992 (.A1(n13086), .A2(N5506), .ZN(N35864));
    NANDX1 U22993 (.A1(N6617), .A2(N1170), .ZN(N35865));
    INVX1 U22994 (.I(n29642), .ZN(n35866));
    INVX1 U22995 (.I(N9160), .ZN(n35867));
    INVX1 U22996 (.I(n28238), .ZN(N35868));
    NANDX1 U22997 (.A1(N334), .A2(N6896), .ZN(N35869));
    NANDX1 U22998 (.A1(n27661), .A2(n20976), .ZN(N35870));
    NANDX1 U22999 (.A1(N231), .A2(n18399), .ZN(n35871));
    NANDX1 U23000 (.A1(N6082), .A2(n18976), .ZN(N35872));
    NANDX1 U23001 (.A1(N846), .A2(n22719), .ZN(n35873));
    INVX1 U23002 (.I(N12313), .ZN(n35874));
    NANDX1 U23003 (.A1(N8989), .A2(N9900), .ZN(N35875));
    NANDX1 U23004 (.A1(N3055), .A2(n21659), .ZN(N35876));
    INVX1 U23005 (.I(N4224), .ZN(n35877));
    NOR2X1 U23006 (.A1(n15714), .A2(n28382), .ZN(N35878));
    NANDX1 U23007 (.A1(n20045), .A2(n26482), .ZN(n35879));
    INVX1 U23008 (.I(N8940), .ZN(N35880));
    NOR2X1 U23009 (.A1(N1305), .A2(N6463), .ZN(n35881));
    NANDX1 U23010 (.A1(N12712), .A2(N6694), .ZN(n35882));
    NOR2X1 U23011 (.A1(n25117), .A2(N12775), .ZN(n35883));
    NOR2X1 U23012 (.A1(n26840), .A2(N2181), .ZN(N35884));
    NOR2X1 U23013 (.A1(n27245), .A2(n14494), .ZN(N35885));
    NOR2X1 U23014 (.A1(n24794), .A2(n12954), .ZN(n35886));
    INVX1 U23015 (.I(n16410), .ZN(n35887));
    NANDX1 U23016 (.A1(N4769), .A2(N9194), .ZN(n35888));
    NOR2X1 U23017 (.A1(N9043), .A2(N7438), .ZN(N35889));
    NANDX1 U23018 (.A1(n29088), .A2(n22480), .ZN(n35890));
    NANDX1 U23019 (.A1(n26588), .A2(n25720), .ZN(N35891));
    INVX1 U23020 (.I(N2913), .ZN(N35892));
    INVX1 U23021 (.I(N10287), .ZN(N35893));
    NOR2X1 U23022 (.A1(n28094), .A2(n23964), .ZN(N35894));
    NANDX1 U23023 (.A1(N6530), .A2(N9228), .ZN(N35895));
    NOR2X1 U23024 (.A1(N7684), .A2(N6335), .ZN(N35896));
    NANDX1 U23025 (.A1(n16786), .A2(n19690), .ZN(N35897));
    INVX1 U23026 (.I(N5345), .ZN(N35898));
    INVX1 U23027 (.I(N10725), .ZN(N35899));
    INVX1 U23028 (.I(n15155), .ZN(N35900));
    NOR2X1 U23029 (.A1(N7716), .A2(N11154), .ZN(N35901));
    INVX1 U23030 (.I(n25364), .ZN(n35902));
    INVX1 U23031 (.I(n19286), .ZN(N35903));
    NOR2X1 U23032 (.A1(n17776), .A2(n16860), .ZN(n35904));
    NOR2X1 U23033 (.A1(n14695), .A2(n15707), .ZN(N35905));
    NANDX1 U23034 (.A1(N1212), .A2(N9534), .ZN(N35906));
    NANDX1 U23035 (.A1(N7741), .A2(n18761), .ZN(N35907));
    INVX1 U23036 (.I(N3986), .ZN(N35908));
    NANDX1 U23037 (.A1(n17374), .A2(N9332), .ZN(n35909));
    INVX1 U23038 (.I(n23624), .ZN(N35910));
    NOR2X1 U23039 (.A1(n27867), .A2(n22909), .ZN(N35911));
    INVX1 U23040 (.I(n12885), .ZN(n35912));
    NOR2X1 U23041 (.A1(n28324), .A2(N12599), .ZN(N35913));
    NOR2X1 U23042 (.A1(N12111), .A2(n16094), .ZN(N35914));
    NOR2X1 U23043 (.A1(n22486), .A2(N3733), .ZN(n35915));
    NANDX1 U23044 (.A1(n24334), .A2(n18427), .ZN(n35916));
    NANDX1 U23045 (.A1(n24348), .A2(n19639), .ZN(N35917));
    NANDX1 U23046 (.A1(N5166), .A2(n15940), .ZN(N35918));
    NANDX1 U23047 (.A1(N6364), .A2(N8486), .ZN(N35919));
    INVX1 U23048 (.I(N12298), .ZN(n35920));
    NANDX1 U23049 (.A1(N958), .A2(N5784), .ZN(N35921));
    NANDX1 U23050 (.A1(n28825), .A2(n28693), .ZN(n35922));
    NOR2X1 U23051 (.A1(N133), .A2(n15659), .ZN(N35923));
    INVX1 U23052 (.I(N12731), .ZN(N35924));
    INVX1 U23053 (.I(n17641), .ZN(n35925));
    NANDX1 U23054 (.A1(N1890), .A2(n28687), .ZN(N35926));
    INVX1 U23055 (.I(n13698), .ZN(N35927));
    NOR2X1 U23056 (.A1(N9407), .A2(n22514), .ZN(n35928));
    INVX1 U23057 (.I(n17606), .ZN(N35929));
    NOR2X1 U23058 (.A1(N10820), .A2(N3408), .ZN(n35930));
    NANDX1 U23059 (.A1(n17184), .A2(N455), .ZN(N35931));
    NANDX1 U23060 (.A1(n29481), .A2(N6833), .ZN(N35932));
    NANDX1 U23061 (.A1(n23826), .A2(n16447), .ZN(N35933));
    NOR2X1 U23062 (.A1(N10942), .A2(N5093), .ZN(N35934));
    NANDX1 U23063 (.A1(n26600), .A2(n22062), .ZN(N35935));
    NOR2X1 U23064 (.A1(N10662), .A2(n28264), .ZN(N35936));
    NANDX1 U23065 (.A1(N1112), .A2(n26813), .ZN(n35937));
    NOR2X1 U23066 (.A1(n14809), .A2(N8120), .ZN(N35938));
    NANDX1 U23067 (.A1(n25884), .A2(n13774), .ZN(n35939));
    INVX1 U23068 (.I(N6473), .ZN(N35940));
    NOR2X1 U23069 (.A1(n28241), .A2(n19991), .ZN(N35941));
    NOR2X1 U23070 (.A1(n28695), .A2(N12562), .ZN(n35942));
    INVX1 U23071 (.I(n24088), .ZN(N35943));
    NANDX1 U23072 (.A1(N11930), .A2(N10398), .ZN(N35944));
    INVX1 U23073 (.I(n22871), .ZN(n35945));
    NOR2X1 U23074 (.A1(n16609), .A2(n19333), .ZN(n35946));
    INVX1 U23075 (.I(n17506), .ZN(N35947));
    NANDX1 U23076 (.A1(n24239), .A2(n17089), .ZN(N35948));
    NANDX1 U23077 (.A1(N9475), .A2(n26350), .ZN(N35949));
    NOR2X1 U23078 (.A1(n17594), .A2(n14880), .ZN(N35950));
    NANDX1 U23079 (.A1(N1230), .A2(n21015), .ZN(n35951));
    INVX1 U23080 (.I(n25823), .ZN(N35952));
    NOR2X1 U23081 (.A1(n22367), .A2(n14583), .ZN(N35953));
    NANDX1 U23082 (.A1(N4791), .A2(N2687), .ZN(N35954));
    NOR2X1 U23083 (.A1(N10880), .A2(n14616), .ZN(N35955));
    INVX1 U23084 (.I(n16443), .ZN(n35956));
    NOR2X1 U23085 (.A1(n21894), .A2(n21612), .ZN(N35957));
    INVX1 U23086 (.I(n17869), .ZN(N35958));
    NOR2X1 U23087 (.A1(n22358), .A2(N531), .ZN(N35959));
    NOR2X1 U23088 (.A1(N448), .A2(N10006), .ZN(n35960));
    INVX1 U23089 (.I(N12044), .ZN(N35961));
    NOR2X1 U23090 (.A1(n25721), .A2(n19387), .ZN(N35962));
    NOR2X1 U23091 (.A1(N5160), .A2(n21762), .ZN(n35963));
    INVX1 U23092 (.I(N12839), .ZN(n35964));
    NANDX1 U23093 (.A1(n27657), .A2(n26334), .ZN(N35965));
    NOR2X1 U23094 (.A1(n18905), .A2(n15082), .ZN(N35966));
    NOR2X1 U23095 (.A1(N3383), .A2(N2788), .ZN(n35967));
    NOR2X1 U23096 (.A1(n29430), .A2(n24682), .ZN(n35968));
    NOR2X1 U23097 (.A1(n14534), .A2(N974), .ZN(n35969));
    NOR2X1 U23098 (.A1(N6754), .A2(N1505), .ZN(n35970));
    NOR2X1 U23099 (.A1(n25899), .A2(N71), .ZN(N35971));
    INVX1 U23100 (.I(N7806), .ZN(N35972));
    NOR2X1 U23101 (.A1(n14593), .A2(n15753), .ZN(N35973));
    NANDX1 U23102 (.A1(n19752), .A2(n26075), .ZN(N35974));
    NOR2X1 U23103 (.A1(n21151), .A2(n28627), .ZN(N35975));
    NANDX1 U23104 (.A1(n17348), .A2(N5831), .ZN(n35976));
    INVX1 U23105 (.I(n20990), .ZN(N35977));
    NANDX1 U23106 (.A1(n13484), .A2(N12339), .ZN(n35978));
    NANDX1 U23107 (.A1(N12776), .A2(n25581), .ZN(N35979));
    NOR2X1 U23108 (.A1(n15871), .A2(n26554), .ZN(N35980));
    NANDX1 U23109 (.A1(N11185), .A2(n16619), .ZN(N35981));
    NANDX1 U23110 (.A1(N6947), .A2(n16689), .ZN(N35982));
    NANDX1 U23111 (.A1(N3313), .A2(N2782), .ZN(N35983));
    NOR2X1 U23112 (.A1(n19065), .A2(n24961), .ZN(N35984));
    NANDX1 U23113 (.A1(N3563), .A2(n30078), .ZN(n35985));
    INVX1 U23114 (.I(N2052), .ZN(N35986));
    NOR2X1 U23115 (.A1(N11004), .A2(n26581), .ZN(N35987));
    INVX1 U23116 (.I(N1856), .ZN(N35988));
    NANDX1 U23117 (.A1(n14722), .A2(N2755), .ZN(N35989));
    NOR2X1 U23118 (.A1(n27498), .A2(n28335), .ZN(n35990));
    NANDX1 U23119 (.A1(N1792), .A2(n13313), .ZN(n35991));
    INVX1 U23120 (.I(n12976), .ZN(N35992));
    NOR2X1 U23121 (.A1(n20152), .A2(n19922), .ZN(n35993));
    NOR2X1 U23122 (.A1(n22768), .A2(n23234), .ZN(N35994));
    NANDX1 U23123 (.A1(N9839), .A2(N722), .ZN(N35995));
    NANDX1 U23124 (.A1(n23920), .A2(N4285), .ZN(N35996));
    NANDX1 U23125 (.A1(n29015), .A2(n25034), .ZN(n35997));
    INVX1 U23126 (.I(N9881), .ZN(N35998));
    INVX1 U23127 (.I(n13661), .ZN(n35999));
    INVX1 U23128 (.I(n19093), .ZN(N36000));
    NANDX1 U23129 (.A1(N3052), .A2(n18228), .ZN(N36001));
    NOR2X1 U23130 (.A1(N1250), .A2(N3441), .ZN(N36002));
    NANDX1 U23131 (.A1(n14562), .A2(n28547), .ZN(N36003));
    NANDX1 U23132 (.A1(N2916), .A2(N7123), .ZN(N36004));
    INVX1 U23133 (.I(N7959), .ZN(N36005));
    INVX1 U23134 (.I(n19210), .ZN(N36006));
    NANDX1 U23135 (.A1(n16850), .A2(n19932), .ZN(n36007));
    NANDX1 U23136 (.A1(N10632), .A2(N12777), .ZN(N36008));
    NOR2X1 U23137 (.A1(n28208), .A2(N7673), .ZN(n36009));
    NANDX1 U23138 (.A1(N7951), .A2(n29150), .ZN(n36010));
    NANDX1 U23139 (.A1(N8248), .A2(N6666), .ZN(N36011));
    NOR2X1 U23140 (.A1(n29998), .A2(n13454), .ZN(n36012));
    NOR2X1 U23141 (.A1(N1110), .A2(n16895), .ZN(N36013));
    INVX1 U23142 (.I(n15671), .ZN(n36014));
    NANDX1 U23143 (.A1(N1862), .A2(N7147), .ZN(n36015));
    INVX1 U23144 (.I(n27975), .ZN(N36016));
    INVX1 U23145 (.I(n17998), .ZN(N36017));
    INVX1 U23146 (.I(N8010), .ZN(n36018));
    NANDX1 U23147 (.A1(n25539), .A2(n22260), .ZN(N36019));
    INVX1 U23148 (.I(N8178), .ZN(N36020));
    INVX1 U23149 (.I(N1973), .ZN(n36021));
    INVX1 U23150 (.I(n22602), .ZN(N36022));
    NANDX1 U23151 (.A1(N3424), .A2(N12507), .ZN(n36023));
    NANDX1 U23152 (.A1(n28787), .A2(N7917), .ZN(N36024));
    NOR2X1 U23153 (.A1(N12104), .A2(N6190), .ZN(N36025));
    NOR2X1 U23154 (.A1(n28998), .A2(N9119), .ZN(N36026));
    INVX1 U23155 (.I(n21423), .ZN(N36027));
    INVX1 U23156 (.I(N7639), .ZN(n36028));
    INVX1 U23157 (.I(n27515), .ZN(N36029));
    NOR2X1 U23158 (.A1(N8831), .A2(N2985), .ZN(N36030));
    INVX1 U23159 (.I(n13541), .ZN(N36031));
    NANDX1 U23160 (.A1(N11437), .A2(N6004), .ZN(n36032));
    INVX1 U23161 (.I(n27656), .ZN(n36033));
    NANDX1 U23162 (.A1(N10975), .A2(n20120), .ZN(n36034));
    NOR2X1 U23163 (.A1(n14398), .A2(N2490), .ZN(N36035));
    NANDX1 U23164 (.A1(N1609), .A2(n29104), .ZN(N36036));
    NANDX1 U23165 (.A1(n13712), .A2(N5156), .ZN(N36037));
    INVX1 U23166 (.I(N1133), .ZN(N36038));
    NOR2X1 U23167 (.A1(N12354), .A2(n22555), .ZN(n36039));
    NOR2X1 U23168 (.A1(n19993), .A2(n13388), .ZN(n36040));
    NOR2X1 U23169 (.A1(N1160), .A2(n22219), .ZN(N36041));
    NANDX1 U23170 (.A1(n20474), .A2(n24320), .ZN(N36042));
    INVX1 U23171 (.I(N1774), .ZN(N36043));
    NOR2X1 U23172 (.A1(n14945), .A2(n17990), .ZN(N36044));
    INVX1 U23173 (.I(n25920), .ZN(n36045));
    NOR2X1 U23174 (.A1(n21878), .A2(n28878), .ZN(n36046));
    NANDX1 U23175 (.A1(n23629), .A2(N349), .ZN(N36047));
    NANDX1 U23176 (.A1(n20531), .A2(N2621), .ZN(N36048));
    INVX1 U23177 (.I(N2256), .ZN(n36049));
    NOR2X1 U23178 (.A1(n24677), .A2(N3170), .ZN(N36050));
    INVX1 U23179 (.I(n15612), .ZN(N36051));
    NOR2X1 U23180 (.A1(n28256), .A2(n15364), .ZN(N36052));
    NOR2X1 U23181 (.A1(N8898), .A2(N6661), .ZN(N36053));
    INVX1 U23182 (.I(n21778), .ZN(n36054));
    INVX1 U23183 (.I(n23690), .ZN(N36055));
    NANDX1 U23184 (.A1(n29986), .A2(N11543), .ZN(n36056));
    NANDX1 U23185 (.A1(n14329), .A2(N8076), .ZN(N36057));
    INVX1 U23186 (.I(n13070), .ZN(N36058));
    INVX1 U23187 (.I(N11175), .ZN(N36059));
    NOR2X1 U23188 (.A1(n23784), .A2(n20266), .ZN(N36060));
    NANDX1 U23189 (.A1(N4049), .A2(N11082), .ZN(N36061));
    INVX1 U23190 (.I(n17286), .ZN(n36062));
    NOR2X1 U23191 (.A1(n23220), .A2(N2761), .ZN(N36063));
    NOR2X1 U23192 (.A1(n21339), .A2(N6685), .ZN(n36064));
    NANDX1 U23193 (.A1(n18797), .A2(N1906), .ZN(N36065));
    INVX1 U23194 (.I(N10438), .ZN(N36066));
    INVX1 U23195 (.I(N12749), .ZN(n36067));
    INVX1 U23196 (.I(n16795), .ZN(N36068));
    NANDX1 U23197 (.A1(N5328), .A2(N987), .ZN(N36069));
    INVX1 U23198 (.I(n23011), .ZN(N36070));
    INVX1 U23199 (.I(n28024), .ZN(n36071));
    NOR2X1 U23200 (.A1(N4595), .A2(N10231), .ZN(N36072));
    INVX1 U23201 (.I(N9194), .ZN(N36073));
    NANDX1 U23202 (.A1(n23956), .A2(N6107), .ZN(N36074));
    NOR2X1 U23203 (.A1(n26768), .A2(n29326), .ZN(n36075));
    NANDX1 U23204 (.A1(n22604), .A2(N9088), .ZN(N36076));
    NANDX1 U23205 (.A1(N1186), .A2(n16446), .ZN(N36077));
    NANDX1 U23206 (.A1(n20382), .A2(n26883), .ZN(n36078));
    NOR2X1 U23207 (.A1(N2993), .A2(n24965), .ZN(n36079));
    NOR2X1 U23208 (.A1(n15845), .A2(N155), .ZN(N36080));
    INVX1 U23209 (.I(n25332), .ZN(N36081));
    INVX1 U23210 (.I(n15803), .ZN(n36082));
    INVX1 U23211 (.I(n15773), .ZN(N36083));
    INVX1 U23212 (.I(n22010), .ZN(n36084));
    NANDX1 U23213 (.A1(n18152), .A2(N6152), .ZN(n36085));
    INVX1 U23214 (.I(n24258), .ZN(N36086));
    NANDX1 U23215 (.A1(N7656), .A2(N12007), .ZN(N36087));
    INVX1 U23216 (.I(N122), .ZN(n36088));
    NOR2X1 U23217 (.A1(n29898), .A2(n20005), .ZN(N36089));
    INVX1 U23218 (.I(N1098), .ZN(n36090));
    NANDX1 U23219 (.A1(N11407), .A2(n19382), .ZN(N36091));
    NANDX1 U23220 (.A1(N6234), .A2(n12884), .ZN(N36092));
    NOR2X1 U23221 (.A1(N6389), .A2(n26070), .ZN(N36093));
    INVX1 U23222 (.I(n18114), .ZN(N36094));
    NANDX1 U23223 (.A1(n13181), .A2(N3750), .ZN(n36095));
    NANDX1 U23224 (.A1(N5054), .A2(n20957), .ZN(n36096));
    NANDX1 U23225 (.A1(n29903), .A2(n20543), .ZN(N36097));
    NOR2X1 U23226 (.A1(n26043), .A2(n28198), .ZN(N36098));
    INVX1 U23227 (.I(n26371), .ZN(n36099));
    INVX1 U23228 (.I(N1610), .ZN(N36100));
    NANDX1 U23229 (.A1(n25446), .A2(n27710), .ZN(n36101));
    INVX1 U23230 (.I(n24255), .ZN(N36102));
    NOR2X1 U23231 (.A1(n23731), .A2(n26057), .ZN(N36103));
    NOR2X1 U23232 (.A1(n25175), .A2(N2127), .ZN(n36104));
    NANDX1 U23233 (.A1(N9668), .A2(N3529), .ZN(N36105));
    NANDX1 U23234 (.A1(N9963), .A2(N5270), .ZN(N36106));
    NANDX1 U23235 (.A1(n19216), .A2(n29021), .ZN(N36107));
    NANDX1 U23236 (.A1(n16482), .A2(n28787), .ZN(N36108));
    NANDX1 U23237 (.A1(n26567), .A2(n24692), .ZN(N36109));
    INVX1 U23238 (.I(n18521), .ZN(n36110));
    NANDX1 U23239 (.A1(N5309), .A2(n20130), .ZN(N36111));
    NOR2X1 U23240 (.A1(n19315), .A2(N6263), .ZN(N36112));
    NANDX1 U23241 (.A1(n13433), .A2(n15241), .ZN(N36113));
    NANDX1 U23242 (.A1(N9352), .A2(n19013), .ZN(N36114));
    NOR2X1 U23243 (.A1(N11479), .A2(n29174), .ZN(N36115));
    NANDX1 U23244 (.A1(N3568), .A2(n15872), .ZN(N36116));
    NOR2X1 U23245 (.A1(N8837), .A2(N6319), .ZN(N36117));
    NOR2X1 U23246 (.A1(N7721), .A2(n17722), .ZN(N36118));
    INVX1 U23247 (.I(n25068), .ZN(n36119));
    NOR2X1 U23248 (.A1(n27337), .A2(N8183), .ZN(n36120));
    INVX1 U23249 (.I(N4281), .ZN(N36121));
    INVX1 U23250 (.I(N1828), .ZN(N36122));
    INVX1 U23251 (.I(N269), .ZN(N36123));
    NOR2X1 U23252 (.A1(n19233), .A2(n17356), .ZN(N36124));
    INVX1 U23253 (.I(n23034), .ZN(N36125));
    NOR2X1 U23254 (.A1(N2350), .A2(N11910), .ZN(n36126));
    NANDX1 U23255 (.A1(N2389), .A2(n29644), .ZN(N36127));
    NOR2X1 U23256 (.A1(N5956), .A2(n15378), .ZN(n36128));
    NANDX1 U23257 (.A1(N3354), .A2(n21696), .ZN(n36129));
    NANDX1 U23258 (.A1(n29772), .A2(n27978), .ZN(N36130));
    NOR2X1 U23259 (.A1(n24702), .A2(N5931), .ZN(N36131));
    NOR2X1 U23260 (.A1(N2747), .A2(N2450), .ZN(n36132));
    NOR2X1 U23261 (.A1(N8976), .A2(n22975), .ZN(N36133));
    INVX1 U23262 (.I(n27943), .ZN(N36134));
    NANDX1 U23263 (.A1(n28777), .A2(n15161), .ZN(N36135));
    NOR2X1 U23264 (.A1(n21673), .A2(N1621), .ZN(n36136));
    INVX1 U23265 (.I(N3445), .ZN(n36137));
    NOR2X1 U23266 (.A1(N277), .A2(n21649), .ZN(N36138));
    NOR2X1 U23267 (.A1(n24931), .A2(N6889), .ZN(N36139));
    NANDX1 U23268 (.A1(n16845), .A2(n17145), .ZN(N36140));
    INVX1 U23269 (.I(n16479), .ZN(N36141));
    NANDX1 U23270 (.A1(n20611), .A2(n29741), .ZN(n36142));
    INVX1 U23271 (.I(n12903), .ZN(N36143));
    INVX1 U23272 (.I(N11925), .ZN(n36144));
    INVX1 U23273 (.I(n30024), .ZN(N36145));
    NANDX1 U23274 (.A1(n19020), .A2(n16390), .ZN(N36146));
    INVX1 U23275 (.I(n17659), .ZN(n36147));
    NOR2X1 U23276 (.A1(N2842), .A2(N9194), .ZN(N36148));
    NOR2X1 U23277 (.A1(N730), .A2(N1200), .ZN(n36149));
    NANDX1 U23278 (.A1(n19704), .A2(n22848), .ZN(N36150));
    NANDX1 U23279 (.A1(n14497), .A2(n18298), .ZN(N36151));
    NANDX1 U23280 (.A1(N1204), .A2(N5305), .ZN(n36152));
    NOR2X1 U23281 (.A1(N6243), .A2(N8851), .ZN(N36153));
    INVX1 U23282 (.I(N5846), .ZN(N36154));
    NOR2X1 U23283 (.A1(n19784), .A2(n26894), .ZN(N36155));
    NOR2X1 U23284 (.A1(n17821), .A2(n15341), .ZN(n36156));
    NANDX1 U23285 (.A1(N6703), .A2(N1593), .ZN(n36157));
    NANDX1 U23286 (.A1(n12922), .A2(n21703), .ZN(N36158));
    INVX1 U23287 (.I(n22115), .ZN(N36159));
    NOR2X1 U23288 (.A1(N129), .A2(n23314), .ZN(N36160));
    NANDX1 U23289 (.A1(n19833), .A2(N4586), .ZN(N36161));
    INVX1 U23290 (.I(N4192), .ZN(n36162));
    INVX1 U23291 (.I(N3393), .ZN(N36163));
    NOR2X1 U23292 (.A1(n16748), .A2(N1103), .ZN(N36164));
    NANDX1 U23293 (.A1(n25598), .A2(N7984), .ZN(n36165));
    NANDX1 U23294 (.A1(N2348), .A2(n16329), .ZN(n36166));
    NANDX1 U23295 (.A1(N9720), .A2(N4012), .ZN(n36167));
    NANDX1 U23296 (.A1(n21854), .A2(N10714), .ZN(n36168));
    NANDX1 U23297 (.A1(n29851), .A2(n23635), .ZN(N36169));
    NANDX1 U23298 (.A1(N10553), .A2(N4173), .ZN(N36170));
    NOR2X1 U23299 (.A1(N10681), .A2(n16048), .ZN(n36171));
    INVX1 U23300 (.I(n19074), .ZN(N36172));
    NANDX1 U23301 (.A1(N8727), .A2(n23266), .ZN(n36173));
    NOR2X1 U23302 (.A1(N12120), .A2(n17222), .ZN(N36174));
    NOR2X1 U23303 (.A1(n13222), .A2(N5981), .ZN(N36175));
    INVX1 U23304 (.I(N9767), .ZN(N36176));
    NANDX1 U23305 (.A1(n23753), .A2(n26095), .ZN(N36177));
    INVX1 U23306 (.I(N3335), .ZN(N36178));
    NOR2X1 U23307 (.A1(N10087), .A2(n13749), .ZN(n36179));
    NOR2X1 U23308 (.A1(n18380), .A2(N2023), .ZN(N36180));
    INVX1 U23309 (.I(N6800), .ZN(N36181));
    NOR2X1 U23310 (.A1(n15610), .A2(N8516), .ZN(N36182));
    NANDX1 U23311 (.A1(N1520), .A2(N8921), .ZN(n36183));
    NOR2X1 U23312 (.A1(N10713), .A2(n17647), .ZN(n36184));
    NOR2X1 U23313 (.A1(N12651), .A2(n18327), .ZN(n36185));
    NANDX1 U23314 (.A1(N1200), .A2(N1412), .ZN(N36186));
    NOR2X1 U23315 (.A1(n22605), .A2(N11178), .ZN(N36187));
    INVX1 U23316 (.I(n16220), .ZN(N36188));
    INVX1 U23317 (.I(n28313), .ZN(N36189));
    NOR2X1 U23318 (.A1(n25801), .A2(N8262), .ZN(n36190));
    INVX1 U23319 (.I(n25043), .ZN(N36191));
    NANDX1 U23320 (.A1(N12446), .A2(N6343), .ZN(N36192));
    NANDX1 U23321 (.A1(n13582), .A2(n21952), .ZN(N36193));
    INVX1 U23322 (.I(n25398), .ZN(N36194));
    INVX1 U23323 (.I(n16559), .ZN(N36195));
    INVX1 U23324 (.I(n22745), .ZN(N36196));
    INVX1 U23325 (.I(n15851), .ZN(N36197));
    NOR2X1 U23326 (.A1(N10956), .A2(N4074), .ZN(N36198));
    NANDX1 U23327 (.A1(N928), .A2(n16976), .ZN(n36199));
    INVX1 U23328 (.I(N666), .ZN(n36200));
    NANDX1 U23329 (.A1(n22403), .A2(n26498), .ZN(N36201));
    INVX1 U23330 (.I(n19078), .ZN(N36202));
    INVX1 U23331 (.I(N6763), .ZN(n36203));
    NANDX1 U23332 (.A1(N5627), .A2(n21965), .ZN(n36204));
    NOR2X1 U23333 (.A1(N11969), .A2(n21088), .ZN(N36205));
    NANDX1 U23334 (.A1(n22481), .A2(n28726), .ZN(N36206));
    NOR2X1 U23335 (.A1(N4376), .A2(N3708), .ZN(n36207));
    NANDX1 U23336 (.A1(n27121), .A2(n26474), .ZN(n36208));
    NOR2X1 U23337 (.A1(N2242), .A2(n25990), .ZN(N36209));
    NOR2X1 U23338 (.A1(n15958), .A2(n26917), .ZN(N36210));
    NOR2X1 U23339 (.A1(n22141), .A2(n16143), .ZN(n36211));
    INVX1 U23340 (.I(n14406), .ZN(N36212));
    NANDX1 U23341 (.A1(n29511), .A2(N3346), .ZN(n36213));
    NOR2X1 U23342 (.A1(N6136), .A2(N2709), .ZN(N36214));
    NOR2X1 U23343 (.A1(n16662), .A2(N3078), .ZN(N36215));
    INVX1 U23344 (.I(N7612), .ZN(N36216));
    NANDX1 U23345 (.A1(N10283), .A2(N6201), .ZN(n36217));
    NANDX1 U23346 (.A1(n14659), .A2(n28606), .ZN(n36218));
    NOR2X1 U23347 (.A1(N11642), .A2(n24942), .ZN(N36219));
    NOR2X1 U23348 (.A1(N2444), .A2(n20794), .ZN(n36220));
    NOR2X1 U23349 (.A1(n18401), .A2(N6134), .ZN(n36221));
    NOR2X1 U23350 (.A1(N10404), .A2(n22276), .ZN(N36222));
    NOR2X1 U23351 (.A1(n13370), .A2(n23339), .ZN(n36223));
    INVX1 U23352 (.I(n16715), .ZN(N36224));
    NOR2X1 U23353 (.A1(n14873), .A2(N7984), .ZN(N36225));
    NANDX1 U23354 (.A1(n20095), .A2(N11061), .ZN(N36226));
    NOR2X1 U23355 (.A1(n16268), .A2(n28089), .ZN(N36227));
    NOR2X1 U23356 (.A1(N11029), .A2(n24191), .ZN(N36228));
    NANDX1 U23357 (.A1(N9497), .A2(n21335), .ZN(N36229));
    NANDX1 U23358 (.A1(N4302), .A2(n16675), .ZN(N36230));
    INVX1 U23359 (.I(n13656), .ZN(N36231));
    NANDX1 U23360 (.A1(N7349), .A2(N8351), .ZN(N36232));
    INVX1 U23361 (.I(N6313), .ZN(N36233));
    NANDX1 U23362 (.A1(n24880), .A2(n19682), .ZN(N36234));
    NOR2X1 U23363 (.A1(N3480), .A2(n24957), .ZN(N36235));
    NOR2X1 U23364 (.A1(n18352), .A2(N2803), .ZN(N36236));
    NANDX1 U23365 (.A1(n27008), .A2(N2424), .ZN(n36237));
    NANDX1 U23366 (.A1(n13138), .A2(N376), .ZN(N36238));
    INVX1 U23367 (.I(n24166), .ZN(N36239));
    INVX1 U23368 (.I(n19354), .ZN(n36240));
    NOR2X1 U23369 (.A1(n23022), .A2(N5859), .ZN(N36241));
    NOR2X1 U23370 (.A1(N9559), .A2(n24944), .ZN(N36242));
    NANDX1 U23371 (.A1(n19661), .A2(n20853), .ZN(n36243));
    NANDX1 U23372 (.A1(N12298), .A2(n15726), .ZN(n36244));
    INVX1 U23373 (.I(n25738), .ZN(n36245));
    NOR2X1 U23374 (.A1(N1132), .A2(n29217), .ZN(N36246));
    NANDX1 U23375 (.A1(n29945), .A2(N5993), .ZN(N36247));
    NOR2X1 U23376 (.A1(n20879), .A2(N2863), .ZN(n36248));
    NOR2X1 U23377 (.A1(N3312), .A2(N4561), .ZN(N36249));
    INVX1 U23378 (.I(N6226), .ZN(N36250));
    NOR2X1 U23379 (.A1(n14636), .A2(n25579), .ZN(N36251));
    NANDX1 U23380 (.A1(N7520), .A2(n19999), .ZN(N36252));
    NOR2X1 U23381 (.A1(N5640), .A2(N3366), .ZN(n36253));
    NANDX1 U23382 (.A1(n13861), .A2(n24219), .ZN(n36254));
    NOR2X1 U23383 (.A1(n26159), .A2(N9807), .ZN(n36255));
    NOR2X1 U23384 (.A1(N10320), .A2(N3638), .ZN(N36256));
    INVX1 U23385 (.I(n28098), .ZN(N36257));
    NANDX1 U23386 (.A1(N12436), .A2(N3953), .ZN(n36258));
    NOR2X1 U23387 (.A1(n21875), .A2(n25513), .ZN(N36259));
    NANDX1 U23388 (.A1(n13747), .A2(n30073), .ZN(N36260));
    NOR2X1 U23389 (.A1(n19972), .A2(n17222), .ZN(N36261));
    INVX1 U23390 (.I(N3975), .ZN(N36262));
    NANDX1 U23391 (.A1(N8536), .A2(N12534), .ZN(N36263));
    NANDX1 U23392 (.A1(N2736), .A2(n15899), .ZN(N36264));
    NOR2X1 U23393 (.A1(n16597), .A2(N9980), .ZN(N36265));
    NANDX1 U23394 (.A1(N1179), .A2(N8348), .ZN(N36266));
    NOR2X1 U23395 (.A1(N11498), .A2(N546), .ZN(N36267));
    NOR2X1 U23396 (.A1(N9458), .A2(N11530), .ZN(n36268));
    NOR2X1 U23397 (.A1(N1971), .A2(n13966), .ZN(n36269));
    NANDX1 U23398 (.A1(n16044), .A2(n28975), .ZN(n36270));
    NOR2X1 U23399 (.A1(n15979), .A2(n15356), .ZN(N36271));
    INVX1 U23400 (.I(N3063), .ZN(N36272));
    NOR2X1 U23401 (.A1(N9086), .A2(N10958), .ZN(N36273));
    NANDX1 U23402 (.A1(n21619), .A2(n17351), .ZN(N36274));
    NANDX1 U23403 (.A1(N7380), .A2(N9408), .ZN(N36275));
    NOR2X1 U23404 (.A1(N5921), .A2(n28397), .ZN(N36276));
    INVX1 U23405 (.I(N2829), .ZN(N36277));
    NANDX1 U23406 (.A1(N11159), .A2(N3374), .ZN(N36278));
    INVX1 U23407 (.I(N9177), .ZN(N36279));
    INVX1 U23408 (.I(N2681), .ZN(n36280));
    INVX1 U23409 (.I(n17430), .ZN(N36281));
    NANDX1 U23410 (.A1(n27191), .A2(n16267), .ZN(N36282));
    NANDX1 U23411 (.A1(N1594), .A2(n20184), .ZN(n36283));
    NANDX1 U23412 (.A1(n23354), .A2(n25116), .ZN(N36284));
    INVX1 U23413 (.I(n22872), .ZN(N36285));
    INVX1 U23414 (.I(N10647), .ZN(N36286));
    INVX1 U23415 (.I(n20471), .ZN(n36287));
    NOR2X1 U23416 (.A1(N8054), .A2(n18953), .ZN(N36288));
    NOR2X1 U23417 (.A1(n25011), .A2(n30053), .ZN(N36289));
    NANDX1 U23418 (.A1(N12181), .A2(n29772), .ZN(n36290));
    NOR2X1 U23419 (.A1(N12327), .A2(N8811), .ZN(n36291));
    NANDX1 U23420 (.A1(n15008), .A2(n19958), .ZN(n36292));
    NANDX1 U23421 (.A1(N520), .A2(N5573), .ZN(N36293));
    NANDX1 U23422 (.A1(N5489), .A2(n25864), .ZN(N36294));
    INVX1 U23423 (.I(n15569), .ZN(N36295));
    NOR2X1 U23424 (.A1(n18014), .A2(N4597), .ZN(N36296));
    INVX1 U23425 (.I(N3582), .ZN(n36297));
    INVX1 U23426 (.I(n29159), .ZN(N36298));
    INVX1 U23427 (.I(N3132), .ZN(n36299));
    INVX1 U23428 (.I(N1429), .ZN(N36300));
    INVX1 U23429 (.I(N1948), .ZN(N36301));
    NANDX1 U23430 (.A1(N836), .A2(n14128), .ZN(n36302));
    NOR2X1 U23431 (.A1(N8104), .A2(n15016), .ZN(n36303));
    NOR2X1 U23432 (.A1(N138), .A2(n18584), .ZN(N36304));
    NANDX1 U23433 (.A1(n28299), .A2(n19103), .ZN(n36305));
    NANDX1 U23434 (.A1(N12453), .A2(n13153), .ZN(n36306));
    NANDX1 U23435 (.A1(N5350), .A2(n28721), .ZN(N36307));
    NANDX1 U23436 (.A1(n23363), .A2(n21879), .ZN(N36308));
    NANDX1 U23437 (.A1(n15506), .A2(N6984), .ZN(N36309));
    NANDX1 U23438 (.A1(n16679), .A2(n28813), .ZN(n36310));
    NOR2X1 U23439 (.A1(n18107), .A2(N2875), .ZN(n36311));
    NOR2X1 U23440 (.A1(n26709), .A2(N3710), .ZN(n36312));
    INVX1 U23441 (.I(N4808), .ZN(N36313));
    INVX1 U23442 (.I(N7610), .ZN(n36314));
    NANDX1 U23443 (.A1(n19210), .A2(n14754), .ZN(N36315));
    NOR2X1 U23444 (.A1(n17371), .A2(N3720), .ZN(n36316));
    NANDX1 U23445 (.A1(n18384), .A2(n16872), .ZN(N36317));
    NOR2X1 U23446 (.A1(n23734), .A2(N4016), .ZN(N36318));
    INVX1 U23447 (.I(N5520), .ZN(N36319));
    NANDX1 U23448 (.A1(n15757), .A2(n21025), .ZN(n36320));
    NANDX1 U23449 (.A1(n26778), .A2(N7567), .ZN(n36321));
    INVX1 U23450 (.I(n14737), .ZN(N36322));
    NANDX1 U23451 (.A1(n22988), .A2(N4643), .ZN(n36323));
    NANDX1 U23452 (.A1(n15258), .A2(n27374), .ZN(n36324));
    NOR2X1 U23453 (.A1(n15632), .A2(n23545), .ZN(N36325));
    INVX1 U23454 (.I(n23402), .ZN(N36326));
    NANDX1 U23455 (.A1(N8993), .A2(N10635), .ZN(n36327));
    NOR2X1 U23456 (.A1(n23095), .A2(n17580), .ZN(N36328));
    NOR2X1 U23457 (.A1(N3786), .A2(N11176), .ZN(N36329));
    NANDX1 U23458 (.A1(n26240), .A2(N5256), .ZN(N36330));
    NOR2X1 U23459 (.A1(N420), .A2(n26281), .ZN(N36331));
    NANDX1 U23460 (.A1(n27197), .A2(n22408), .ZN(n36332));
    NOR2X1 U23461 (.A1(N11796), .A2(n25202), .ZN(N36333));
    NANDX1 U23462 (.A1(N4999), .A2(n24568), .ZN(n36334));
    NANDX1 U23463 (.A1(n20934), .A2(N5864), .ZN(n36335));
    NOR2X1 U23464 (.A1(n14341), .A2(N9013), .ZN(N36336));
    NOR2X1 U23465 (.A1(N11062), .A2(N6567), .ZN(N36337));
    NANDX1 U23466 (.A1(N64), .A2(n18222), .ZN(N36338));
    NANDX1 U23467 (.A1(N5936), .A2(N10569), .ZN(N36339));
    NOR2X1 U23468 (.A1(N4385), .A2(n25369), .ZN(n36340));
    NANDX1 U23469 (.A1(n17289), .A2(n25788), .ZN(N36341));
    NOR2X1 U23470 (.A1(n21493), .A2(n22847), .ZN(N36342));
    NANDX1 U23471 (.A1(N4235), .A2(N4506), .ZN(n36343));
    INVX1 U23472 (.I(N9965), .ZN(N36344));
    NANDX1 U23473 (.A1(n13938), .A2(N815), .ZN(N36345));
    NANDX1 U23474 (.A1(n19801), .A2(n14555), .ZN(N36346));
    NOR2X1 U23475 (.A1(n17374), .A2(N2861), .ZN(N36347));
    NOR2X1 U23476 (.A1(N12501), .A2(N9060), .ZN(N36348));
    NOR2X1 U23477 (.A1(N586), .A2(n14141), .ZN(n36349));
    NOR2X1 U23478 (.A1(N11154), .A2(N7518), .ZN(n36350));
    NANDX1 U23479 (.A1(N6385), .A2(N6151), .ZN(N36351));
    INVX1 U23480 (.I(N2035), .ZN(n36352));
    INVX1 U23481 (.I(n17670), .ZN(N36353));
    NANDX1 U23482 (.A1(N6671), .A2(N10466), .ZN(N36354));
    NOR2X1 U23483 (.A1(N7480), .A2(n20430), .ZN(N36355));
    NANDX1 U23484 (.A1(N9978), .A2(N9805), .ZN(N36356));
    NOR2X1 U23485 (.A1(n29778), .A2(n24359), .ZN(n36357));
    NOR2X1 U23486 (.A1(n17014), .A2(n15780), .ZN(N36358));
    NOR2X1 U23487 (.A1(n29515), .A2(n24839), .ZN(n36359));
    NOR2X1 U23488 (.A1(n18661), .A2(n27540), .ZN(n36360));
    NOR2X1 U23489 (.A1(n29814), .A2(N4921), .ZN(n36361));
    INVX1 U23490 (.I(n24759), .ZN(N36362));
    INVX1 U23491 (.I(N748), .ZN(N36363));
    NOR2X1 U23492 (.A1(N559), .A2(N6979), .ZN(N36364));
    INVX1 U23493 (.I(N7229), .ZN(N36365));
    NANDX1 U23494 (.A1(n16605), .A2(N3269), .ZN(N36366));
    INVX1 U23495 (.I(N9738), .ZN(N36367));
    NANDX1 U23496 (.A1(N6101), .A2(N3170), .ZN(N36368));
    NOR2X1 U23497 (.A1(n19020), .A2(N7062), .ZN(n36369));
    INVX1 U23498 (.I(N4662), .ZN(n36370));
    NANDX1 U23499 (.A1(n25097), .A2(n29500), .ZN(N36371));
    NANDX1 U23500 (.A1(n13620), .A2(n15464), .ZN(N36372));
    NANDX1 U23501 (.A1(N1857), .A2(n20384), .ZN(N36373));
    NANDX1 U23502 (.A1(n26615), .A2(n20015), .ZN(N36374));
    INVX1 U23503 (.I(n23270), .ZN(n36375));
    INVX1 U23504 (.I(n22859), .ZN(N36376));
    INVX1 U23505 (.I(n16363), .ZN(n36377));
    NANDX1 U23506 (.A1(n27092), .A2(N8192), .ZN(N36378));
    NANDX1 U23507 (.A1(N6692), .A2(N9999), .ZN(n36379));
    INVX1 U23508 (.I(n28560), .ZN(N36380));
    NOR2X1 U23509 (.A1(N8702), .A2(n24182), .ZN(N36381));
    NOR2X1 U23510 (.A1(N1924), .A2(n26520), .ZN(n36382));
    NOR2X1 U23511 (.A1(n19984), .A2(n15580), .ZN(N36383));
    NOR2X1 U23512 (.A1(N5310), .A2(N7444), .ZN(n36384));
    NOR2X1 U23513 (.A1(n14254), .A2(n15318), .ZN(N36385));
    NOR2X1 U23514 (.A1(n22830), .A2(N1061), .ZN(n36386));
    NOR2X1 U23515 (.A1(n13265), .A2(n23919), .ZN(N36387));
    NANDX1 U23516 (.A1(n18188), .A2(n22644), .ZN(N36388));
    NOR2X1 U23517 (.A1(n14941), .A2(N6226), .ZN(n36389));
    NANDX1 U23518 (.A1(n13500), .A2(n26045), .ZN(N36390));
    NOR2X1 U23519 (.A1(n24944), .A2(n23307), .ZN(N36391));
    NANDX1 U23520 (.A1(N1834), .A2(n13791), .ZN(n36392));
    INVX1 U23521 (.I(N3819), .ZN(N36393));
    NANDX1 U23522 (.A1(n28711), .A2(N7985), .ZN(N36394));
    INVX1 U23523 (.I(N6017), .ZN(N36395));
    NANDX1 U23524 (.A1(N11761), .A2(N9895), .ZN(N36396));
    NOR2X1 U23525 (.A1(N4453), .A2(N10955), .ZN(n36397));
    NANDX1 U23526 (.A1(N6279), .A2(n23434), .ZN(N36398));
    NOR2X1 U23527 (.A1(n13027), .A2(n15940), .ZN(n36399));
    INVX1 U23528 (.I(n16528), .ZN(N36400));
    INVX1 U23529 (.I(N8212), .ZN(N36401));
    INVX1 U23530 (.I(N6633), .ZN(n36402));
    NOR2X1 U23531 (.A1(n13395), .A2(n29939), .ZN(N36403));
    NANDX1 U23532 (.A1(N3789), .A2(n13592), .ZN(N36404));
    NOR2X1 U23533 (.A1(n26305), .A2(N5790), .ZN(n36405));
    NANDX1 U23534 (.A1(N4152), .A2(N3297), .ZN(N36406));
    NANDX1 U23535 (.A1(n18158), .A2(N3618), .ZN(n36407));
    NOR2X1 U23536 (.A1(n15964), .A2(n26769), .ZN(N36408));
    NANDX1 U23537 (.A1(n28098), .A2(n21608), .ZN(n36409));
    NANDX1 U23538 (.A1(n16214), .A2(N4497), .ZN(N36410));
    NOR2X1 U23539 (.A1(N7402), .A2(n21025), .ZN(n36411));
    NANDX1 U23540 (.A1(N4174), .A2(N9475), .ZN(N36412));
    NOR2X1 U23541 (.A1(n16391), .A2(n22869), .ZN(N36413));
    NOR2X1 U23542 (.A1(n26658), .A2(n26657), .ZN(n36414));
    INVX1 U23543 (.I(n19919), .ZN(N36415));
    NOR2X1 U23544 (.A1(N7281), .A2(N314), .ZN(N36416));
    INVX1 U23545 (.I(n29275), .ZN(n36417));
    NANDX1 U23546 (.A1(n14996), .A2(n21454), .ZN(n36418));
    NANDX1 U23547 (.A1(n19520), .A2(n18085), .ZN(N36419));
    NOR2X1 U23548 (.A1(n17481), .A2(N9555), .ZN(N36420));
    NANDX1 U23549 (.A1(N3557), .A2(N2612), .ZN(N36421));
    NANDX1 U23550 (.A1(n29656), .A2(N12197), .ZN(N36422));
    INVX1 U23551 (.I(n22390), .ZN(N36423));
    NANDX1 U23552 (.A1(N2867), .A2(N8643), .ZN(N36424));
    INVX1 U23553 (.I(n20904), .ZN(N36425));
    NANDX1 U23554 (.A1(n29621), .A2(n22396), .ZN(N36426));
    INVX1 U23555 (.I(n22308), .ZN(N36427));
    NANDX1 U23556 (.A1(N2517), .A2(N7707), .ZN(N36428));
    NANDX1 U23557 (.A1(n19379), .A2(N11264), .ZN(N36429));
    INVX1 U23558 (.I(n21108), .ZN(N36430));
    INVX1 U23559 (.I(n15336), .ZN(N36431));
    NOR2X1 U23560 (.A1(N6687), .A2(n13451), .ZN(N36432));
    INVX1 U23561 (.I(N10243), .ZN(N36433));
    NANDX1 U23562 (.A1(N132), .A2(n28459), .ZN(N36434));
    INVX1 U23563 (.I(n22159), .ZN(N36435));
    NANDX1 U23564 (.A1(N8354), .A2(n13587), .ZN(N36436));
    NOR2X1 U23565 (.A1(n22756), .A2(n23051), .ZN(N36437));
    NANDX1 U23566 (.A1(n22239), .A2(N3870), .ZN(n36438));
    NOR2X1 U23567 (.A1(N2970), .A2(n22107), .ZN(N36439));
    NANDX1 U23568 (.A1(N10677), .A2(n28042), .ZN(n36440));
    INVX1 U23569 (.I(n21940), .ZN(n36441));
    NOR2X1 U23570 (.A1(n22526), .A2(N11146), .ZN(N36442));
    NANDX1 U23571 (.A1(n29745), .A2(n17833), .ZN(N36443));
    NANDX1 U23572 (.A1(N755), .A2(n16636), .ZN(n36444));
    NOR2X1 U23573 (.A1(n19584), .A2(N3519), .ZN(n36445));
    INVX1 U23574 (.I(N167), .ZN(n36446));
    INVX1 U23575 (.I(N720), .ZN(n36447));
    NOR2X1 U23576 (.A1(N567), .A2(N12037), .ZN(N36448));
    NOR2X1 U23577 (.A1(N765), .A2(n22836), .ZN(n36449));
    NANDX1 U23578 (.A1(N3166), .A2(n25806), .ZN(n36450));
    NOR2X1 U23579 (.A1(N8083), .A2(N6345), .ZN(N36451));
    NANDX1 U23580 (.A1(N9501), .A2(n16845), .ZN(N36452));
    INVX1 U23581 (.I(N1890), .ZN(N36453));
    NOR2X1 U23582 (.A1(n27831), .A2(n20195), .ZN(n36454));
    INVX1 U23583 (.I(n28893), .ZN(N36455));
    INVX1 U23584 (.I(n20882), .ZN(N36456));
    INVX1 U23585 (.I(n29094), .ZN(N36457));
    INVX1 U23586 (.I(n26944), .ZN(N36458));
    INVX1 U23587 (.I(N7052), .ZN(n36459));
    NOR2X1 U23588 (.A1(N1436), .A2(N7618), .ZN(n36460));
    NANDX1 U23589 (.A1(n15360), .A2(N8382), .ZN(n36461));
    NANDX1 U23590 (.A1(n14456), .A2(N108), .ZN(n36462));
    NOR2X1 U23591 (.A1(N12780), .A2(N8191), .ZN(N36463));
    NANDX1 U23592 (.A1(N9008), .A2(n17691), .ZN(N36464));
    NANDX1 U23593 (.A1(N7650), .A2(N8141), .ZN(N36465));
    NANDX1 U23594 (.A1(N5343), .A2(n28336), .ZN(N36466));
    NOR2X1 U23595 (.A1(n22796), .A2(n19147), .ZN(N36467));
    NANDX1 U23596 (.A1(n15797), .A2(N6664), .ZN(N36468));
    NOR2X1 U23597 (.A1(N1164), .A2(N5786), .ZN(N36469));
    INVX1 U23598 (.I(n17387), .ZN(N36470));
    INVX1 U23599 (.I(n14530), .ZN(N36471));
    INVX1 U23600 (.I(n22581), .ZN(N36472));
    INVX1 U23601 (.I(N6331), .ZN(N36473));
    NANDX1 U23602 (.A1(N11580), .A2(n22957), .ZN(N36474));
    INVX1 U23603 (.I(n19770), .ZN(N36475));
    NOR2X1 U23604 (.A1(N5808), .A2(n26021), .ZN(n36476));
    INVX1 U23605 (.I(N2019), .ZN(N36477));
    NANDX1 U23606 (.A1(n24636), .A2(n26059), .ZN(N36478));
    NOR2X1 U23607 (.A1(N2094), .A2(N7279), .ZN(n36479));
    NANDX1 U23608 (.A1(N433), .A2(n23075), .ZN(N36480));
    INVX1 U23609 (.I(N11732), .ZN(N36481));
    NOR2X1 U23610 (.A1(N10940), .A2(n18644), .ZN(N36482));
    INVX1 U23611 (.I(N6722), .ZN(N36483));
    NOR2X1 U23612 (.A1(n15557), .A2(n17863), .ZN(N36484));
    INVX1 U23613 (.I(N10448), .ZN(n36485));
    NANDX1 U23614 (.A1(n26086), .A2(N3267), .ZN(n36486));
    NANDX1 U23615 (.A1(N4279), .A2(n26315), .ZN(n36487));
    NANDX1 U23616 (.A1(N163), .A2(N6025), .ZN(N36488));
    INVX1 U23617 (.I(n22885), .ZN(N36489));
    INVX1 U23618 (.I(n21128), .ZN(N36490));
    INVX1 U23619 (.I(n21315), .ZN(N36491));
    INVX1 U23620 (.I(N12158), .ZN(N36492));
    NANDX1 U23621 (.A1(N9904), .A2(n17312), .ZN(N36493));
    INVX1 U23622 (.I(n22702), .ZN(n36494));
    INVX1 U23623 (.I(N10546), .ZN(n36495));
    NOR2X1 U23624 (.A1(N4836), .A2(N2142), .ZN(n36496));
    INVX1 U23625 (.I(n22698), .ZN(N36497));
    NOR2X1 U23626 (.A1(n25876), .A2(n24580), .ZN(N36498));
    INVX1 U23627 (.I(n17703), .ZN(N36499));
    NANDX1 U23628 (.A1(n16876), .A2(N2442), .ZN(N36500));
    NOR2X1 U23629 (.A1(N5599), .A2(N8466), .ZN(N36501));
    NOR2X1 U23630 (.A1(n17044), .A2(n16248), .ZN(N36502));
    NANDX1 U23631 (.A1(N574), .A2(N7426), .ZN(N36503));
    INVX1 U23632 (.I(N12731), .ZN(n36504));
    NOR2X1 U23633 (.A1(n25063), .A2(n30043), .ZN(N36505));
    NOR2X1 U23634 (.A1(N6189), .A2(n16718), .ZN(N36506));
    NOR2X1 U23635 (.A1(n17499), .A2(n21553), .ZN(N36507));
    NANDX1 U23636 (.A1(N2789), .A2(N2674), .ZN(n36508));
    INVX1 U23637 (.I(n28664), .ZN(n36509));
    INVX1 U23638 (.I(N5812), .ZN(n36510));
    NOR2X1 U23639 (.A1(n27637), .A2(N11248), .ZN(n36511));
    NOR2X1 U23640 (.A1(n21072), .A2(N5407), .ZN(N36512));
    NOR2X1 U23641 (.A1(n21015), .A2(n22450), .ZN(n36513));
    INVX1 U23642 (.I(n19208), .ZN(n36514));
    NANDX1 U23643 (.A1(n16492), .A2(n15669), .ZN(N36515));
    NANDX1 U23644 (.A1(n22786), .A2(N10594), .ZN(N36516));
    INVX1 U23645 (.I(N9543), .ZN(n36517));
    INVX1 U23646 (.I(N10799), .ZN(N36518));
    INVX1 U23647 (.I(n22841), .ZN(N36519));
    INVX1 U23648 (.I(n13550), .ZN(n36520));
    NOR2X1 U23649 (.A1(N12146), .A2(N6764), .ZN(N36521));
    INVX1 U23650 (.I(n27960), .ZN(N36522));
    NOR2X1 U23651 (.A1(N6068), .A2(n14020), .ZN(n36523));
    NANDX1 U23652 (.A1(n13299), .A2(N4955), .ZN(N36524));
    INVX1 U23653 (.I(n17557), .ZN(N36525));
    NOR2X1 U23654 (.A1(N10101), .A2(n26623), .ZN(N36526));
    NOR2X1 U23655 (.A1(N2986), .A2(n12977), .ZN(N36527));
    INVX1 U23656 (.I(n27300), .ZN(N36528));
    NOR2X1 U23657 (.A1(n18423), .A2(N9942), .ZN(N36529));
    NOR2X1 U23658 (.A1(n23765), .A2(n20741), .ZN(n36530));
    INVX1 U23659 (.I(n16469), .ZN(N36531));
    NOR2X1 U23660 (.A1(N1245), .A2(N522), .ZN(N36532));
    NOR2X1 U23661 (.A1(N8008), .A2(N1799), .ZN(n36533));
    INVX1 U23662 (.I(N9144), .ZN(N36534));
    NOR2X1 U23663 (.A1(N12624), .A2(n21526), .ZN(n36535));
    NANDX1 U23664 (.A1(N6139), .A2(N9178), .ZN(N36536));
    NANDX1 U23665 (.A1(N9230), .A2(n19278), .ZN(N36537));
    NANDX1 U23666 (.A1(N12829), .A2(N10825), .ZN(n36538));
    NOR2X1 U23667 (.A1(n20658), .A2(N7987), .ZN(N36539));
    NOR2X1 U23668 (.A1(n27641), .A2(n17928), .ZN(N36540));
    NOR2X1 U23669 (.A1(n21268), .A2(n27229), .ZN(n36541));
    INVX1 U23670 (.I(n26297), .ZN(N36542));
    NANDX1 U23671 (.A1(N12156), .A2(n26818), .ZN(N36543));
    NANDX1 U23672 (.A1(N8724), .A2(n28617), .ZN(n36544));
    NOR2X1 U23673 (.A1(n17867), .A2(N6346), .ZN(N36545));
    NOR2X1 U23674 (.A1(N9256), .A2(n16071), .ZN(N36546));
    INVX1 U23675 (.I(N6994), .ZN(n36547));
    NOR2X1 U23676 (.A1(n24545), .A2(n26271), .ZN(N36548));
    INVX1 U23677 (.I(N7236), .ZN(N36549));
    NANDX1 U23678 (.A1(N2012), .A2(n16454), .ZN(n36550));
    INVX1 U23679 (.I(n21500), .ZN(n36551));
    NANDX1 U23680 (.A1(n28692), .A2(N3140), .ZN(N36552));
    NOR2X1 U23681 (.A1(n25783), .A2(N2612), .ZN(N36553));
    NOR2X1 U23682 (.A1(n22950), .A2(N3328), .ZN(N36554));
    INVX1 U23683 (.I(n20899), .ZN(n36555));
    NANDX1 U23684 (.A1(N3666), .A2(n28891), .ZN(N36556));
    NANDX1 U23685 (.A1(n28709), .A2(N7931), .ZN(N36557));
    INVX1 U23686 (.I(n14642), .ZN(N36558));
    NOR2X1 U23687 (.A1(N4590), .A2(n16418), .ZN(n36559));
    NOR2X1 U23688 (.A1(n19422), .A2(N11824), .ZN(N36560));
    NOR2X1 U23689 (.A1(n14940), .A2(N2396), .ZN(N36561));
    INVX1 U23690 (.I(N7006), .ZN(N36562));
    INVX1 U23691 (.I(N2283), .ZN(N36563));
    INVX1 U23692 (.I(n15596), .ZN(N36564));
    NOR2X1 U23693 (.A1(n19903), .A2(n18207), .ZN(N36565));
    NOR2X1 U23694 (.A1(N1277), .A2(n21535), .ZN(N36566));
    INVX1 U23695 (.I(n22175), .ZN(N36567));
    NOR2X1 U23696 (.A1(n13288), .A2(n20929), .ZN(n36568));
    INVX1 U23697 (.I(N420), .ZN(N36569));
    NOR2X1 U23698 (.A1(N8085), .A2(N3622), .ZN(N36570));
    NANDX1 U23699 (.A1(N1235), .A2(n20040), .ZN(N36571));
    NANDX1 U23700 (.A1(N9217), .A2(N1726), .ZN(n36572));
    INVX1 U23701 (.I(n24157), .ZN(n36573));
    NANDX1 U23702 (.A1(n29954), .A2(n19723), .ZN(n36574));
    NOR2X1 U23703 (.A1(n20798), .A2(n13843), .ZN(N36575));
    NOR2X1 U23704 (.A1(N5289), .A2(N3608), .ZN(N36576));
    INVX1 U23705 (.I(n28423), .ZN(N36577));
    NOR2X1 U23706 (.A1(n18897), .A2(N7908), .ZN(N36578));
    NANDX1 U23707 (.A1(N10906), .A2(N9756), .ZN(n36579));
    NOR2X1 U23708 (.A1(n21393), .A2(n28873), .ZN(N36580));
    NANDX1 U23709 (.A1(n18038), .A2(N2358), .ZN(n36581));
    INVX1 U23710 (.I(N7834), .ZN(n36582));
    NANDX1 U23711 (.A1(n13701), .A2(n17050), .ZN(N36583));
    INVX1 U23712 (.I(n13752), .ZN(N36584));
    INVX1 U23713 (.I(N5364), .ZN(N36585));
    NANDX1 U23714 (.A1(N7913), .A2(n21939), .ZN(n36586));
    INVX1 U23715 (.I(n21755), .ZN(N36587));
    NANDX1 U23716 (.A1(n28215), .A2(n13924), .ZN(N36588));
    NOR2X1 U23717 (.A1(n26501), .A2(N7368), .ZN(n36589));
    INVX1 U23718 (.I(n22969), .ZN(n36590));
    NANDX1 U23719 (.A1(N9560), .A2(n21286), .ZN(n36591));
    INVX1 U23720 (.I(N815), .ZN(N36592));
    NANDX1 U23721 (.A1(n23089), .A2(N7414), .ZN(n36593));
    INVX1 U23722 (.I(N8610), .ZN(N36594));
    NANDX1 U23723 (.A1(N3198), .A2(N10871), .ZN(N36595));
    INVX1 U23724 (.I(N4441), .ZN(N36596));
    NANDX1 U23725 (.A1(n20487), .A2(N9804), .ZN(N36597));
    NOR2X1 U23726 (.A1(n28399), .A2(n20304), .ZN(N36598));
    INVX1 U23727 (.I(n20017), .ZN(N36599));
    INVX1 U23728 (.I(n17618), .ZN(N36600));
    NOR2X1 U23729 (.A1(N1156), .A2(n13981), .ZN(N36601));
    NOR2X1 U23730 (.A1(n18508), .A2(n25511), .ZN(N36602));
    NANDX1 U23731 (.A1(n16628), .A2(N5220), .ZN(N36603));
    NANDX1 U23732 (.A1(N6003), .A2(n13801), .ZN(N36604));
    NANDX1 U23733 (.A1(n13416), .A2(n24740), .ZN(N36605));
    NANDX1 U23734 (.A1(n28662), .A2(n27937), .ZN(n36606));
    INVX1 U23735 (.I(n19382), .ZN(N36607));
    NANDX1 U23736 (.A1(n17455), .A2(N9731), .ZN(N36608));
    NOR2X1 U23737 (.A1(n14069), .A2(N7992), .ZN(N36609));
    NANDX1 U23738 (.A1(N3472), .A2(n16569), .ZN(N36610));
    NANDX1 U23739 (.A1(n21089), .A2(N8932), .ZN(N36611));
    NANDX1 U23740 (.A1(n23631), .A2(N8663), .ZN(n36612));
    NOR2X1 U23741 (.A1(N7565), .A2(N1243), .ZN(N36613));
    INVX1 U23742 (.I(N12784), .ZN(n36614));
    NANDX1 U23743 (.A1(n20143), .A2(n26584), .ZN(N36615));
    INVX1 U23744 (.I(N3421), .ZN(n36616));
    NOR2X1 U23745 (.A1(N8670), .A2(n20644), .ZN(N36617));
    NANDX1 U23746 (.A1(n20200), .A2(N9888), .ZN(N36618));
    NOR2X1 U23747 (.A1(N7517), .A2(N8179), .ZN(N36619));
    NOR2X1 U23748 (.A1(N10146), .A2(N4731), .ZN(n36620));
    NANDX1 U23749 (.A1(n13617), .A2(n21300), .ZN(N36621));
    INVX1 U23750 (.I(N4568), .ZN(N36622));
    NANDX1 U23751 (.A1(n25551), .A2(n16759), .ZN(N36623));
    NANDX1 U23752 (.A1(n23063), .A2(n24323), .ZN(N36624));
    NANDX1 U23753 (.A1(N7066), .A2(N6969), .ZN(N36625));
    NANDX1 U23754 (.A1(n15769), .A2(n22114), .ZN(N36626));
    NOR2X1 U23755 (.A1(n19189), .A2(n13162), .ZN(N36627));
    NANDX1 U23756 (.A1(n28393), .A2(N9269), .ZN(n36628));
    NANDX1 U23757 (.A1(n26841), .A2(n26314), .ZN(N36629));
    INVX1 U23758 (.I(N4882), .ZN(N36630));
    INVX1 U23759 (.I(N423), .ZN(n36631));
    INVX1 U23760 (.I(n29506), .ZN(n36632));
    INVX1 U23761 (.I(n19473), .ZN(N36633));
    INVX1 U23762 (.I(n25866), .ZN(N36634));
    NOR2X1 U23763 (.A1(n29887), .A2(N12487), .ZN(N36635));
    NANDX1 U23764 (.A1(n22813), .A2(N6673), .ZN(N36636));
    INVX1 U23765 (.I(n18439), .ZN(n36637));
    NANDX1 U23766 (.A1(n21599), .A2(N4070), .ZN(N36638));
    INVX1 U23767 (.I(n17069), .ZN(N36639));
    NANDX1 U23768 (.A1(n26038), .A2(N9768), .ZN(N36640));
    NOR2X1 U23769 (.A1(N5169), .A2(n22667), .ZN(n36641));
    NOR2X1 U23770 (.A1(n20044), .A2(n12944), .ZN(N36642));
    NANDX1 U23771 (.A1(N3733), .A2(N1928), .ZN(n36643));
    NOR2X1 U23772 (.A1(n21799), .A2(N4527), .ZN(N36644));
    NOR2X1 U23773 (.A1(n26135), .A2(N255), .ZN(N36645));
    NOR2X1 U23774 (.A1(n14446), .A2(N12742), .ZN(N36646));
    INVX1 U23775 (.I(n25819), .ZN(N36647));
    INVX1 U23776 (.I(n19818), .ZN(n36648));
    NANDX1 U23777 (.A1(N10176), .A2(N11279), .ZN(N36649));
    INVX1 U23778 (.I(N4354), .ZN(N36650));
    INVX1 U23779 (.I(N7129), .ZN(N36651));
    INVX1 U23780 (.I(n26676), .ZN(n36652));
    NOR2X1 U23781 (.A1(n24120), .A2(n19205), .ZN(N36653));
    NOR2X1 U23782 (.A1(n14026), .A2(n20709), .ZN(N36654));
    NANDX1 U23783 (.A1(N6319), .A2(n22636), .ZN(N36655));
    INVX1 U23784 (.I(n16678), .ZN(N36656));
    NOR2X1 U23785 (.A1(N9221), .A2(N1237), .ZN(N36657));
    INVX1 U23786 (.I(N12334), .ZN(n36658));
    NANDX1 U23787 (.A1(N5841), .A2(N9452), .ZN(n36659));
    INVX1 U23788 (.I(n13815), .ZN(n36660));
    INVX1 U23789 (.I(N2604), .ZN(N36661));
    INVX1 U23790 (.I(N10410), .ZN(N36662));
    NOR2X1 U23791 (.A1(n16905), .A2(n27318), .ZN(N36663));
    NOR2X1 U23792 (.A1(N5719), .A2(N12417), .ZN(N36664));
    NOR2X1 U23793 (.A1(n18399), .A2(N1484), .ZN(N36665));
    NOR2X1 U23794 (.A1(n20986), .A2(n22192), .ZN(N36666));
    INVX1 U23795 (.I(n15865), .ZN(N36667));
    NANDX1 U23796 (.A1(N7664), .A2(n21104), .ZN(N36668));
    INVX1 U23797 (.I(n16884), .ZN(N36669));
    NOR2X1 U23798 (.A1(N12074), .A2(n29217), .ZN(n36670));
    NANDX1 U23799 (.A1(n17915), .A2(n27229), .ZN(N36671));
    NOR2X1 U23800 (.A1(N1592), .A2(n26360), .ZN(N36672));
    NANDX1 U23801 (.A1(n14143), .A2(n25331), .ZN(N36673));
    NANDX1 U23802 (.A1(n19608), .A2(N11072), .ZN(N36674));
    NANDX1 U23803 (.A1(n13887), .A2(n23488), .ZN(N36675));
    INVX1 U23804 (.I(n20847), .ZN(n36676));
    INVX1 U23805 (.I(n16277), .ZN(N36677));
    INVX1 U23806 (.I(N5586), .ZN(N36678));
    NANDX1 U23807 (.A1(N4681), .A2(N8837), .ZN(N36679));
    NOR2X1 U23808 (.A1(n25784), .A2(n16372), .ZN(N36680));
    INVX1 U23809 (.I(n17986), .ZN(n36681));
    NANDX1 U23810 (.A1(n21894), .A2(N2991), .ZN(N36682));
    INVX1 U23811 (.I(n18985), .ZN(N36683));
    NANDX1 U23812 (.A1(N6375), .A2(N3769), .ZN(N36684));
    NOR2X1 U23813 (.A1(N9079), .A2(n29099), .ZN(n36685));
    NANDX1 U23814 (.A1(n17247), .A2(N10033), .ZN(N36686));
    INVX1 U23815 (.I(n19695), .ZN(N36687));
    INVX1 U23816 (.I(n12944), .ZN(N36688));
    INVX1 U23817 (.I(n16914), .ZN(N36689));
    NOR2X1 U23818 (.A1(N10659), .A2(N11060), .ZN(n36690));
    INVX1 U23819 (.I(N3900), .ZN(N36691));
    NANDX1 U23820 (.A1(n14721), .A2(n29684), .ZN(n36692));
    INVX1 U23821 (.I(n18836), .ZN(n36693));
    INVX1 U23822 (.I(N11698), .ZN(n36694));
    NANDX1 U23823 (.A1(N9084), .A2(n16481), .ZN(N36695));
    NANDX1 U23824 (.A1(n27139), .A2(n22856), .ZN(n36696));
    INVX1 U23825 (.I(n25467), .ZN(N36697));
    INVX1 U23826 (.I(n28126), .ZN(n36698));
    NANDX1 U23827 (.A1(N7604), .A2(N8021), .ZN(N36699));
    NANDX1 U23828 (.A1(n27298), .A2(n18662), .ZN(n36700));
    INVX1 U23829 (.I(n26262), .ZN(N36701));
    NANDX1 U23830 (.A1(n14220), .A2(n25481), .ZN(N36702));
    INVX1 U23831 (.I(N11570), .ZN(N36703));
    INVX1 U23832 (.I(n13515), .ZN(n36704));
    NANDX1 U23833 (.A1(n28927), .A2(N8207), .ZN(N36705));
    NANDX1 U23834 (.A1(N4882), .A2(N8465), .ZN(N36706));
    INVX1 U23835 (.I(N2526), .ZN(N36707));
    INVX1 U23836 (.I(n28098), .ZN(n36708));
    INVX1 U23837 (.I(n17664), .ZN(N36709));
    NOR2X1 U23838 (.A1(n13555), .A2(n26719), .ZN(n36710));
    NANDX1 U23839 (.A1(N11353), .A2(N4185), .ZN(N36711));
    NOR2X1 U23840 (.A1(n13546), .A2(n20044), .ZN(n36712));
    INVX1 U23841 (.I(n28682), .ZN(N36713));
    INVX1 U23842 (.I(N4216), .ZN(n36714));
    INVX1 U23843 (.I(N73), .ZN(N36715));
    INVX1 U23844 (.I(N1455), .ZN(N36716));
    NANDX1 U23845 (.A1(n22788), .A2(n27745), .ZN(N36717));
    NANDX1 U23846 (.A1(n19555), .A2(n19855), .ZN(N36718));
    NANDX1 U23847 (.A1(n28020), .A2(N11117), .ZN(N36719));
    NOR2X1 U23848 (.A1(n22828), .A2(N9078), .ZN(N36720));
    NOR2X1 U23849 (.A1(n29052), .A2(N6065), .ZN(N36721));
    INVX1 U23850 (.I(n14194), .ZN(N36722));
    INVX1 U23851 (.I(n25765), .ZN(N36723));
    INVX1 U23852 (.I(N11295), .ZN(N36724));
    NOR2X1 U23853 (.A1(n26982), .A2(n21513), .ZN(N36725));
    INVX1 U23854 (.I(N1574), .ZN(n36726));
    NOR2X1 U23855 (.A1(n16300), .A2(N1646), .ZN(N36727));
    INVX1 U23856 (.I(N6316), .ZN(n36728));
    NOR2X1 U23857 (.A1(n16213), .A2(N3923), .ZN(N36729));
    INVX1 U23858 (.I(n24328), .ZN(N36730));
    INVX1 U23859 (.I(n16568), .ZN(n36731));
    NOR2X1 U23860 (.A1(n23454), .A2(n17899), .ZN(n36732));
    NANDX1 U23861 (.A1(n21092), .A2(n18757), .ZN(N36733));
    NOR2X1 U23862 (.A1(n27157), .A2(N3032), .ZN(N36734));
    NOR2X1 U23863 (.A1(n16758), .A2(n17358), .ZN(N36735));
    NANDX1 U23864 (.A1(n16613), .A2(n15091), .ZN(n36736));
    NANDX1 U23865 (.A1(N7988), .A2(n30067), .ZN(N36737));
    NANDX1 U23866 (.A1(n22277), .A2(N4790), .ZN(N36738));
    NOR2X1 U23867 (.A1(n15701), .A2(N11105), .ZN(n36739));
    NANDX1 U23868 (.A1(n20474), .A2(N3588), .ZN(N36740));
    NOR2X1 U23869 (.A1(n14665), .A2(n15925), .ZN(n36741));
    NOR2X1 U23870 (.A1(n25435), .A2(n27940), .ZN(N36742));
    NANDX1 U23871 (.A1(n28896), .A2(n18894), .ZN(N36743));
    INVX1 U23872 (.I(N8392), .ZN(N36744));
    NOR2X1 U23873 (.A1(n25731), .A2(n13521), .ZN(n36745));
    NOR2X1 U23874 (.A1(n12951), .A2(n25588), .ZN(N36746));
    NOR2X1 U23875 (.A1(n28042), .A2(n23060), .ZN(N36747));
    NOR2X1 U23876 (.A1(n16532), .A2(N10667), .ZN(N36748));
    NOR2X1 U23877 (.A1(n21321), .A2(n30055), .ZN(N36749));
    NANDX1 U23878 (.A1(n20987), .A2(n27526), .ZN(n36750));
    NANDX1 U23879 (.A1(n13135), .A2(n19880), .ZN(n36751));
    INVX1 U23880 (.I(n17621), .ZN(N36752));
    NOR2X1 U23881 (.A1(n19652), .A2(n15423), .ZN(n36753));
    NOR2X1 U23882 (.A1(N6971), .A2(N4179), .ZN(N36754));
    NOR2X1 U23883 (.A1(N3923), .A2(N8653), .ZN(N36755));
    NANDX1 U23884 (.A1(n17443), .A2(N7005), .ZN(N36756));
    NOR2X1 U23885 (.A1(N1454), .A2(N3272), .ZN(n36757));
    NANDX1 U23886 (.A1(n13075), .A2(n26225), .ZN(N36758));
    NOR2X1 U23887 (.A1(N12302), .A2(n29877), .ZN(n36759));
    NANDX1 U23888 (.A1(N12219), .A2(n19093), .ZN(N36760));
    NOR2X1 U23889 (.A1(n28305), .A2(n28783), .ZN(n36761));
    NANDX1 U23890 (.A1(n18048), .A2(N11560), .ZN(n36762));
    NANDX1 U23891 (.A1(N5273), .A2(n19772), .ZN(n36763));
    INVX1 U23892 (.I(N7880), .ZN(N36764));
    INVX1 U23893 (.I(n16219), .ZN(N36765));
    NOR2X1 U23894 (.A1(n19226), .A2(n13432), .ZN(n36766));
    NOR2X1 U23895 (.A1(N6531), .A2(n20437), .ZN(N36767));
    NOR2X1 U23896 (.A1(n26683), .A2(N12269), .ZN(N36768));
    INVX1 U23897 (.I(n28318), .ZN(N36769));
    NOR2X1 U23898 (.A1(N5851), .A2(N10482), .ZN(N36770));
    NOR2X1 U23899 (.A1(n22441), .A2(N11261), .ZN(N36771));
    NOR2X1 U23900 (.A1(n18442), .A2(N9429), .ZN(n36772));
    NANDX1 U23901 (.A1(n27577), .A2(n16037), .ZN(N36773));
    INVX1 U23902 (.I(n24195), .ZN(N36774));
    NOR2X1 U23903 (.A1(N4149), .A2(N6098), .ZN(n36775));
    INVX1 U23904 (.I(n19452), .ZN(n36776));
    NANDX1 U23905 (.A1(N9359), .A2(N8540), .ZN(N36777));
    NANDX1 U23906 (.A1(N3170), .A2(N3631), .ZN(N36778));
    NANDX1 U23907 (.A1(N694), .A2(N176), .ZN(N36779));
    INVX1 U23908 (.I(n18533), .ZN(N36780));
    INVX1 U23909 (.I(N915), .ZN(n36781));
    NANDX1 U23910 (.A1(N8837), .A2(n16269), .ZN(N36782));
    NANDX1 U23911 (.A1(n20098), .A2(N1880), .ZN(N36783));
    NANDX1 U23912 (.A1(n18087), .A2(N4835), .ZN(N36784));
    NOR2X1 U23913 (.A1(N3986), .A2(n19349), .ZN(N36785));
    NOR2X1 U23914 (.A1(N2416), .A2(N12058), .ZN(N36786));
    INVX1 U23915 (.I(N8726), .ZN(N36787));
    NANDX1 U23916 (.A1(n27978), .A2(N6646), .ZN(N36788));
    NANDX1 U23917 (.A1(n29408), .A2(n28513), .ZN(N36789));
    NOR2X1 U23918 (.A1(n21137), .A2(n29207), .ZN(n36790));
    INVX1 U23919 (.I(n13696), .ZN(N36791));
    NANDX1 U23920 (.A1(n19332), .A2(N3171), .ZN(n36792));
    NANDX1 U23921 (.A1(n16729), .A2(n19439), .ZN(N36793));
    INVX1 U23922 (.I(n25387), .ZN(n36794));
    NANDX1 U23923 (.A1(n20984), .A2(n13336), .ZN(N36795));
    NANDX1 U23924 (.A1(N7794), .A2(N5882), .ZN(n36796));
    INVX1 U23925 (.I(n18798), .ZN(N36797));
    NOR2X1 U23926 (.A1(N4543), .A2(N5762), .ZN(N36798));
    NANDX1 U23927 (.A1(n24612), .A2(n22300), .ZN(N36799));
    INVX1 U23928 (.I(N4386), .ZN(n36800));
    NANDX1 U23929 (.A1(N10605), .A2(N6488), .ZN(n36801));
    NOR2X1 U23930 (.A1(n28372), .A2(N8765), .ZN(n36802));
    INVX1 U23931 (.I(n23095), .ZN(N36803));
    NOR2X1 U23932 (.A1(n17996), .A2(n19323), .ZN(N36804));
    NANDX1 U23933 (.A1(N7297), .A2(N9359), .ZN(N36805));
    NOR2X1 U23934 (.A1(N5737), .A2(N205), .ZN(N36806));
    NOR2X1 U23935 (.A1(N9010), .A2(n26696), .ZN(N36807));
    INVX1 U23936 (.I(n20193), .ZN(N36808));
    NANDX1 U23937 (.A1(N3134), .A2(n13296), .ZN(N36809));
    NOR2X1 U23938 (.A1(N8718), .A2(N7770), .ZN(N36810));
    INVX1 U23939 (.I(N9507), .ZN(N36811));
    NANDX1 U23940 (.A1(n23411), .A2(n20111), .ZN(N36812));
    NANDX1 U23941 (.A1(n24541), .A2(N6906), .ZN(N36813));
    INVX1 U23942 (.I(N9230), .ZN(n36814));
    NOR2X1 U23943 (.A1(n21185), .A2(n27225), .ZN(n36815));
    NOR2X1 U23944 (.A1(n24433), .A2(n23083), .ZN(N36816));
    INVX1 U23945 (.I(n22931), .ZN(N36817));
    NOR2X1 U23946 (.A1(N5871), .A2(N4627), .ZN(N36818));
    NOR2X1 U23947 (.A1(N2430), .A2(N10902), .ZN(n36819));
    NANDX1 U23948 (.A1(n17785), .A2(N2597), .ZN(N36820));
    INVX1 U23949 (.I(n27463), .ZN(N36821));
    INVX1 U23950 (.I(n26070), .ZN(N36822));
    INVX1 U23951 (.I(n20820), .ZN(N36823));
    INVX1 U23952 (.I(n22576), .ZN(N36824));
    NANDX1 U23953 (.A1(N3851), .A2(n16979), .ZN(N36825));
    NANDX1 U23954 (.A1(n27077), .A2(n14769), .ZN(n36826));
    INVX1 U23955 (.I(n18124), .ZN(n36827));
    NOR2X1 U23956 (.A1(n21129), .A2(N12420), .ZN(N36828));
    NANDX1 U23957 (.A1(N8097), .A2(n23911), .ZN(N36829));
    NANDX1 U23958 (.A1(N2528), .A2(n28537), .ZN(n36830));
    INVX1 U23959 (.I(N4957), .ZN(N36831));
    INVX1 U23960 (.I(N11998), .ZN(n36832));
    NOR2X1 U23961 (.A1(N458), .A2(N160), .ZN(n36833));
    NANDX1 U23962 (.A1(N332), .A2(n26229), .ZN(N36834));
    NOR2X1 U23963 (.A1(N9713), .A2(n22877), .ZN(N36835));
    NANDX1 U23964 (.A1(n27765), .A2(n15288), .ZN(n36836));
    INVX1 U23965 (.I(n22585), .ZN(n36837));
    INVX1 U23966 (.I(n20539), .ZN(n36838));
    NOR2X1 U23967 (.A1(n18911), .A2(n20956), .ZN(N36839));
    INVX1 U23968 (.I(n19891), .ZN(N36840));
    NANDX1 U23969 (.A1(N12176), .A2(n13664), .ZN(n36841));
    NOR2X1 U23970 (.A1(n14703), .A2(N624), .ZN(N36842));
    NOR2X1 U23971 (.A1(n19660), .A2(n17184), .ZN(n36843));
    NOR2X1 U23972 (.A1(N825), .A2(N6202), .ZN(n36844));
    NANDX1 U23973 (.A1(N9452), .A2(n25232), .ZN(N36845));
    INVX1 U23974 (.I(n17244), .ZN(N36846));
    NANDX1 U23975 (.A1(n24678), .A2(n17474), .ZN(n36847));
    NANDX1 U23976 (.A1(n28526), .A2(n23243), .ZN(N36848));
    INVX1 U23977 (.I(n29313), .ZN(n36849));
    NOR2X1 U23978 (.A1(N7969), .A2(n18087), .ZN(N36850));
    NANDX1 U23979 (.A1(n23487), .A2(n26538), .ZN(N36851));
    NOR2X1 U23980 (.A1(N5525), .A2(N10065), .ZN(N36852));
    NOR2X1 U23981 (.A1(n20228), .A2(n29386), .ZN(N36853));
    NOR2X1 U23982 (.A1(N9750), .A2(n16432), .ZN(N36854));
    NOR2X1 U23983 (.A1(n29272), .A2(N11195), .ZN(N36855));
    INVX1 U23984 (.I(N8586), .ZN(n36856));
    INVX1 U23985 (.I(N1618), .ZN(n36857));
    INVX1 U23986 (.I(n29793), .ZN(N36858));
    INVX1 U23987 (.I(N1726), .ZN(N36859));
    INVX1 U23988 (.I(n13245), .ZN(n36860));
    NANDX1 U23989 (.A1(N4228), .A2(N12420), .ZN(N36861));
    NANDX1 U23990 (.A1(N12197), .A2(n19067), .ZN(N36862));
    INVX1 U23991 (.I(N5546), .ZN(N36863));
    INVX1 U23992 (.I(n23355), .ZN(N36864));
    NOR2X1 U23993 (.A1(n14093), .A2(N9996), .ZN(N36865));
    NOR2X1 U23994 (.A1(n13341), .A2(n13069), .ZN(N36866));
    NOR2X1 U23995 (.A1(n18334), .A2(n14434), .ZN(N36867));
    NOR2X1 U23996 (.A1(n18089), .A2(n21508), .ZN(n36868));
    NOR2X1 U23997 (.A1(n24377), .A2(N11686), .ZN(N36869));
    INVX1 U23998 (.I(N12593), .ZN(N36870));
    INVX1 U23999 (.I(n19124), .ZN(N36871));
    NOR2X1 U24000 (.A1(n28347), .A2(N2515), .ZN(N36872));
    NANDX1 U24001 (.A1(N10629), .A2(N6809), .ZN(N36873));
    INVX1 U24002 (.I(n29696), .ZN(N36874));
    NANDX1 U24003 (.A1(n13772), .A2(N3587), .ZN(n36875));
    NOR2X1 U24004 (.A1(n13403), .A2(n17679), .ZN(n36876));
    NANDX1 U24005 (.A1(n21822), .A2(n19580), .ZN(n36877));
    NOR2X1 U24006 (.A1(n28551), .A2(N7776), .ZN(n36878));
    NOR2X1 U24007 (.A1(N4277), .A2(n14425), .ZN(N36879));
    NOR2X1 U24008 (.A1(n18725), .A2(n27362), .ZN(N36880));
    NOR2X1 U24009 (.A1(N5986), .A2(N9817), .ZN(N36881));
    INVX1 U24010 (.I(n25109), .ZN(N36882));
    NANDX1 U24011 (.A1(n16890), .A2(n16184), .ZN(n36883));
    NANDX1 U24012 (.A1(n27518), .A2(N11554), .ZN(n36884));
    NANDX1 U24013 (.A1(n15637), .A2(n15679), .ZN(n36885));
    NOR2X1 U24014 (.A1(n19223), .A2(N1582), .ZN(N36886));
    INVX1 U24015 (.I(N6764), .ZN(N36887));
    NOR2X1 U24016 (.A1(n17472), .A2(n26344), .ZN(N36888));
    NOR2X1 U24017 (.A1(N4446), .A2(n22680), .ZN(N36889));
    NANDX1 U24018 (.A1(N8722), .A2(N6968), .ZN(N36890));
    NOR2X1 U24019 (.A1(n16007), .A2(n22890), .ZN(N36891));
    NANDX1 U24020 (.A1(n21992), .A2(N2570), .ZN(N36892));
    NOR2X1 U24021 (.A1(N5524), .A2(n15627), .ZN(N36893));
    INVX1 U24022 (.I(N10269), .ZN(n36894));
    INVX1 U24023 (.I(n27029), .ZN(n36895));
    NANDX1 U24024 (.A1(n16070), .A2(N12529), .ZN(N36896));
    INVX1 U24025 (.I(n28455), .ZN(N36897));
    INVX1 U24026 (.I(n16203), .ZN(N36898));
    NANDX1 U24027 (.A1(n27076), .A2(N2243), .ZN(n36899));
    NOR2X1 U24028 (.A1(N11843), .A2(n23208), .ZN(N36900));
    NANDX1 U24029 (.A1(n23083), .A2(n14557), .ZN(n36901));
    NANDX1 U24030 (.A1(n18611), .A2(n27936), .ZN(N36902));
    NANDX1 U24031 (.A1(N11364), .A2(N3317), .ZN(n36903));
    INVX1 U24032 (.I(n13933), .ZN(n36904));
    INVX1 U24033 (.I(n22373), .ZN(n36905));
    NANDX1 U24034 (.A1(n27026), .A2(N2504), .ZN(N36906));
    NOR2X1 U24035 (.A1(n23918), .A2(n12886), .ZN(N36907));
    NOR2X1 U24036 (.A1(n25007), .A2(N8809), .ZN(N36908));
    NOR2X1 U24037 (.A1(n15181), .A2(n25011), .ZN(N36909));
    NANDX1 U24038 (.A1(N680), .A2(n15814), .ZN(N36910));
    NANDX1 U24039 (.A1(N1083), .A2(N8884), .ZN(N36911));
    NOR2X1 U24040 (.A1(n24166), .A2(n23441), .ZN(N36912));
    NANDX1 U24041 (.A1(N1200), .A2(n21239), .ZN(n36913));
    NOR2X1 U24042 (.A1(N12563), .A2(n13117), .ZN(n36914));
    NANDX1 U24043 (.A1(n15056), .A2(N10494), .ZN(N36915));
    NANDX1 U24044 (.A1(N3039), .A2(N7383), .ZN(N36916));
    NOR2X1 U24045 (.A1(n27174), .A2(n19861), .ZN(N36917));
    NOR2X1 U24046 (.A1(N7104), .A2(n14730), .ZN(N36918));
    INVX1 U24047 (.I(n22747), .ZN(n36919));
    NOR2X1 U24048 (.A1(N4480), .A2(n20920), .ZN(N36920));
    NOR2X1 U24049 (.A1(N8854), .A2(n26352), .ZN(N36921));
    NOR2X1 U24050 (.A1(n17738), .A2(N6093), .ZN(N36922));
    INVX1 U24051 (.I(n29739), .ZN(N36923));
    INVX1 U24052 (.I(n15461), .ZN(n36924));
    NOR2X1 U24053 (.A1(N1285), .A2(n16584), .ZN(N36925));
    NOR2X1 U24054 (.A1(N5899), .A2(n20201), .ZN(N36926));
    NANDX1 U24055 (.A1(n21446), .A2(n23239), .ZN(n36927));
    NANDX1 U24056 (.A1(n20798), .A2(n20275), .ZN(N36928));
    INVX1 U24057 (.I(n21596), .ZN(N36929));
    NOR2X1 U24058 (.A1(n21967), .A2(N1065), .ZN(N36930));
    INVX1 U24059 (.I(N10300), .ZN(N36931));
    NOR2X1 U24060 (.A1(n18028), .A2(n29450), .ZN(N36932));
    INVX1 U24061 (.I(n14242), .ZN(N36933));
    NOR2X1 U24062 (.A1(N9256), .A2(N8895), .ZN(N36934));
    NOR2X1 U24063 (.A1(N8857), .A2(N3716), .ZN(n36935));
    NANDX1 U24064 (.A1(n18258), .A2(n23698), .ZN(N36936));
    NANDX1 U24065 (.A1(n29335), .A2(n29596), .ZN(N36937));
    INVX1 U24066 (.I(n20769), .ZN(N36938));
    NOR2X1 U24067 (.A1(n26136), .A2(N8146), .ZN(N36939));
    INVX1 U24068 (.I(n16273), .ZN(n36940));
    NANDX1 U24069 (.A1(N10281), .A2(n20772), .ZN(n36941));
    INVX1 U24070 (.I(n30043), .ZN(n36942));
    NANDX1 U24071 (.A1(N6073), .A2(n24147), .ZN(n36943));
    NANDX1 U24072 (.A1(n24083), .A2(n15665), .ZN(n36944));
    NOR2X1 U24073 (.A1(n13491), .A2(n24921), .ZN(n36945));
    NOR2X1 U24074 (.A1(N5721), .A2(n22338), .ZN(N36946));
    INVX1 U24075 (.I(N1971), .ZN(n36947));
    NANDX1 U24076 (.A1(N3304), .A2(n14805), .ZN(N36948));
    INVX1 U24077 (.I(n21460), .ZN(N36949));
    INVX1 U24078 (.I(N7546), .ZN(N36950));
    NANDX1 U24079 (.A1(N2261), .A2(N4253), .ZN(N36951));
    NANDX1 U24080 (.A1(N7094), .A2(N8196), .ZN(N36952));
    NOR2X1 U24081 (.A1(n27865), .A2(N3969), .ZN(n36953));
    NOR2X1 U24082 (.A1(n15608), .A2(n28739), .ZN(N36954));
    INVX1 U24083 (.I(n21378), .ZN(N36955));
    NOR2X1 U24084 (.A1(n28028), .A2(n29950), .ZN(N36956));
    INVX1 U24085 (.I(n22811), .ZN(n36957));
    NOR2X1 U24086 (.A1(N319), .A2(n15012), .ZN(N36958));
    INVX1 U24087 (.I(N2289), .ZN(N36959));
    NANDX1 U24088 (.A1(N7448), .A2(n17094), .ZN(N36960));
    NOR2X1 U24089 (.A1(n17468), .A2(n23356), .ZN(N36961));
    INVX1 U24090 (.I(n18254), .ZN(N36962));
    NOR2X1 U24091 (.A1(N12605), .A2(N7725), .ZN(n36963));
    INVX1 U24092 (.I(n20800), .ZN(N36964));
    NANDX1 U24093 (.A1(N7560), .A2(n13329), .ZN(n36965));
    INVX1 U24094 (.I(n23167), .ZN(n36966));
    NANDX1 U24095 (.A1(n19495), .A2(N2968), .ZN(N36967));
    NOR2X1 U24096 (.A1(n17386), .A2(n21478), .ZN(n36968));
    NOR2X1 U24097 (.A1(N10059), .A2(n15880), .ZN(n36969));
    NOR2X1 U24098 (.A1(n25070), .A2(n20024), .ZN(N36970));
    NOR2X1 U24099 (.A1(n27661), .A2(n16033), .ZN(n36971));
    INVX1 U24100 (.I(n28467), .ZN(N36972));
    NANDX1 U24101 (.A1(n26511), .A2(N6682), .ZN(n36973));
    NOR2X1 U24102 (.A1(n29249), .A2(N7847), .ZN(n36974));
    INVX1 U24103 (.I(N8943), .ZN(n36975));
    NOR2X1 U24104 (.A1(n25378), .A2(n16502), .ZN(n36976));
    INVX1 U24105 (.I(N2372), .ZN(N36977));
    NOR2X1 U24106 (.A1(N890), .A2(n21867), .ZN(N36978));
    NANDX1 U24107 (.A1(N1186), .A2(N9115), .ZN(n36979));
    INVX1 U24108 (.I(N7519), .ZN(N36980));
    INVX1 U24109 (.I(n15538), .ZN(N36981));
    INVX1 U24110 (.I(n21365), .ZN(N36982));
    NOR2X1 U24111 (.A1(N11670), .A2(n18888), .ZN(n36983));
    NOR2X1 U24112 (.A1(n14825), .A2(n17217), .ZN(n36984));
    NOR2X1 U24113 (.A1(n29896), .A2(N12460), .ZN(N36985));
    NANDX1 U24114 (.A1(n17568), .A2(N8867), .ZN(n36986));
    NANDX1 U24115 (.A1(n26510), .A2(n26074), .ZN(n36987));
    NANDX1 U24116 (.A1(n12875), .A2(n26473), .ZN(n36988));
    NANDX1 U24117 (.A1(n29664), .A2(n15923), .ZN(n36989));
    INVX1 U24118 (.I(n19284), .ZN(N36990));
    NOR2X1 U24119 (.A1(n17035), .A2(n18942), .ZN(N36991));
    NANDX1 U24120 (.A1(n24768), .A2(N4342), .ZN(N36992));
    NANDX1 U24121 (.A1(n15995), .A2(N9765), .ZN(n36993));
    NANDX1 U24122 (.A1(n23443), .A2(n19782), .ZN(n36994));
    NOR2X1 U24123 (.A1(n29221), .A2(n21722), .ZN(N36995));
    INVX1 U24124 (.I(N11543), .ZN(n36996));
    INVX1 U24125 (.I(N6720), .ZN(n36997));
    NANDX1 U24126 (.A1(n15022), .A2(N3093), .ZN(N36998));
    NANDX1 U24127 (.A1(N10144), .A2(N4528), .ZN(N36999));
    NOR2X1 U24128 (.A1(N7637), .A2(N4054), .ZN(N37000));
    NOR2X1 U24129 (.A1(N4118), .A2(n23337), .ZN(N37001));
    NOR2X1 U24130 (.A1(n21152), .A2(N12141), .ZN(N37002));
    INVX1 U24131 (.I(N4343), .ZN(N37003));
    INVX1 U24132 (.I(N10358), .ZN(N37004));
    NANDX1 U24133 (.A1(n14808), .A2(n26504), .ZN(n37005));
    NANDX1 U24134 (.A1(n23150), .A2(n15899), .ZN(N37006));
    INVX1 U24135 (.I(n14734), .ZN(n37007));
    INVX1 U24136 (.I(n20088), .ZN(n37008));
    NOR2X1 U24137 (.A1(N332), .A2(n29058), .ZN(n37009));
    NANDX1 U24138 (.A1(n22122), .A2(N3827), .ZN(n37010));
    NOR2X1 U24139 (.A1(n15210), .A2(n23766), .ZN(N37011));
    NOR2X1 U24140 (.A1(n19263), .A2(n18051), .ZN(n37012));
    NOR2X1 U24141 (.A1(N1024), .A2(n18004), .ZN(N37013));
    INVX1 U24142 (.I(N1725), .ZN(N37014));
    INVX1 U24143 (.I(n16392), .ZN(n37015));
    NANDX1 U24144 (.A1(N11363), .A2(n25290), .ZN(N37016));
    NANDX1 U24145 (.A1(n26427), .A2(N4615), .ZN(N37017));
    INVX1 U24146 (.I(N749), .ZN(N37018));
    NANDX1 U24147 (.A1(N6442), .A2(n24498), .ZN(N37019));
    NOR2X1 U24148 (.A1(n24876), .A2(n13390), .ZN(N37020));
    INVX1 U24149 (.I(n28194), .ZN(N37021));
    NOR2X1 U24150 (.A1(N5857), .A2(N80), .ZN(n37022));
    NANDX1 U24151 (.A1(n18183), .A2(n28436), .ZN(N37023));
    NANDX1 U24152 (.A1(N6096), .A2(N12075), .ZN(N37024));
    INVX1 U24153 (.I(n24099), .ZN(N37025));
    NANDX1 U24154 (.A1(n19715), .A2(n25104), .ZN(N37026));
    NANDX1 U24155 (.A1(n15043), .A2(n25027), .ZN(n37027));
    INVX1 U24156 (.I(n25178), .ZN(N37028));
    NANDX1 U24157 (.A1(n28842), .A2(n16886), .ZN(N37029));
    NANDX1 U24158 (.A1(N11865), .A2(n23327), .ZN(n37030));
    NANDX1 U24159 (.A1(n26414), .A2(n18065), .ZN(N37031));
    INVX1 U24160 (.I(n28445), .ZN(N37032));
    INVX1 U24161 (.I(n23748), .ZN(n37033));
    NOR2X1 U24162 (.A1(N4761), .A2(N2754), .ZN(n37034));
    NOR2X1 U24163 (.A1(N3060), .A2(N1023), .ZN(N37035));
    NOR2X1 U24164 (.A1(N3695), .A2(n19012), .ZN(n37036));
    NOR2X1 U24165 (.A1(n16378), .A2(n27287), .ZN(N37037));
    INVX1 U24166 (.I(n15316), .ZN(N37038));
    NOR2X1 U24167 (.A1(N8080), .A2(N9405), .ZN(N37039));
    NANDX1 U24168 (.A1(n17957), .A2(n26807), .ZN(n37040));
    NANDX1 U24169 (.A1(n28582), .A2(N8534), .ZN(n37041));
    NANDX1 U24170 (.A1(N3431), .A2(n23509), .ZN(N37042));
    NANDX1 U24171 (.A1(N10366), .A2(N10377), .ZN(N37043));
    NOR2X1 U24172 (.A1(n22675), .A2(n21799), .ZN(N37044));
    INVX1 U24173 (.I(n25428), .ZN(n37045));
    NANDX1 U24174 (.A1(n13554), .A2(n15011), .ZN(N37046));
    NANDX1 U24175 (.A1(n17248), .A2(n22584), .ZN(n37047));
    NANDX1 U24176 (.A1(n22187), .A2(n19733), .ZN(N37048));
    NOR2X1 U24177 (.A1(N7365), .A2(n20486), .ZN(n37049));
    NANDX1 U24178 (.A1(N5330), .A2(n27717), .ZN(n37050));
    INVX1 U24179 (.I(N2000), .ZN(n37051));
    NOR2X1 U24180 (.A1(n29708), .A2(n29231), .ZN(N37052));
    INVX1 U24181 (.I(n21699), .ZN(N37053));
    NOR2X1 U24182 (.A1(n28616), .A2(N1927), .ZN(N37054));
    NANDX1 U24183 (.A1(n15652), .A2(n24601), .ZN(N37055));
    NANDX1 U24184 (.A1(N7448), .A2(N8453), .ZN(n37056));
    INVX1 U24185 (.I(n21002), .ZN(n37057));
    NOR2X1 U24186 (.A1(N1023), .A2(n26810), .ZN(n37058));
    NANDX1 U24187 (.A1(n15939), .A2(n18859), .ZN(N37059));
    INVX1 U24188 (.I(n13908), .ZN(n37060));
    NOR2X1 U24189 (.A1(N3112), .A2(N8516), .ZN(N37061));
    NOR2X1 U24190 (.A1(n19389), .A2(n21081), .ZN(n37062));
    NANDX1 U24191 (.A1(n18207), .A2(n20651), .ZN(N37063));
    NOR2X1 U24192 (.A1(n22892), .A2(N12212), .ZN(n37064));
    NOR2X1 U24193 (.A1(n21370), .A2(n14138), .ZN(N37065));
    NANDX1 U24194 (.A1(N6884), .A2(n27300), .ZN(N37066));
    NOR2X1 U24195 (.A1(N2892), .A2(N5615), .ZN(N37067));
    NANDX1 U24196 (.A1(n23893), .A2(N6199), .ZN(N37068));
    NANDX1 U24197 (.A1(N9127), .A2(N10669), .ZN(n37069));
    INVX1 U24198 (.I(n27985), .ZN(N37070));
    NANDX1 U24199 (.A1(n26412), .A2(N12632), .ZN(N37071));
    INVX1 U24200 (.I(N4790), .ZN(n37072));
    NOR2X1 U24201 (.A1(n23053), .A2(n14431), .ZN(n37073));
    NANDX1 U24202 (.A1(n29821), .A2(N4944), .ZN(n37074));
    INVX1 U24203 (.I(n22575), .ZN(N37075));
    NANDX1 U24204 (.A1(N2400), .A2(n13807), .ZN(n37076));
    NANDX1 U24205 (.A1(N3292), .A2(N9251), .ZN(n37077));
    NANDX1 U24206 (.A1(N5944), .A2(N12142), .ZN(n37078));
    INVX1 U24207 (.I(n12926), .ZN(N37079));
    INVX1 U24208 (.I(N5950), .ZN(n37080));
    NOR2X1 U24209 (.A1(N3585), .A2(N5179), .ZN(n37081));
    INVX1 U24210 (.I(n20130), .ZN(n37082));
    INVX1 U24211 (.I(N6831), .ZN(N37083));
    NOR2X1 U24212 (.A1(n20835), .A2(N181), .ZN(N37084));
    NOR2X1 U24213 (.A1(N2312), .A2(n14612), .ZN(N37085));
    INVX1 U24214 (.I(N1995), .ZN(n37086));
    NANDX1 U24215 (.A1(n18680), .A2(n24569), .ZN(N37087));
    INVX1 U24216 (.I(n21079), .ZN(N37088));
    NANDX1 U24217 (.A1(N3548), .A2(n24370), .ZN(N37089));
    INVX1 U24218 (.I(N9124), .ZN(N37090));
    NANDX1 U24219 (.A1(N6751), .A2(n27573), .ZN(N37091));
    NOR2X1 U24220 (.A1(N1209), .A2(N3385), .ZN(N37092));
    NOR2X1 U24221 (.A1(N4793), .A2(N8564), .ZN(N37093));
    NOR2X1 U24222 (.A1(n24923), .A2(n25734), .ZN(N37094));
    NANDX1 U24223 (.A1(n16107), .A2(N4993), .ZN(n37095));
    NOR2X1 U24224 (.A1(N9899), .A2(N7304), .ZN(n37096));
    NANDX1 U24225 (.A1(N5531), .A2(N9298), .ZN(N37097));
    NOR2X1 U24226 (.A1(n24210), .A2(n22427), .ZN(n37098));
    INVX1 U24227 (.I(N3713), .ZN(N37099));
    INVX1 U24228 (.I(n23069), .ZN(N37100));
    NOR2X1 U24229 (.A1(n13834), .A2(n20753), .ZN(n37101));
    NANDX1 U24230 (.A1(n20584), .A2(n18188), .ZN(n37102));
    NOR2X1 U24231 (.A1(N10354), .A2(n21573), .ZN(N37103));
    NANDX1 U24232 (.A1(n15146), .A2(n30136), .ZN(n37104));
    NOR2X1 U24233 (.A1(n28629), .A2(n14293), .ZN(n37105));
    INVX1 U24234 (.I(N3160), .ZN(n37106));
    NOR2X1 U24235 (.A1(N5653), .A2(N1619), .ZN(n37107));
    NANDX1 U24236 (.A1(n14667), .A2(N7149), .ZN(N37108));
    INVX1 U24237 (.I(n20358), .ZN(N37109));
    INVX1 U24238 (.I(N5296), .ZN(n37110));
    NOR2X1 U24239 (.A1(n23632), .A2(n13081), .ZN(N37111));
    INVX1 U24240 (.I(N10137), .ZN(n37112));
    NOR2X1 U24241 (.A1(n23426), .A2(n15517), .ZN(N37113));
    NOR2X1 U24242 (.A1(N11477), .A2(n22559), .ZN(n37114));
    NANDX1 U24243 (.A1(N2912), .A2(n17876), .ZN(N37115));
    NANDX1 U24244 (.A1(N2910), .A2(n23464), .ZN(n37116));
    INVX1 U24245 (.I(n17202), .ZN(N37117));
    INVX1 U24246 (.I(N10193), .ZN(n37118));
    NANDX1 U24247 (.A1(n28927), .A2(N11811), .ZN(n37119));
    NOR2X1 U24248 (.A1(N2018), .A2(N7520), .ZN(N37120));
    NANDX1 U24249 (.A1(N10936), .A2(n16000), .ZN(N37121));
    NANDX1 U24250 (.A1(N1979), .A2(n28192), .ZN(n37122));
    INVX1 U24251 (.I(N4652), .ZN(N37123));
    NANDX1 U24252 (.A1(n26779), .A2(n28078), .ZN(N37124));
    NOR2X1 U24253 (.A1(N2563), .A2(n28115), .ZN(N37125));
    INVX1 U24254 (.I(n18837), .ZN(n37126));
    NANDX1 U24255 (.A1(n22565), .A2(N8681), .ZN(n37127));
    NANDX1 U24256 (.A1(N4453), .A2(n15714), .ZN(N37128));
    NOR2X1 U24257 (.A1(n27727), .A2(n25906), .ZN(n37129));
    INVX1 U24258 (.I(n15077), .ZN(n37130));
    NANDX1 U24259 (.A1(N3090), .A2(N5655), .ZN(N37131));
    INVX1 U24260 (.I(n14716), .ZN(n37132));
    NANDX1 U24261 (.A1(N8220), .A2(n12939), .ZN(n37133));
    NOR2X1 U24262 (.A1(N6274), .A2(N12804), .ZN(n37134));
    INVX1 U24263 (.I(n14465), .ZN(n37135));
    INVX1 U24264 (.I(n16980), .ZN(n37136));
    NOR2X1 U24265 (.A1(N569), .A2(n14957), .ZN(N37137));
    INVX1 U24266 (.I(n19406), .ZN(n37138));
    INVX1 U24267 (.I(N972), .ZN(N37139));
    NOR2X1 U24268 (.A1(n26901), .A2(N5424), .ZN(N37140));
    NOR2X1 U24269 (.A1(n25022), .A2(n21711), .ZN(N37141));
    INVX1 U24270 (.I(n18052), .ZN(N37142));
    NANDX1 U24271 (.A1(n24267), .A2(N9702), .ZN(n37143));
    NANDX1 U24272 (.A1(n16486), .A2(n24417), .ZN(N37144));
    NOR2X1 U24273 (.A1(n24705), .A2(n25917), .ZN(N37145));
    NOR2X1 U24274 (.A1(N842), .A2(n27281), .ZN(n37146));
    NANDX1 U24275 (.A1(N3867), .A2(n25287), .ZN(n37147));
    NOR2X1 U24276 (.A1(n19161), .A2(n25856), .ZN(N37148));
    NOR2X1 U24277 (.A1(N9006), .A2(N3685), .ZN(N37149));
    NOR2X1 U24278 (.A1(n28675), .A2(n20331), .ZN(N37150));
    NANDX1 U24279 (.A1(N3961), .A2(n22553), .ZN(n37151));
    INVX1 U24280 (.I(n14232), .ZN(N37152));
    NANDX1 U24281 (.A1(n13771), .A2(n28141), .ZN(N37153));
    INVX1 U24282 (.I(N12034), .ZN(N37154));
    NOR2X1 U24283 (.A1(n19718), .A2(n25011), .ZN(N37155));
    NANDX1 U24284 (.A1(n14286), .A2(n20790), .ZN(N37156));
    NOR2X1 U24285 (.A1(N3688), .A2(N6495), .ZN(N37157));
    INVX1 U24286 (.I(n26252), .ZN(N37158));
    NANDX1 U24287 (.A1(N605), .A2(n15275), .ZN(N37159));
    NOR2X1 U24288 (.A1(N271), .A2(N12842), .ZN(n37160));
    NANDX1 U24289 (.A1(n15782), .A2(N11379), .ZN(N37161));
    NOR2X1 U24290 (.A1(n16617), .A2(N3901), .ZN(N37162));
    NANDX1 U24291 (.A1(N12336), .A2(n18132), .ZN(N37163));
    NOR2X1 U24292 (.A1(n14667), .A2(n16135), .ZN(N37164));
    NOR2X1 U24293 (.A1(n26700), .A2(N3564), .ZN(N37165));
    NOR2X1 U24294 (.A1(n21574), .A2(n15707), .ZN(N37166));
    NANDX1 U24295 (.A1(N787), .A2(n18116), .ZN(N37167));
    NANDX1 U24296 (.A1(n25979), .A2(N11133), .ZN(n37168));
    NANDX1 U24297 (.A1(n27623), .A2(N298), .ZN(N37169));
    INVX1 U24298 (.I(N2106), .ZN(N37170));
    NANDX1 U24299 (.A1(N12153), .A2(n29109), .ZN(N37171));
    NOR2X1 U24300 (.A1(N12092), .A2(n27606), .ZN(n37172));
    NANDX1 U24301 (.A1(n15992), .A2(N7080), .ZN(N37173));
    INVX1 U24302 (.I(N3987), .ZN(n37174));
    NANDX1 U24303 (.A1(N6952), .A2(N8682), .ZN(n37175));
    NOR2X1 U24304 (.A1(N3515), .A2(N807), .ZN(N37176));
    NOR2X1 U24305 (.A1(n13649), .A2(N5074), .ZN(N37177));
    INVX1 U24306 (.I(N2996), .ZN(n37178));
    INVX1 U24307 (.I(N12724), .ZN(N37179));
    NANDX1 U24308 (.A1(n22882), .A2(n15458), .ZN(N37180));
    NOR2X1 U24309 (.A1(n23179), .A2(n14769), .ZN(N37181));
    INVX1 U24310 (.I(n23747), .ZN(N37182));
    NOR2X1 U24311 (.A1(N4658), .A2(n28657), .ZN(n37183));
    INVX1 U24312 (.I(n20825), .ZN(n37184));
    NANDX1 U24313 (.A1(n13428), .A2(n16465), .ZN(N37185));
    NOR2X1 U24314 (.A1(N5975), .A2(N12120), .ZN(N37186));
    NOR2X1 U24315 (.A1(N3218), .A2(n29721), .ZN(N37187));
    INVX1 U24316 (.I(n22722), .ZN(n37188));
    INVX1 U24317 (.I(n13567), .ZN(n37189));
    NOR2X1 U24318 (.A1(N11936), .A2(N5123), .ZN(n37190));
    INVX1 U24319 (.I(n13220), .ZN(n37191));
    NANDX1 U24320 (.A1(n20849), .A2(n28678), .ZN(N37192));
    NANDX1 U24321 (.A1(N2451), .A2(N1870), .ZN(N37193));
    NOR2X1 U24322 (.A1(n14759), .A2(N5913), .ZN(N37194));
    INVX1 U24323 (.I(N1839), .ZN(N37195));
    NOR2X1 U24324 (.A1(n27270), .A2(N10446), .ZN(N37196));
    INVX1 U24325 (.I(n13597), .ZN(N37197));
    NOR2X1 U24326 (.A1(n30010), .A2(n14278), .ZN(N37198));
    NOR2X1 U24327 (.A1(N3090), .A2(N2422), .ZN(N37199));
    NOR2X1 U24328 (.A1(n14372), .A2(n19694), .ZN(N37200));
    INVX1 U24329 (.I(N12029), .ZN(N37201));
    NANDX1 U24330 (.A1(n14909), .A2(N9996), .ZN(N37202));
    NOR2X1 U24331 (.A1(N7429), .A2(n19405), .ZN(n37203));
    INVX1 U24332 (.I(N3531), .ZN(N37204));
    INVX1 U24333 (.I(N10941), .ZN(N37205));
    INVX1 U24334 (.I(N6476), .ZN(N37206));
    NANDX1 U24335 (.A1(N11764), .A2(N8315), .ZN(n37207));
    INVX1 U24336 (.I(n27595), .ZN(n37208));
    NANDX1 U24337 (.A1(N2660), .A2(n29752), .ZN(n37209));
    INVX1 U24338 (.I(N2532), .ZN(n37210));
    INVX1 U24339 (.I(n26398), .ZN(N37211));
    NOR2X1 U24340 (.A1(N4875), .A2(n22617), .ZN(N37212));
    NANDX1 U24341 (.A1(n13129), .A2(N2266), .ZN(N37213));
    INVX1 U24342 (.I(N3181), .ZN(N37214));
    NOR2X1 U24343 (.A1(N7698), .A2(n25151), .ZN(N37215));
    INVX1 U24344 (.I(n15663), .ZN(N37216));
    INVX1 U24345 (.I(n16693), .ZN(n37217));
    NANDX1 U24346 (.A1(N3587), .A2(n22011), .ZN(N37218));
    NANDX1 U24347 (.A1(N9000), .A2(n22336), .ZN(n37219));
    NOR2X1 U24348 (.A1(N6323), .A2(n19793), .ZN(N37220));
    INVX1 U24349 (.I(n27680), .ZN(n37221));
    NANDX1 U24350 (.A1(n13829), .A2(n18772), .ZN(N37222));
    INVX1 U24351 (.I(n28787), .ZN(n37223));
    INVX1 U24352 (.I(n26734), .ZN(n37224));
    INVX1 U24353 (.I(N10066), .ZN(n37225));
    INVX1 U24354 (.I(n23532), .ZN(N37226));
    INVX1 U24355 (.I(N1466), .ZN(n37227));
    NANDX1 U24356 (.A1(N4026), .A2(n15178), .ZN(N37228));
    NANDX1 U24357 (.A1(n19688), .A2(N7823), .ZN(n37229));
    NOR2X1 U24358 (.A1(n15628), .A2(n30107), .ZN(N37230));
    INVX1 U24359 (.I(N6605), .ZN(N37231));
    INVX1 U24360 (.I(N1616), .ZN(N37232));
    NANDX1 U24361 (.A1(N3853), .A2(n21408), .ZN(n37233));
    NANDX1 U24362 (.A1(n20093), .A2(n29376), .ZN(N37234));
    INVX1 U24363 (.I(N8727), .ZN(N37235));
    NANDX1 U24364 (.A1(n24985), .A2(N10240), .ZN(n37236));
    NOR2X1 U24365 (.A1(N4675), .A2(n20305), .ZN(N37237));
    INVX1 U24366 (.I(n28206), .ZN(N37238));
    NOR2X1 U24367 (.A1(N6005), .A2(n27334), .ZN(N37239));
    NOR2X1 U24368 (.A1(n21182), .A2(n28186), .ZN(n37240));
    NANDX1 U24369 (.A1(n29005), .A2(n15593), .ZN(n37241));
    NOR2X1 U24370 (.A1(n28974), .A2(n25010), .ZN(N37242));
    NOR2X1 U24371 (.A1(n26504), .A2(n26626), .ZN(N37243));
    INVX1 U24372 (.I(n18917), .ZN(N37244));
    NANDX1 U24373 (.A1(n16525), .A2(N8872), .ZN(N37245));
    NOR2X1 U24374 (.A1(N1284), .A2(n17598), .ZN(n37246));
    INVX1 U24375 (.I(n14829), .ZN(N37247));
    NOR2X1 U24376 (.A1(N2909), .A2(n19504), .ZN(N37248));
    NANDX1 U24377 (.A1(N7448), .A2(n17572), .ZN(N37249));
    NANDX1 U24378 (.A1(n13453), .A2(N3330), .ZN(n37250));
    NANDX1 U24379 (.A1(n23195), .A2(N1378), .ZN(N37251));
    NOR2X1 U24380 (.A1(n22062), .A2(n16970), .ZN(N37252));
    NOR2X1 U24381 (.A1(N9460), .A2(N403), .ZN(N37253));
    NOR2X1 U24382 (.A1(N5826), .A2(n15589), .ZN(N37254));
    INVX1 U24383 (.I(n13304), .ZN(n37255));
    NANDX1 U24384 (.A1(N11227), .A2(n22175), .ZN(N37256));
    NANDX1 U24385 (.A1(N12510), .A2(n28334), .ZN(n37257));
    INVX1 U24386 (.I(n15900), .ZN(n37258));
    INVX1 U24387 (.I(n23123), .ZN(n37259));
    INVX1 U24388 (.I(n21159), .ZN(N37260));
    INVX1 U24389 (.I(N11398), .ZN(n37261));
    INVX1 U24390 (.I(N2447), .ZN(n37262));
    NOR2X1 U24391 (.A1(N12316), .A2(n25641), .ZN(n37263));
    INVX1 U24392 (.I(N1922), .ZN(N37264));
    NOR2X1 U24393 (.A1(N10195), .A2(n13183), .ZN(N37265));
    NOR2X1 U24394 (.A1(N10598), .A2(n22566), .ZN(N37266));
    NANDX1 U24395 (.A1(n14747), .A2(n17269), .ZN(N37267));
    INVX1 U24396 (.I(N6655), .ZN(n37268));
    INVX1 U24397 (.I(N3874), .ZN(N37269));
    NANDX1 U24398 (.A1(n29566), .A2(N2070), .ZN(n37270));
    NANDX1 U24399 (.A1(n15328), .A2(n16663), .ZN(N37271));
    INVX1 U24400 (.I(N9154), .ZN(N37272));
    INVX1 U24401 (.I(n25149), .ZN(N37273));
    INVX1 U24402 (.I(n17722), .ZN(N37274));
    INVX1 U24403 (.I(n23839), .ZN(N37275));
    NOR2X1 U24404 (.A1(N11660), .A2(n17064), .ZN(N37276));
    NANDX1 U24405 (.A1(N6347), .A2(n27259), .ZN(N37277));
    NOR2X1 U24406 (.A1(n21932), .A2(n26417), .ZN(N37278));
    NANDX1 U24407 (.A1(N1766), .A2(N11026), .ZN(N37279));
    NOR2X1 U24408 (.A1(n13602), .A2(N6242), .ZN(N37280));
    INVX1 U24409 (.I(n17475), .ZN(n37281));
    NOR2X1 U24410 (.A1(n18306), .A2(N8105), .ZN(N37282));
    NANDX1 U24411 (.A1(n22194), .A2(n24767), .ZN(n37283));
    NANDX1 U24412 (.A1(N1210), .A2(n21012), .ZN(N37284));
    INVX1 U24413 (.I(n21760), .ZN(N37285));
    NANDX1 U24414 (.A1(n13657), .A2(N4022), .ZN(N37286));
    INVX1 U24415 (.I(n13877), .ZN(n37287));
    NANDX1 U24416 (.A1(n17574), .A2(n20223), .ZN(N37288));
    NOR2X1 U24417 (.A1(n21138), .A2(N578), .ZN(N37289));
    INVX1 U24418 (.I(N5692), .ZN(N37290));
    INVX1 U24419 (.I(N2633), .ZN(n37291));
    INVX1 U24420 (.I(N4506), .ZN(n37292));
    INVX1 U24421 (.I(n26390), .ZN(n37293));
    NOR2X1 U24422 (.A1(n15192), .A2(n14558), .ZN(N37294));
    NOR2X1 U24423 (.A1(N4405), .A2(N6614), .ZN(n37295));
    INVX1 U24424 (.I(N6895), .ZN(n37296));
    NOR2X1 U24425 (.A1(N11407), .A2(N4396), .ZN(N37297));
    INVX1 U24426 (.I(N8563), .ZN(n37298));
    NOR2X1 U24427 (.A1(N10726), .A2(N5618), .ZN(N37299));
    NOR2X1 U24428 (.A1(n20372), .A2(n23192), .ZN(N37300));
    NANDX1 U24429 (.A1(n27139), .A2(N2753), .ZN(n37301));
    INVX1 U24430 (.I(n18746), .ZN(N37302));
    NANDX1 U24431 (.A1(N9316), .A2(n21379), .ZN(n37303));
    NOR2X1 U24432 (.A1(N2382), .A2(n18813), .ZN(N37304));
    NANDX1 U24433 (.A1(N1483), .A2(N3868), .ZN(N37305));
    NOR2X1 U24434 (.A1(n20127), .A2(n26970), .ZN(N37306));
    NANDX1 U24435 (.A1(n21961), .A2(N3727), .ZN(N37307));
    NANDX1 U24436 (.A1(n21929), .A2(N8122), .ZN(N37308));
    NOR2X1 U24437 (.A1(N354), .A2(N3296), .ZN(N37309));
    INVX1 U24438 (.I(N5972), .ZN(N37310));
    INVX1 U24439 (.I(N10370), .ZN(N37311));
    NOR2X1 U24440 (.A1(N42), .A2(n26069), .ZN(N37312));
    NANDX1 U24441 (.A1(n18453), .A2(N3239), .ZN(N37313));
    INVX1 U24442 (.I(n16329), .ZN(n37314));
    NOR2X1 U24443 (.A1(N10559), .A2(N7271), .ZN(n37315));
    INVX1 U24444 (.I(n30026), .ZN(N37316));
    INVX1 U24445 (.I(N5720), .ZN(n37317));
    INVX1 U24446 (.I(n17440), .ZN(n37318));
    NOR2X1 U24447 (.A1(N10099), .A2(n27962), .ZN(N37319));
    NANDX1 U24448 (.A1(n24243), .A2(n19753), .ZN(N37320));
    NOR2X1 U24449 (.A1(n14954), .A2(n20106), .ZN(N37321));
    INVX1 U24450 (.I(N4951), .ZN(N37322));
    INVX1 U24451 (.I(N7163), .ZN(n37323));
    NANDX1 U24452 (.A1(N2224), .A2(N7204), .ZN(N37324));
    NANDX1 U24453 (.A1(n22700), .A2(n14218), .ZN(N37325));
    INVX1 U24454 (.I(n28741), .ZN(N37326));
    NANDX1 U24455 (.A1(n16228), .A2(N9162), .ZN(N37327));
    INVX1 U24456 (.I(n18080), .ZN(N37328));
    INVX1 U24457 (.I(N4993), .ZN(n37329));
    INVX1 U24458 (.I(n20086), .ZN(n37330));
    NANDX1 U24459 (.A1(N3474), .A2(N47), .ZN(N37331));
    INVX1 U24460 (.I(n28450), .ZN(n37332));
    NANDX1 U24461 (.A1(n28570), .A2(n19972), .ZN(n37333));
    INVX1 U24462 (.I(n18538), .ZN(N37334));
    NANDX1 U24463 (.A1(N2616), .A2(N3039), .ZN(N37335));
    NOR2X1 U24464 (.A1(n17936), .A2(N5262), .ZN(N37336));
    NOR2X1 U24465 (.A1(n17748), .A2(n16522), .ZN(n37337));
    NOR2X1 U24466 (.A1(n20798), .A2(n15125), .ZN(N37338));
    INVX1 U24467 (.I(N6888), .ZN(N37339));
    NOR2X1 U24468 (.A1(n17142), .A2(n13528), .ZN(n37340));
    NANDX1 U24469 (.A1(N10696), .A2(n14449), .ZN(N37341));
    INVX1 U24470 (.I(n21689), .ZN(N37342));
    NOR2X1 U24471 (.A1(N11891), .A2(N369), .ZN(N37343));
    NANDX1 U24472 (.A1(n24740), .A2(n28938), .ZN(n37344));
    NANDX1 U24473 (.A1(n22405), .A2(n17338), .ZN(N37345));
    NANDX1 U24474 (.A1(n13581), .A2(N8937), .ZN(N37346));
    NANDX1 U24475 (.A1(N1379), .A2(N2760), .ZN(N37347));
    NANDX1 U24476 (.A1(N7687), .A2(n19281), .ZN(N37348));
    INVX1 U24477 (.I(n17045), .ZN(N37349));
    NANDX1 U24478 (.A1(N68), .A2(N12493), .ZN(N37350));
    INVX1 U24479 (.I(N5770), .ZN(N37351));
    NANDX1 U24480 (.A1(n27572), .A2(n16465), .ZN(N37352));
    NANDX1 U24481 (.A1(N9279), .A2(N8016), .ZN(N37353));
    NOR2X1 U24482 (.A1(N9730), .A2(N8384), .ZN(N37354));
    INVX1 U24483 (.I(n23030), .ZN(N37355));
    NANDX1 U24484 (.A1(N4800), .A2(N3858), .ZN(n37356));
    NOR2X1 U24485 (.A1(n21477), .A2(n17439), .ZN(n37357));
    NOR2X1 U24486 (.A1(n29968), .A2(N7378), .ZN(N37358));
    INVX1 U24487 (.I(n26036), .ZN(N37359));
    INVX1 U24488 (.I(N2483), .ZN(N37360));
    NOR2X1 U24489 (.A1(n20670), .A2(n25449), .ZN(n37361));
    NANDX1 U24490 (.A1(N3026), .A2(N987), .ZN(n37362));
    NANDX1 U24491 (.A1(n17607), .A2(n28559), .ZN(N37363));
    NOR2X1 U24492 (.A1(n27938), .A2(n26398), .ZN(n37364));
    NANDX1 U24493 (.A1(N3176), .A2(N5991), .ZN(N37365));
    NANDX1 U24494 (.A1(n13346), .A2(n17581), .ZN(N37366));
    NOR2X1 U24495 (.A1(n18146), .A2(n21439), .ZN(n37367));
    NANDX1 U24496 (.A1(n28183), .A2(N8740), .ZN(N37368));
    NOR2X1 U24497 (.A1(n28013), .A2(n16117), .ZN(n37369));
    NOR2X1 U24498 (.A1(n23912), .A2(n19742), .ZN(n37370));
    NANDX1 U24499 (.A1(N6235), .A2(N10275), .ZN(N37371));
    INVX1 U24500 (.I(n18762), .ZN(n37372));
    NANDX1 U24501 (.A1(n22411), .A2(n25619), .ZN(N37373));
    NANDX1 U24502 (.A1(n20832), .A2(N106), .ZN(N37374));
    INVX1 U24503 (.I(n17092), .ZN(N37375));
    NOR2X1 U24504 (.A1(N9004), .A2(N11643), .ZN(N37376));
    INVX1 U24505 (.I(n22349), .ZN(N37377));
    NOR2X1 U24506 (.A1(n16219), .A2(n29055), .ZN(N37378));
    INVX1 U24507 (.I(N4493), .ZN(N37379));
    INVX1 U24508 (.I(n17825), .ZN(N37380));
    NOR2X1 U24509 (.A1(n24976), .A2(n22502), .ZN(N37381));
    NOR2X1 U24510 (.A1(N7311), .A2(N668), .ZN(N37382));
    NANDX1 U24511 (.A1(N2106), .A2(N10942), .ZN(N37383));
    NANDX1 U24512 (.A1(n20867), .A2(N1363), .ZN(n37384));
    INVX1 U24513 (.I(N4910), .ZN(n37385));
    NANDX1 U24514 (.A1(n15903), .A2(N5015), .ZN(N37386));
    NANDX1 U24515 (.A1(n21556), .A2(n25019), .ZN(N37387));
    INVX1 U24516 (.I(N3061), .ZN(N37388));
    INVX1 U24517 (.I(n16432), .ZN(N37389));
    NANDX1 U24518 (.A1(n29250), .A2(n15349), .ZN(N37390));
    NANDX1 U24519 (.A1(N3605), .A2(N12312), .ZN(N37391));
    NANDX1 U24520 (.A1(n18389), .A2(n25849), .ZN(N37392));
    NANDX1 U24521 (.A1(n15227), .A2(n21720), .ZN(N37393));
    INVX1 U24522 (.I(n19480), .ZN(N37394));
    NOR2X1 U24523 (.A1(n17410), .A2(N3581), .ZN(n37395));
    NANDX1 U24524 (.A1(n18772), .A2(n28789), .ZN(n37396));
    NANDX1 U24525 (.A1(N9463), .A2(n14555), .ZN(n37397));
    NOR2X1 U24526 (.A1(n24679), .A2(N5973), .ZN(n37398));
    NANDX1 U24527 (.A1(N64), .A2(N9033), .ZN(N37399));
    INVX1 U24528 (.I(n16495), .ZN(n37400));
    INVX1 U24529 (.I(N8625), .ZN(N37401));
    NOR2X1 U24530 (.A1(N6792), .A2(N790), .ZN(N37402));
    NANDX1 U24531 (.A1(n12970), .A2(N7739), .ZN(N37403));
    INVX1 U24532 (.I(N73), .ZN(N37404));
    NOR2X1 U24533 (.A1(N8570), .A2(N6541), .ZN(N37405));
    INVX1 U24534 (.I(N2258), .ZN(n37406));
    INVX1 U24535 (.I(N4449), .ZN(N37407));
    NOR2X1 U24536 (.A1(N1145), .A2(N3100), .ZN(N37408));
    INVX1 U24537 (.I(n29305), .ZN(N37409));
    INVX1 U24538 (.I(n14998), .ZN(N37410));
    NOR2X1 U24539 (.A1(N12187), .A2(N41), .ZN(N37411));
    INVX1 U24540 (.I(N9781), .ZN(n37412));
    INVX1 U24541 (.I(n17525), .ZN(n37413));
    NANDX1 U24542 (.A1(n25436), .A2(N7792), .ZN(N37414));
    INVX1 U24543 (.I(n14786), .ZN(N37415));
    INVX1 U24544 (.I(N6403), .ZN(n37416));
    NANDX1 U24545 (.A1(n15918), .A2(n25173), .ZN(N37417));
    INVX1 U24546 (.I(n13048), .ZN(N37418));
    INVX1 U24547 (.I(N4780), .ZN(N37419));
    NANDX1 U24548 (.A1(N2647), .A2(n27926), .ZN(N37420));
    NANDX1 U24549 (.A1(N3791), .A2(N889), .ZN(N37421));
    NOR2X1 U24550 (.A1(n21656), .A2(n25801), .ZN(n37422));
    INVX1 U24551 (.I(N3926), .ZN(n37423));
    NOR2X1 U24552 (.A1(n22056), .A2(N4956), .ZN(N37424));
    INVX1 U24553 (.I(n20169), .ZN(N37425));
    NANDX1 U24554 (.A1(N4273), .A2(N4028), .ZN(N37426));
    INVX1 U24555 (.I(n27843), .ZN(N37427));
    NANDX1 U24556 (.A1(N6324), .A2(n22807), .ZN(N37428));
    NOR2X1 U24557 (.A1(N10802), .A2(n17842), .ZN(n37429));
    INVX1 U24558 (.I(n23849), .ZN(N37430));
    NOR2X1 U24559 (.A1(n19890), .A2(n16276), .ZN(n37431));
    NOR2X1 U24560 (.A1(n17678), .A2(n14076), .ZN(N37432));
    INVX1 U24561 (.I(N7127), .ZN(N37433));
    NANDX1 U24562 (.A1(n13193), .A2(N2791), .ZN(N37434));
    NANDX1 U24563 (.A1(N5679), .A2(n29339), .ZN(N37435));
    NANDX1 U24564 (.A1(N10635), .A2(N5393), .ZN(n37436));
    NOR2X1 U24565 (.A1(N2978), .A2(n28363), .ZN(N37437));
    INVX1 U24566 (.I(N10371), .ZN(N37438));
    INVX1 U24567 (.I(N10501), .ZN(N37439));
    NOR2X1 U24568 (.A1(N7298), .A2(N10260), .ZN(N37440));
    NANDX1 U24569 (.A1(n25140), .A2(n13930), .ZN(n37441));
    INVX1 U24570 (.I(n21679), .ZN(N37442));
    NANDX1 U24571 (.A1(n26043), .A2(N9425), .ZN(N37443));
    INVX1 U24572 (.I(n28679), .ZN(N37444));
    NOR2X1 U24573 (.A1(N5608), .A2(N12376), .ZN(N37445));
    INVX1 U24574 (.I(n27096), .ZN(N37446));
    INVX1 U24575 (.I(n19833), .ZN(n37447));
    NOR2X1 U24576 (.A1(n27157), .A2(n19028), .ZN(N37448));
    NOR2X1 U24577 (.A1(n14818), .A2(N10566), .ZN(n37449));
    NOR2X1 U24578 (.A1(n25204), .A2(n20936), .ZN(N37450));
    NANDX1 U24579 (.A1(n24265), .A2(n26190), .ZN(n37451));
    INVX1 U24580 (.I(N4387), .ZN(n37452));
    INVX1 U24581 (.I(N5266), .ZN(N37453));
    NOR2X1 U24582 (.A1(n21875), .A2(n15505), .ZN(N37454));
    NANDX1 U24583 (.A1(N6341), .A2(n24930), .ZN(N37455));
    NANDX1 U24584 (.A1(N4882), .A2(n25891), .ZN(n37456));
    INVX1 U24585 (.I(N5819), .ZN(N37457));
    NANDX1 U24586 (.A1(N167), .A2(n23906), .ZN(n37458));
    NOR2X1 U24587 (.A1(n15025), .A2(n20926), .ZN(n37459));
    NANDX1 U24588 (.A1(N5137), .A2(n24304), .ZN(N37460));
    INVX1 U24589 (.I(n23612), .ZN(n37461));
    INVX1 U24590 (.I(n15815), .ZN(n37462));
    INVX1 U24591 (.I(N2059), .ZN(N37463));
    INVX1 U24592 (.I(n18143), .ZN(N37464));
    INVX1 U24593 (.I(N12536), .ZN(n37465));
    NANDX1 U24594 (.A1(N1884), .A2(N4273), .ZN(N37466));
    NOR2X1 U24595 (.A1(N1003), .A2(n29311), .ZN(N37467));
    NANDX1 U24596 (.A1(n28741), .A2(N4056), .ZN(n37468));
    INVX1 U24597 (.I(N1812), .ZN(N37469));
    NOR2X1 U24598 (.A1(N12308), .A2(n20676), .ZN(N37470));
    NOR2X1 U24599 (.A1(n19170), .A2(N5563), .ZN(n37471));
    NANDX1 U24600 (.A1(N3484), .A2(N10700), .ZN(n37472));
    INVX1 U24601 (.I(n17061), .ZN(n37473));
    NANDX1 U24602 (.A1(N3787), .A2(N2738), .ZN(n37474));
    NOR2X1 U24603 (.A1(n24543), .A2(N3166), .ZN(N37475));
    INVX1 U24604 (.I(N8110), .ZN(n37476));
    INVX1 U24605 (.I(n19286), .ZN(N37477));
    NANDX1 U24606 (.A1(N8535), .A2(N5184), .ZN(n37478));
    INVX1 U24607 (.I(n26407), .ZN(N37479));
    NANDX1 U24608 (.A1(n28297), .A2(n19023), .ZN(N37480));
    NANDX1 U24609 (.A1(n18669), .A2(n17457), .ZN(N37481));
    NANDX1 U24610 (.A1(N9207), .A2(N9659), .ZN(N37482));
    INVX1 U24611 (.I(N3331), .ZN(N37483));
    NOR2X1 U24612 (.A1(N11794), .A2(N2591), .ZN(n37484));
    NOR2X1 U24613 (.A1(n28854), .A2(n25462), .ZN(N37485));
    INVX1 U24614 (.I(n20153), .ZN(N37486));
    NOR2X1 U24615 (.A1(N12653), .A2(n23318), .ZN(n37487));
    INVX1 U24616 (.I(n20763), .ZN(N37488));
    NOR2X1 U24617 (.A1(n29799), .A2(n19316), .ZN(n37489));
    NANDX1 U24618 (.A1(n23543), .A2(n18872), .ZN(N37490));
    INVX1 U24619 (.I(n28113), .ZN(n37491));
    NOR2X1 U24620 (.A1(N9830), .A2(n27825), .ZN(N37492));
    NANDX1 U24621 (.A1(n27286), .A2(n28405), .ZN(n37493));
    NOR2X1 U24622 (.A1(N6807), .A2(n18017), .ZN(n37494));
    INVX1 U24623 (.I(n18154), .ZN(n37495));
    NOR2X1 U24624 (.A1(N5070), .A2(n13917), .ZN(N37496));
    INVX1 U24625 (.I(N394), .ZN(N37497));
    INVX1 U24626 (.I(N7103), .ZN(N37498));
    NOR2X1 U24627 (.A1(N3241), .A2(n18982), .ZN(n37499));
    NOR2X1 U24628 (.A1(n24003), .A2(n16424), .ZN(N37500));
    NOR2X1 U24629 (.A1(N1742), .A2(N10962), .ZN(N37501));
    NANDX1 U24630 (.A1(N9175), .A2(n20467), .ZN(N37502));
    INVX1 U24631 (.I(N3327), .ZN(N37503));
    NOR2X1 U24632 (.A1(n28788), .A2(n16148), .ZN(N37504));
    INVX1 U24633 (.I(n27055), .ZN(N37505));
    NANDX1 U24634 (.A1(n22812), .A2(N3495), .ZN(N37506));
    NANDX1 U24635 (.A1(n29526), .A2(n21866), .ZN(n37507));
    INVX1 U24636 (.I(N1867), .ZN(N37508));
    INVX1 U24637 (.I(N11799), .ZN(N37509));
    NANDX1 U24638 (.A1(N4480), .A2(n15388), .ZN(n37510));
    NOR2X1 U24639 (.A1(n23461), .A2(n18050), .ZN(n37511));
    NOR2X1 U24640 (.A1(n28446), .A2(n20374), .ZN(N37512));
    INVX1 U24641 (.I(n27968), .ZN(N37513));
    NANDX1 U24642 (.A1(n19173), .A2(n18298), .ZN(N37514));
    NOR2X1 U24643 (.A1(n22499), .A2(n18456), .ZN(N37515));
    NOR2X1 U24644 (.A1(n27207), .A2(N4324), .ZN(n37516));
    NANDX1 U24645 (.A1(N12366), .A2(n15696), .ZN(N37517));
    NOR2X1 U24646 (.A1(N4), .A2(n15084), .ZN(N37518));
    NOR2X1 U24647 (.A1(N11409), .A2(N5511), .ZN(N37519));
    INVX1 U24648 (.I(n23207), .ZN(N37520));
    NOR2X1 U24649 (.A1(N5532), .A2(n27155), .ZN(N37521));
    NANDX1 U24650 (.A1(n17553), .A2(n15068), .ZN(n37522));
    NOR2X1 U24651 (.A1(n15861), .A2(n24002), .ZN(N37523));
    NOR2X1 U24652 (.A1(n13692), .A2(n17225), .ZN(N37524));
    NOR2X1 U24653 (.A1(N1852), .A2(n22851), .ZN(n37525));
    INVX1 U24654 (.I(N8868), .ZN(N37526));
    NANDX1 U24655 (.A1(N9077), .A2(N1752), .ZN(N37527));
    NANDX1 U24656 (.A1(n21442), .A2(n17447), .ZN(N37528));
    INVX1 U24657 (.I(N10007), .ZN(N37529));
    NANDX1 U24658 (.A1(n21061), .A2(n21415), .ZN(n37530));
    NANDX1 U24659 (.A1(n22113), .A2(n14485), .ZN(N37531));
    INVX1 U24660 (.I(n16205), .ZN(N37532));
    NOR2X1 U24661 (.A1(N6785), .A2(N3620), .ZN(N37533));
    NOR2X1 U24662 (.A1(n27397), .A2(N8042), .ZN(N37534));
    INVX1 U24663 (.I(N9172), .ZN(N37535));
    INVX1 U24664 (.I(n14780), .ZN(N37536));
    NOR2X1 U24665 (.A1(N706), .A2(N7493), .ZN(N37537));
    NOR2X1 U24666 (.A1(N9573), .A2(n23179), .ZN(N37538));
    NANDX1 U24667 (.A1(N11325), .A2(n28619), .ZN(n37539));
    NANDX1 U24668 (.A1(n17332), .A2(n15868), .ZN(N37540));
    NANDX1 U24669 (.A1(N8286), .A2(N6792), .ZN(n37541));
    NOR2X1 U24670 (.A1(N4751), .A2(n17465), .ZN(N37542));
    INVX1 U24671 (.I(n17877), .ZN(N37543));
    NOR2X1 U24672 (.A1(n22717), .A2(n24661), .ZN(n37544));
    NOR2X1 U24673 (.A1(n26407), .A2(n21920), .ZN(N37545));
    INVX1 U24674 (.I(n23962), .ZN(N37546));
    INVX1 U24675 (.I(n21305), .ZN(N37547));
    NOR2X1 U24676 (.A1(n25590), .A2(n22010), .ZN(N37548));
    NANDX1 U24677 (.A1(n24837), .A2(n20144), .ZN(N37549));
    INVX1 U24678 (.I(n21720), .ZN(N37550));
    INVX1 U24679 (.I(n14878), .ZN(N37551));
    INVX1 U24680 (.I(N7223), .ZN(N37552));
    NANDX1 U24681 (.A1(n15361), .A2(n15509), .ZN(N37553));
    INVX1 U24682 (.I(n23531), .ZN(N37554));
    INVX1 U24683 (.I(N1985), .ZN(n37555));
    INVX1 U24684 (.I(n26696), .ZN(N37556));
    NOR2X1 U24685 (.A1(n15885), .A2(N9781), .ZN(N37557));
    NOR2X1 U24686 (.A1(N716), .A2(n20261), .ZN(N37558));
    INVX1 U24687 (.I(n24677), .ZN(N37559));
    NOR2X1 U24688 (.A1(N10666), .A2(N10402), .ZN(n37560));
    NOR2X1 U24689 (.A1(n21236), .A2(N3619), .ZN(n37561));
    NOR2X1 U24690 (.A1(N11242), .A2(n20014), .ZN(n37562));
    NOR2X1 U24691 (.A1(N1133), .A2(n23452), .ZN(N37563));
    INVX1 U24692 (.I(N8356), .ZN(N37564));
    INVX1 U24693 (.I(n19857), .ZN(N37565));
    NANDX1 U24694 (.A1(n27278), .A2(N1811), .ZN(N37566));
    NANDX1 U24695 (.A1(n29263), .A2(n25116), .ZN(n37567));
    NANDX1 U24696 (.A1(N11900), .A2(N10864), .ZN(n37568));
    INVX1 U24697 (.I(N8947), .ZN(n37569));
    NANDX1 U24698 (.A1(N6267), .A2(n17006), .ZN(n37570));
    INVX1 U24699 (.I(N4603), .ZN(N37571));
    NOR2X1 U24700 (.A1(N5080), .A2(n28528), .ZN(N37572));
    NANDX1 U24701 (.A1(N8698), .A2(N5577), .ZN(N37573));
    INVX1 U24702 (.I(n17272), .ZN(N37574));
    NANDX1 U24703 (.A1(n19704), .A2(N10587), .ZN(N37575));
    NANDX1 U24704 (.A1(n16620), .A2(n23207), .ZN(N37576));
    INVX1 U24705 (.I(n29044), .ZN(n37577));
    NOR2X1 U24706 (.A1(N7628), .A2(n20150), .ZN(N37578));
    NANDX1 U24707 (.A1(N2607), .A2(n26513), .ZN(N37579));
    INVX1 U24708 (.I(n13470), .ZN(N37580));
    NANDX1 U24709 (.A1(N6001), .A2(n13609), .ZN(N37581));
    INVX1 U24710 (.I(n23006), .ZN(N37582));
    INVX1 U24711 (.I(n23386), .ZN(N37583));
    NOR2X1 U24712 (.A1(n20625), .A2(N10338), .ZN(N37584));
    NOR2X1 U24713 (.A1(n17883), .A2(n15914), .ZN(N37585));
    NOR2X1 U24714 (.A1(N5017), .A2(N8819), .ZN(N37586));
    NOR2X1 U24715 (.A1(n15603), .A2(N6219), .ZN(n37587));
    NANDX1 U24716 (.A1(n27370), .A2(n23476), .ZN(N37588));
    NANDX1 U24717 (.A1(N6141), .A2(N966), .ZN(n37589));
    INVX1 U24718 (.I(N2734), .ZN(N37590));
    INVX1 U24719 (.I(N3603), .ZN(N37591));
    NOR2X1 U24720 (.A1(N5602), .A2(N4681), .ZN(N37592));
    NOR2X1 U24721 (.A1(N7771), .A2(N12026), .ZN(N37593));
    NOR2X1 U24722 (.A1(N4618), .A2(N5274), .ZN(n37594));
    NOR2X1 U24723 (.A1(n25242), .A2(n15611), .ZN(N37595));
    NANDX1 U24724 (.A1(n12987), .A2(n20085), .ZN(N37596));
    INVX1 U24725 (.I(N6565), .ZN(n37597));
    INVX1 U24726 (.I(N600), .ZN(N37598));
    NOR2X1 U24727 (.A1(N4985), .A2(N210), .ZN(n37599));
    NANDX1 U24728 (.A1(n17021), .A2(n28864), .ZN(N37600));
    NANDX1 U24729 (.A1(N6547), .A2(n24652), .ZN(N37601));
    INVX1 U24730 (.I(N10119), .ZN(N37602));
    NOR2X1 U24731 (.A1(N12442), .A2(N4281), .ZN(N37603));
    NOR2X1 U24732 (.A1(N6791), .A2(N613), .ZN(N37604));
    INVX1 U24733 (.I(n24145), .ZN(N37605));
    NOR2X1 U24734 (.A1(n27355), .A2(N9023), .ZN(n37606));
    NANDX1 U24735 (.A1(N1389), .A2(N10330), .ZN(N37607));
    INVX1 U24736 (.I(n21474), .ZN(N37608));
    NOR2X1 U24737 (.A1(n27144), .A2(N8800), .ZN(N37609));
    NANDX1 U24738 (.A1(n26433), .A2(n13784), .ZN(N37610));
    INVX1 U24739 (.I(n22954), .ZN(N37611));
    INVX1 U24740 (.I(N4596), .ZN(N37612));
    NANDX1 U24741 (.A1(n25912), .A2(n29247), .ZN(N37613));
    NANDX1 U24742 (.A1(n24591), .A2(n15924), .ZN(N37614));
    INVX1 U24743 (.I(n17432), .ZN(n37615));
    NANDX1 U24744 (.A1(n15923), .A2(n18044), .ZN(N37616));
    NOR2X1 U24745 (.A1(n28629), .A2(N11835), .ZN(N37617));
    INVX1 U24746 (.I(N7514), .ZN(N37618));
    NANDX1 U24747 (.A1(n27968), .A2(n17844), .ZN(n37619));
    NOR2X1 U24748 (.A1(N7865), .A2(N4206), .ZN(N37620));
    INVX1 U24749 (.I(n16664), .ZN(N37621));
    NANDX1 U24750 (.A1(n21870), .A2(n19009), .ZN(N37622));
    INVX1 U24751 (.I(n14686), .ZN(N37623));
    INVX1 U24752 (.I(N1633), .ZN(N37624));
    NOR2X1 U24753 (.A1(N4010), .A2(N743), .ZN(N37625));
    NANDX1 U24754 (.A1(n28600), .A2(N5227), .ZN(n37626));
    NOR2X1 U24755 (.A1(N4456), .A2(N1069), .ZN(n37627));
    INVX1 U24756 (.I(n22499), .ZN(N37628));
    NOR2X1 U24757 (.A1(N7522), .A2(N4196), .ZN(N37629));
    INVX1 U24758 (.I(n15036), .ZN(N37630));
    NANDX1 U24759 (.A1(N1824), .A2(n21440), .ZN(N37631));
    NOR2X1 U24760 (.A1(N9688), .A2(n14206), .ZN(N37632));
    NOR2X1 U24761 (.A1(n26352), .A2(N5374), .ZN(N37633));
    NOR2X1 U24762 (.A1(N3784), .A2(n21109), .ZN(n37634));
    INVX1 U24763 (.I(N12019), .ZN(N37635));
    INVX1 U24764 (.I(N3933), .ZN(N37636));
    NANDX1 U24765 (.A1(N12044), .A2(n29484), .ZN(n37637));
    INVX1 U24766 (.I(n17271), .ZN(N37638));
    INVX1 U24767 (.I(n26205), .ZN(N37639));
    INVX1 U24768 (.I(N1486), .ZN(n37640));
    NOR2X1 U24769 (.A1(N7193), .A2(N9007), .ZN(n37641));
    NOR2X1 U24770 (.A1(n22626), .A2(N12603), .ZN(n37642));
    NOR2X1 U24771 (.A1(n13010), .A2(N3905), .ZN(N37643));
    NANDX1 U24772 (.A1(n22698), .A2(n18111), .ZN(N37644));
    NANDX1 U24773 (.A1(N7473), .A2(N12045), .ZN(N37645));
    INVX1 U24774 (.I(N11256), .ZN(N37646));
    NANDX1 U24775 (.A1(N2689), .A2(n23274), .ZN(N37647));
    NOR2X1 U24776 (.A1(N6621), .A2(n16424), .ZN(N37648));
    NOR2X1 U24777 (.A1(n24665), .A2(N8037), .ZN(N37649));
    INVX1 U24778 (.I(n17120), .ZN(N37650));
    INVX1 U24779 (.I(n27652), .ZN(N37651));
    NOR2X1 U24780 (.A1(n22670), .A2(N4708), .ZN(n37652));
    NOR2X1 U24781 (.A1(N3856), .A2(n15894), .ZN(n37653));
    INVX1 U24782 (.I(N8664), .ZN(N37654));
    INVX1 U24783 (.I(n21240), .ZN(N37655));
    NANDX1 U24784 (.A1(N10024), .A2(n27911), .ZN(N37656));
    INVX1 U24785 (.I(N6057), .ZN(n37657));
    NOR2X1 U24786 (.A1(n14002), .A2(n17312), .ZN(N37658));
    NANDX1 U24787 (.A1(n16690), .A2(n29147), .ZN(N37659));
    NANDX1 U24788 (.A1(N11871), .A2(n15433), .ZN(N37660));
    NANDX1 U24789 (.A1(n25096), .A2(n23469), .ZN(N37661));
    NOR2X1 U24790 (.A1(N639), .A2(n16134), .ZN(n37662));
    INVX1 U24791 (.I(N7804), .ZN(N37663));
    NANDX1 U24792 (.A1(N590), .A2(N12537), .ZN(N37664));
    NOR2X1 U24793 (.A1(n16483), .A2(n29872), .ZN(n37665));
    NOR2X1 U24794 (.A1(N3810), .A2(N9535), .ZN(N37666));
    INVX1 U24795 (.I(N2394), .ZN(n37667));
    INVX1 U24796 (.I(N1517), .ZN(N37668));
    NOR2X1 U24797 (.A1(n24385), .A2(N4079), .ZN(n37669));
    NOR2X1 U24798 (.A1(n14340), .A2(N9329), .ZN(N37670));
    NOR2X1 U24799 (.A1(n18611), .A2(n21199), .ZN(N37671));
    NOR2X1 U24800 (.A1(n26364), .A2(N4719), .ZN(N37672));
    INVX1 U24801 (.I(N6034), .ZN(N37673));
    NANDX1 U24802 (.A1(n15351), .A2(n13355), .ZN(N37674));
    INVX1 U24803 (.I(N12578), .ZN(n37675));
    NANDX1 U24804 (.A1(n14258), .A2(n13659), .ZN(n37676));
    INVX1 U24805 (.I(n13992), .ZN(N37677));
    NANDX1 U24806 (.A1(N11358), .A2(n23526), .ZN(N37678));
    NOR2X1 U24807 (.A1(n13752), .A2(n19395), .ZN(n37679));
    NANDX1 U24808 (.A1(N10763), .A2(n13643), .ZN(N37680));
    NANDX1 U24809 (.A1(n25085), .A2(n16543), .ZN(n37681));
    INVX1 U24810 (.I(n26978), .ZN(n37682));
    INVX1 U24811 (.I(N2944), .ZN(n37683));
    NOR2X1 U24812 (.A1(n19940), .A2(N7662), .ZN(N37684));
    INVX1 U24813 (.I(n25973), .ZN(n37685));
    NANDX1 U24814 (.A1(n17295), .A2(N9190), .ZN(n37686));
    NANDX1 U24815 (.A1(n29872), .A2(N11695), .ZN(N37687));
    NOR2X1 U24816 (.A1(N1954), .A2(n19244), .ZN(N37688));
    NOR2X1 U24817 (.A1(n25357), .A2(N464), .ZN(n37689));
    NANDX1 U24818 (.A1(N3618), .A2(N2776), .ZN(N37690));
    NANDX1 U24819 (.A1(n13532), .A2(N2099), .ZN(N37691));
    NOR2X1 U24820 (.A1(n27524), .A2(n27184), .ZN(N37692));
    NOR2X1 U24821 (.A1(n20708), .A2(N12585), .ZN(N37693));
    INVX1 U24822 (.I(n23652), .ZN(n37694));
    NANDX1 U24823 (.A1(N4879), .A2(n19874), .ZN(N37695));
    NANDX1 U24824 (.A1(N714), .A2(n21453), .ZN(N37696));
    NOR2X1 U24825 (.A1(n28601), .A2(n24753), .ZN(N37697));
    NOR2X1 U24826 (.A1(n28857), .A2(N12173), .ZN(n37698));
    NANDX1 U24827 (.A1(n17963), .A2(N2145), .ZN(n37699));
    NANDX1 U24828 (.A1(N6987), .A2(N4204), .ZN(n37700));
    NANDX1 U24829 (.A1(n28461), .A2(n25657), .ZN(N37701));
    NANDX1 U24830 (.A1(N422), .A2(N478), .ZN(n37702));
    NOR2X1 U24831 (.A1(n16166), .A2(N10539), .ZN(n37703));
    INVX1 U24832 (.I(n28750), .ZN(n37704));
    INVX1 U24833 (.I(n21714), .ZN(N37705));
    NOR2X1 U24834 (.A1(n19054), .A2(N11451), .ZN(n37706));
    NANDX1 U24835 (.A1(n19767), .A2(N2766), .ZN(N37707));
    NANDX1 U24836 (.A1(N6791), .A2(n16080), .ZN(N37708));
    NANDX1 U24837 (.A1(n24208), .A2(n16813), .ZN(N37709));
    NOR2X1 U24838 (.A1(N12033), .A2(N7519), .ZN(N37710));
    NANDX1 U24839 (.A1(n19020), .A2(N11722), .ZN(N37711));
    INVX1 U24840 (.I(n17343), .ZN(N37712));
    NANDX1 U24841 (.A1(n15330), .A2(N6325), .ZN(N37713));
    NANDX1 U24842 (.A1(N4124), .A2(n22491), .ZN(N37714));
    NOR2X1 U24843 (.A1(n13626), .A2(N9664), .ZN(N37715));
    NOR2X1 U24844 (.A1(N5202), .A2(N12148), .ZN(N37716));
    INVX1 U24845 (.I(N5213), .ZN(N37717));
    NOR2X1 U24846 (.A1(n29674), .A2(n26677), .ZN(n37718));
    INVX1 U24847 (.I(n25025), .ZN(n37719));
    NOR2X1 U24848 (.A1(n22949), .A2(n19096), .ZN(N37720));
    INVX1 U24849 (.I(n18842), .ZN(n37721));
    NOR2X1 U24850 (.A1(n25510), .A2(n19132), .ZN(n37722));
    NOR2X1 U24851 (.A1(N7094), .A2(N1478), .ZN(N37723));
    INVX1 U24852 (.I(N2895), .ZN(N37724));
    INVX1 U24853 (.I(N9360), .ZN(n37725));
    NOR2X1 U24854 (.A1(n28190), .A2(N1713), .ZN(N37726));
    NANDX1 U24855 (.A1(N11678), .A2(n30074), .ZN(N37727));
    NANDX1 U24856 (.A1(N5440), .A2(N12084), .ZN(N37728));
    NANDX1 U24857 (.A1(n29351), .A2(n21090), .ZN(N37729));
    NOR2X1 U24858 (.A1(n25890), .A2(N12668), .ZN(N37730));
    INVX1 U24859 (.I(n27069), .ZN(N37731));
    INVX1 U24860 (.I(n27528), .ZN(n37732));
    NOR2X1 U24861 (.A1(n12882), .A2(n17079), .ZN(n37733));
    NOR2X1 U24862 (.A1(N1876), .A2(n14211), .ZN(N37734));
    INVX1 U24863 (.I(n22051), .ZN(n37735));
    INVX1 U24864 (.I(N8845), .ZN(N37736));
    NANDX1 U24865 (.A1(n15165), .A2(N8017), .ZN(N37737));
    NANDX1 U24866 (.A1(N5438), .A2(n14006), .ZN(N37738));
    NANDX1 U24867 (.A1(N5375), .A2(N10848), .ZN(N37739));
    NOR2X1 U24868 (.A1(N6019), .A2(n17598), .ZN(N37740));
    INVX1 U24869 (.I(n27109), .ZN(n37741));
    INVX1 U24870 (.I(n21933), .ZN(N37742));
    NOR2X1 U24871 (.A1(n20876), .A2(N7425), .ZN(N37743));
    INVX1 U24872 (.I(n18266), .ZN(n37744));
    NOR2X1 U24873 (.A1(N5120), .A2(N5208), .ZN(N37745));
    NANDX1 U24874 (.A1(n25693), .A2(N7979), .ZN(N37746));
    NOR2X1 U24875 (.A1(N6167), .A2(n13784), .ZN(N37747));
    NANDX1 U24876 (.A1(N10707), .A2(n28949), .ZN(N37748));
    NOR2X1 U24877 (.A1(n24737), .A2(N4249), .ZN(N37749));
    NOR2X1 U24878 (.A1(n27567), .A2(n28321), .ZN(N37750));
    NANDX1 U24879 (.A1(n24397), .A2(N4203), .ZN(N37751));
    NANDX1 U24880 (.A1(n20440), .A2(N1174), .ZN(N37752));
    NOR2X1 U24881 (.A1(N796), .A2(n29510), .ZN(N37753));
    NANDX1 U24882 (.A1(N8220), .A2(n21748), .ZN(N37754));
    NANDX1 U24883 (.A1(N7688), .A2(n26868), .ZN(n37755));
    NOR2X1 U24884 (.A1(n17452), .A2(N10984), .ZN(N37756));
    INVX1 U24885 (.I(n21726), .ZN(N37757));
    NANDX1 U24886 (.A1(N1791), .A2(N4707), .ZN(n37758));
    NOR2X1 U24887 (.A1(N602), .A2(n14402), .ZN(N37759));
    NOR2X1 U24888 (.A1(n23548), .A2(n26664), .ZN(n37760));
    NOR2X1 U24889 (.A1(n21732), .A2(N8197), .ZN(N37761));
    NOR2X1 U24890 (.A1(n25934), .A2(n26025), .ZN(n37762));
    NOR2X1 U24891 (.A1(n15668), .A2(n14720), .ZN(N37763));
    NANDX1 U24892 (.A1(n15040), .A2(n24291), .ZN(N37764));
    INVX1 U24893 (.I(n25348), .ZN(n37765));
    NANDX1 U24894 (.A1(n24227), .A2(n22078), .ZN(N37766));
    NANDX1 U24895 (.A1(N11541), .A2(n21623), .ZN(n37767));
    INVX1 U24896 (.I(N3129), .ZN(N37768));
    NOR2X1 U24897 (.A1(n21953), .A2(n26533), .ZN(N37769));
    NOR2X1 U24898 (.A1(N11115), .A2(n29495), .ZN(N37770));
    NOR2X1 U24899 (.A1(N4525), .A2(n14582), .ZN(n37771));
    NOR2X1 U24900 (.A1(n14817), .A2(n22778), .ZN(N37772));
    NOR2X1 U24901 (.A1(n29311), .A2(N7226), .ZN(N37773));
    NOR2X1 U24902 (.A1(n14841), .A2(N10507), .ZN(N37774));
    INVX1 U24903 (.I(n18441), .ZN(N37775));
    INVX1 U24904 (.I(N3709), .ZN(N37776));
    NANDX1 U24905 (.A1(n15211), .A2(n16496), .ZN(N37777));
    NOR2X1 U24906 (.A1(N5791), .A2(n28036), .ZN(N37778));
    NANDX1 U24907 (.A1(n25953), .A2(n19725), .ZN(N37779));
    INVX1 U24908 (.I(n17768), .ZN(N37780));
    INVX1 U24909 (.I(n26584), .ZN(N37781));
    NANDX1 U24910 (.A1(N4038), .A2(n21077), .ZN(N37782));
    NOR2X1 U24911 (.A1(n18620), .A2(N1137), .ZN(N37783));
    INVX1 U24912 (.I(n29958), .ZN(n37784));
    NOR2X1 U24913 (.A1(n24518), .A2(n25745), .ZN(n37785));
    NANDX1 U24914 (.A1(N9222), .A2(N6114), .ZN(N37786));
    INVX1 U24915 (.I(n16223), .ZN(n37787));
    NOR2X1 U24916 (.A1(n21162), .A2(n18435), .ZN(N37788));
    INVX1 U24917 (.I(N7520), .ZN(N37789));
    NOR2X1 U24918 (.A1(N8896), .A2(n24116), .ZN(N37790));
    INVX1 U24919 (.I(n23409), .ZN(N37791));
    NOR2X1 U24920 (.A1(N7016), .A2(n29737), .ZN(N37792));
    NOR2X1 U24921 (.A1(N3462), .A2(n28481), .ZN(N37793));
    NOR2X1 U24922 (.A1(n13099), .A2(N8871), .ZN(n37794));
    NOR2X1 U24923 (.A1(N2796), .A2(N4078), .ZN(N37795));
    NOR2X1 U24924 (.A1(n24093), .A2(n28596), .ZN(N37796));
    INVX1 U24925 (.I(N12800), .ZN(N37797));
    NOR2X1 U24926 (.A1(N8263), .A2(N116), .ZN(N37798));
    NANDX1 U24927 (.A1(n26294), .A2(N9838), .ZN(n37799));
    NANDX1 U24928 (.A1(n17960), .A2(N5918), .ZN(n37800));
    INVX1 U24929 (.I(n15416), .ZN(n37801));
    INVX1 U24930 (.I(n26090), .ZN(n37802));
    NANDX1 U24931 (.A1(N9418), .A2(N2968), .ZN(N37803));
    NANDX1 U24932 (.A1(n16361), .A2(n25128), .ZN(N37804));
    INVX1 U24933 (.I(n15903), .ZN(n37805));
    NANDX1 U24934 (.A1(N4061), .A2(n22624), .ZN(N37806));
    INVX1 U24935 (.I(n26836), .ZN(N37807));
    NOR2X1 U24936 (.A1(n23538), .A2(n25294), .ZN(N37808));
    NOR2X1 U24937 (.A1(n24898), .A2(n21534), .ZN(N37809));
    NANDX1 U24938 (.A1(n25014), .A2(n22558), .ZN(n37810));
    NANDX1 U24939 (.A1(n23412), .A2(N440), .ZN(N37811));
    INVX1 U24940 (.I(n17891), .ZN(n37812));
    NANDX1 U24941 (.A1(n16094), .A2(N6347), .ZN(N37813));
    NOR2X1 U24942 (.A1(n13341), .A2(n15765), .ZN(N37814));
    NOR2X1 U24943 (.A1(n21627), .A2(n20686), .ZN(n37815));
    INVX1 U24944 (.I(N5377), .ZN(N37816));
    INVX1 U24945 (.I(n18864), .ZN(n37817));
    NOR2X1 U24946 (.A1(n17636), .A2(n18309), .ZN(n37818));
    NOR2X1 U24947 (.A1(N5225), .A2(N270), .ZN(N37819));
    INVX1 U24948 (.I(N6403), .ZN(N37820));
    INVX1 U24949 (.I(n18646), .ZN(n37821));
    NOR2X1 U24950 (.A1(N8605), .A2(N11066), .ZN(n37822));
    INVX1 U24951 (.I(N1879), .ZN(n37823));
    NOR2X1 U24952 (.A1(n25195), .A2(n19769), .ZN(n37824));
    INVX1 U24953 (.I(N11151), .ZN(n37825));
    NOR2X1 U24954 (.A1(n26669), .A2(n13052), .ZN(N37826));
    INVX1 U24955 (.I(n23756), .ZN(N37827));
    INVX1 U24956 (.I(N9550), .ZN(N37828));
    NOR2X1 U24957 (.A1(n28616), .A2(N4562), .ZN(n37829));
    NOR2X1 U24958 (.A1(n26613), .A2(N10758), .ZN(N37830));
    NANDX1 U24959 (.A1(n21309), .A2(n15982), .ZN(N37831));
    NOR2X1 U24960 (.A1(n29860), .A2(N10945), .ZN(N37832));
    NOR2X1 U24961 (.A1(n18368), .A2(N3909), .ZN(N37833));
    INVX1 U24962 (.I(n17994), .ZN(n37834));
    NANDX1 U24963 (.A1(n24470), .A2(n18059), .ZN(n37835));
    INVX1 U24964 (.I(N2663), .ZN(n37836));
    NOR2X1 U24965 (.A1(n23193), .A2(N5900), .ZN(N37837));
    NOR2X1 U24966 (.A1(N6108), .A2(n24901), .ZN(N37838));
    NOR2X1 U24967 (.A1(n29346), .A2(N4313), .ZN(n37839));
    NOR2X1 U24968 (.A1(n27824), .A2(n27572), .ZN(N37840));
    NOR2X1 U24969 (.A1(N12861), .A2(n26890), .ZN(N37841));
    NANDX1 U24970 (.A1(N4032), .A2(N12735), .ZN(n37842));
    INVX1 U24971 (.I(n22452), .ZN(n37843));
    INVX1 U24972 (.I(N6751), .ZN(N37844));
    INVX1 U24973 (.I(N4709), .ZN(n37845));
    NANDX1 U24974 (.A1(N5797), .A2(N2997), .ZN(N37846));
    NOR2X1 U24975 (.A1(N12416), .A2(n15039), .ZN(N37847));
    NOR2X1 U24976 (.A1(n28706), .A2(n26793), .ZN(n37848));
    NOR2X1 U24977 (.A1(N11391), .A2(N2763), .ZN(n37849));
    INVX1 U24978 (.I(n17831), .ZN(n37850));
    NOR2X1 U24979 (.A1(N8433), .A2(n17225), .ZN(N37851));
    INVX1 U24980 (.I(n24565), .ZN(N37852));
    NANDX1 U24981 (.A1(n19777), .A2(n21318), .ZN(N37853));
    NOR2X1 U24982 (.A1(N12369), .A2(N3915), .ZN(N37854));
    NOR2X1 U24983 (.A1(n23382), .A2(N4715), .ZN(N37855));
    INVX1 U24984 (.I(n22624), .ZN(n37856));
    INVX1 U24985 (.I(n19659), .ZN(N37857));
    NANDX1 U24986 (.A1(N981), .A2(N1756), .ZN(N37858));
    INVX1 U24987 (.I(n16019), .ZN(N37859));
    NANDX1 U24988 (.A1(n27966), .A2(N12674), .ZN(N37860));
    NANDX1 U24989 (.A1(n27917), .A2(N3997), .ZN(N37861));
    NOR2X1 U24990 (.A1(n15610), .A2(n13227), .ZN(N37862));
    INVX1 U24991 (.I(N2697), .ZN(N37863));
    NANDX1 U24992 (.A1(N10110), .A2(N12436), .ZN(N37864));
    INVX1 U24993 (.I(N1290), .ZN(N37865));
    NOR2X1 U24994 (.A1(N10711), .A2(n23902), .ZN(N37866));
    NOR2X1 U24995 (.A1(N3955), .A2(n28617), .ZN(N37867));
    INVX1 U24996 (.I(n15140), .ZN(N37868));
    INVX1 U24997 (.I(n26919), .ZN(N37869));
    INVX1 U24998 (.I(n27581), .ZN(n37870));
    INVX1 U24999 (.I(n19941), .ZN(N37871));
    NANDX1 U25000 (.A1(n22449), .A2(N6330), .ZN(N37872));
    NOR2X1 U25001 (.A1(N6881), .A2(N4109), .ZN(n37873));
    INVX1 U25002 (.I(n25570), .ZN(N37874));
    NANDX1 U25003 (.A1(N9041), .A2(N11115), .ZN(N37875));
    NANDX1 U25004 (.A1(n17744), .A2(n21225), .ZN(N37876));
    NOR2X1 U25005 (.A1(n16086), .A2(n22514), .ZN(N37877));
    INVX1 U25006 (.I(n15358), .ZN(N37878));
    NOR2X1 U25007 (.A1(N2018), .A2(n19312), .ZN(N37879));
    NOR2X1 U25008 (.A1(N9279), .A2(n23012), .ZN(n37880));
    INVX1 U25009 (.I(n24758), .ZN(n37881));
    INVX1 U25010 (.I(n27362), .ZN(N37882));
    INVX1 U25011 (.I(N3360), .ZN(n37883));
    NANDX1 U25012 (.A1(N4167), .A2(n28387), .ZN(N37884));
    NANDX1 U25013 (.A1(N11048), .A2(N2359), .ZN(N37885));
    NOR2X1 U25014 (.A1(n25178), .A2(n29335), .ZN(n37886));
    NOR2X1 U25015 (.A1(N6156), .A2(n28871), .ZN(N37887));
    NANDX1 U25016 (.A1(n15941), .A2(N10706), .ZN(N37888));
    NOR2X1 U25017 (.A1(n27015), .A2(n14478), .ZN(N37889));
    NOR2X1 U25018 (.A1(N1717), .A2(n16495), .ZN(N37890));
    INVX1 U25019 (.I(N5035), .ZN(N37891));
    NANDX1 U25020 (.A1(n27155), .A2(n23514), .ZN(N37892));
    NOR2X1 U25021 (.A1(N10574), .A2(N9299), .ZN(N37893));
    NOR2X1 U25022 (.A1(N2494), .A2(N8546), .ZN(N37894));
    NOR2X1 U25023 (.A1(N743), .A2(N11049), .ZN(N37895));
    NANDX1 U25024 (.A1(n21799), .A2(N9367), .ZN(N37896));
    NANDX1 U25025 (.A1(n20997), .A2(n16726), .ZN(n37897));
    NOR2X1 U25026 (.A1(n19730), .A2(N11691), .ZN(N37898));
    NOR2X1 U25027 (.A1(n18996), .A2(N11302), .ZN(n37899));
    NANDX1 U25028 (.A1(N3336), .A2(n26271), .ZN(N37900));
    INVX1 U25029 (.I(N8392), .ZN(n37901));
    NANDX1 U25030 (.A1(n29730), .A2(N11286), .ZN(n37902));
    NOR2X1 U25031 (.A1(n23106), .A2(n20240), .ZN(N37903));
    NANDX1 U25032 (.A1(N2268), .A2(n29611), .ZN(N37904));
    NOR2X1 U25033 (.A1(n29511), .A2(n13011), .ZN(N37905));
    INVX1 U25034 (.I(N10422), .ZN(n37906));
    INVX1 U25035 (.I(n28721), .ZN(N37907));
    NANDX1 U25036 (.A1(N4204), .A2(n19580), .ZN(N37908));
    INVX1 U25037 (.I(n25804), .ZN(N37909));
    INVX1 U25038 (.I(n25326), .ZN(n37910));
    NANDX1 U25039 (.A1(n16729), .A2(n25188), .ZN(N37911));
    INVX1 U25040 (.I(N8626), .ZN(N37912));
    INVX1 U25041 (.I(n13346), .ZN(N37913));
    NOR2X1 U25042 (.A1(n28856), .A2(N1499), .ZN(N37914));
    NOR2X1 U25043 (.A1(n21970), .A2(n24604), .ZN(N37915));
    NOR2X1 U25044 (.A1(n25656), .A2(n15432), .ZN(n37916));
    NOR2X1 U25045 (.A1(N1699), .A2(N3366), .ZN(N37917));
    NOR2X1 U25046 (.A1(N8621), .A2(N2349), .ZN(N37918));
    NOR2X1 U25047 (.A1(n25902), .A2(N10698), .ZN(N37919));
    NANDX1 U25048 (.A1(N3906), .A2(n24333), .ZN(N37920));
    INVX1 U25049 (.I(N1639), .ZN(N37921));
    NOR2X1 U25050 (.A1(n25664), .A2(N6928), .ZN(N37922));
    NOR2X1 U25051 (.A1(N2875), .A2(n15553), .ZN(N37923));
    NANDX1 U25052 (.A1(n16220), .A2(n21130), .ZN(N37924));
    INVX1 U25053 (.I(n17718), .ZN(n37925));
    NOR2X1 U25054 (.A1(N10823), .A2(N746), .ZN(n37926));
    NOR2X1 U25055 (.A1(N6342), .A2(N4738), .ZN(N37927));
    NOR2X1 U25056 (.A1(n26738), .A2(N8104), .ZN(N37928));
    NANDX1 U25057 (.A1(N5221), .A2(N10452), .ZN(N37929));
    INVX1 U25058 (.I(n19683), .ZN(N37930));
    INVX1 U25059 (.I(N7208), .ZN(n37931));
    INVX1 U25060 (.I(N3905), .ZN(N37932));
    NOR2X1 U25061 (.A1(n25226), .A2(N11986), .ZN(N37933));
    INVX1 U25062 (.I(n20715), .ZN(N37934));
    INVX1 U25063 (.I(n16764), .ZN(N37935));
    INVX1 U25064 (.I(n16691), .ZN(n37936));
    INVX1 U25065 (.I(n15821), .ZN(N37937));
    NOR2X1 U25066 (.A1(n27823), .A2(N12237), .ZN(N37938));
    NOR2X1 U25067 (.A1(n17129), .A2(n15618), .ZN(N37939));
    NANDX1 U25068 (.A1(n21867), .A2(N2559), .ZN(N37940));
    NANDX1 U25069 (.A1(n18531), .A2(N8948), .ZN(N37941));
    NOR2X1 U25070 (.A1(n17543), .A2(N7925), .ZN(n37942));
    NOR2X1 U25071 (.A1(n27252), .A2(n15132), .ZN(N37943));
    INVX1 U25072 (.I(n19717), .ZN(N37944));
    INVX1 U25073 (.I(n28570), .ZN(N37945));
    INVX1 U25074 (.I(N5808), .ZN(N37946));
    NOR2X1 U25075 (.A1(N5242), .A2(n22572), .ZN(n37947));
    INVX1 U25076 (.I(N10494), .ZN(N37948));
    INVX1 U25077 (.I(n18218), .ZN(N37949));
    NANDX1 U25078 (.A1(N225), .A2(N317), .ZN(N37950));
    INVX1 U25079 (.I(n17354), .ZN(n37951));
    NANDX1 U25080 (.A1(N9356), .A2(n27781), .ZN(N37952));
    NANDX1 U25081 (.A1(N5785), .A2(n16174), .ZN(N37953));
    INVX1 U25082 (.I(n26133), .ZN(n37954));
    NOR2X1 U25083 (.A1(N12485), .A2(N5889), .ZN(n37955));
    INVX1 U25084 (.I(n16178), .ZN(n37956));
    NANDX1 U25085 (.A1(n27668), .A2(N8096), .ZN(N37957));
    NANDX1 U25086 (.A1(n29232), .A2(n13904), .ZN(n37958));
    NANDX1 U25087 (.A1(n23034), .A2(n25036), .ZN(N37959));
    NOR2X1 U25088 (.A1(N3390), .A2(n27575), .ZN(N37960));
    NOR2X1 U25089 (.A1(n26686), .A2(n27799), .ZN(N37961));
    INVX1 U25090 (.I(n24773), .ZN(n37962));
    INVX1 U25091 (.I(n17919), .ZN(n37963));
    INVX1 U25092 (.I(N1219), .ZN(N37964));
    NANDX1 U25093 (.A1(n17034), .A2(n17392), .ZN(N37965));
    NOR2X1 U25094 (.A1(n13029), .A2(n28229), .ZN(N37966));
    NOR2X1 U25095 (.A1(N7478), .A2(N6043), .ZN(N37967));
    INVX1 U25096 (.I(n16710), .ZN(N37968));
    NOR2X1 U25097 (.A1(n13274), .A2(N1495), .ZN(N37969));
    NOR2X1 U25098 (.A1(n27177), .A2(N5427), .ZN(N37970));
    NANDX1 U25099 (.A1(n22075), .A2(N11756), .ZN(N37971));
    NANDX1 U25100 (.A1(n19512), .A2(N6165), .ZN(N37972));
    NANDX1 U25101 (.A1(N5735), .A2(n19589), .ZN(N37973));
    NANDX1 U25102 (.A1(N9310), .A2(N7371), .ZN(n37974));
    NANDX1 U25103 (.A1(N10529), .A2(n20903), .ZN(n37975));
    NOR2X1 U25104 (.A1(n27920), .A2(N8858), .ZN(n37976));
    INVX1 U25105 (.I(n26012), .ZN(N37977));
    NOR2X1 U25106 (.A1(N4608), .A2(n20615), .ZN(n37978));
    INVX1 U25107 (.I(N9878), .ZN(N37979));
    NANDX1 U25108 (.A1(n16311), .A2(N11373), .ZN(N37980));
    INVX1 U25109 (.I(n13350), .ZN(N37981));
    NANDX1 U25110 (.A1(n18237), .A2(n23986), .ZN(N37982));
    NOR2X1 U25111 (.A1(n13010), .A2(N1921), .ZN(N37983));
    INVX1 U25112 (.I(N4331), .ZN(n37984));
    NOR2X1 U25113 (.A1(N1292), .A2(N8985), .ZN(n37985));
    NOR2X1 U25114 (.A1(N8662), .A2(N6190), .ZN(N37986));
    NANDX1 U25115 (.A1(n18125), .A2(n20428), .ZN(N37987));
    NANDX1 U25116 (.A1(n26982), .A2(n17558), .ZN(N37988));
    NOR2X1 U25117 (.A1(n24841), .A2(N10727), .ZN(N37989));
    NANDX1 U25118 (.A1(n27877), .A2(N9165), .ZN(N37990));
    INVX1 U25119 (.I(n14050), .ZN(n37991));
    NANDX1 U25120 (.A1(N5472), .A2(n15961), .ZN(n37992));
    NOR2X1 U25121 (.A1(n23709), .A2(n28507), .ZN(n37993));
    NOR2X1 U25122 (.A1(n25279), .A2(N290), .ZN(N37994));
    INVX1 U25123 (.I(n18170), .ZN(n37995));
    NOR2X1 U25124 (.A1(n21824), .A2(n27154), .ZN(n37996));
    NANDX1 U25125 (.A1(N348), .A2(N3206), .ZN(n37997));
    INVX1 U25126 (.I(n18472), .ZN(N37998));
    INVX1 U25127 (.I(N1782), .ZN(N37999));
    NOR2X1 U25128 (.A1(n29752), .A2(N53), .ZN(N38000));
    NOR2X1 U25129 (.A1(n29039), .A2(N7499), .ZN(n38001));
    NANDX1 U25130 (.A1(N8066), .A2(N8995), .ZN(n38002));
    INVX1 U25131 (.I(N5725), .ZN(N38003));
    INVX1 U25132 (.I(N3451), .ZN(n38004));
    INVX1 U25133 (.I(n26735), .ZN(N38005));
    INVX1 U25134 (.I(n28874), .ZN(N38006));
    INVX1 U25135 (.I(N9369), .ZN(n38007));
    NANDX1 U25136 (.A1(n28606), .A2(N5874), .ZN(n38008));
    NANDX1 U25137 (.A1(n14183), .A2(N7904), .ZN(N38009));
    NOR2X1 U25138 (.A1(N5949), .A2(n25987), .ZN(N38010));
    NANDX1 U25139 (.A1(n18143), .A2(n27768), .ZN(N38011));
    INVX1 U25140 (.I(n17757), .ZN(N38012));
    NANDX1 U25141 (.A1(n28049), .A2(N5219), .ZN(n38013));
    NOR2X1 U25142 (.A1(N1490), .A2(N1845), .ZN(n38014));
    NANDX1 U25143 (.A1(n19117), .A2(N7569), .ZN(N38015));
    NOR2X1 U25144 (.A1(N11129), .A2(n16311), .ZN(N38016));
    NANDX1 U25145 (.A1(N1509), .A2(N3608), .ZN(N38017));
    INVX1 U25146 (.I(N10877), .ZN(n38018));
    NOR2X1 U25147 (.A1(N7085), .A2(N5311), .ZN(N38019));
    NANDX1 U25148 (.A1(N9829), .A2(n13214), .ZN(n38020));
    INVX1 U25149 (.I(n15777), .ZN(n38021));
    NANDX1 U25150 (.A1(N6269), .A2(N3782), .ZN(N38022));
    INVX1 U25151 (.I(N5600), .ZN(N38023));
    NANDX1 U25152 (.A1(N11635), .A2(n22209), .ZN(N38024));
    NANDX1 U25153 (.A1(N5377), .A2(n23698), .ZN(N38025));
    INVX1 U25154 (.I(n15371), .ZN(N38026));
    INVX1 U25155 (.I(n24730), .ZN(N38027));
    INVX1 U25156 (.I(N12367), .ZN(n38028));
    NANDX1 U25157 (.A1(N7874), .A2(N2436), .ZN(N38029));
    NOR2X1 U25158 (.A1(n16490), .A2(N1874), .ZN(N38030));
    NANDX1 U25159 (.A1(N12135), .A2(N7184), .ZN(N38031));
    INVX1 U25160 (.I(n21963), .ZN(N38032));
    NOR2X1 U25161 (.A1(N1954), .A2(N7603), .ZN(N38033));
    NANDX1 U25162 (.A1(N8222), .A2(n30082), .ZN(N38034));
    NOR2X1 U25163 (.A1(N2383), .A2(N10044), .ZN(N38035));
    NOR2X1 U25164 (.A1(n24591), .A2(n25360), .ZN(n38036));
    NOR2X1 U25165 (.A1(n18152), .A2(N945), .ZN(n38037));
    INVX1 U25166 (.I(n19390), .ZN(n38038));
    NOR2X1 U25167 (.A1(N2335), .A2(n20317), .ZN(n38039));
    NANDX1 U25168 (.A1(n28906), .A2(n22752), .ZN(N38040));
    NANDX1 U25169 (.A1(n15258), .A2(n24625), .ZN(N38041));
    INVX1 U25170 (.I(n15953), .ZN(n38042));
    NOR2X1 U25171 (.A1(N6798), .A2(N7779), .ZN(N38043));
    NOR2X1 U25172 (.A1(N8751), .A2(N3942), .ZN(n38044));
    INVX1 U25173 (.I(n16973), .ZN(N38045));
    INVX1 U25174 (.I(N349), .ZN(N38046));
    INVX1 U25175 (.I(N2490), .ZN(N38047));
    INVX1 U25176 (.I(N2369), .ZN(N38048));
    NANDX1 U25177 (.A1(N2528), .A2(N9081), .ZN(N38049));
    INVX1 U25178 (.I(n25305), .ZN(N38050));
    NANDX1 U25179 (.A1(n20151), .A2(n16200), .ZN(N38051));
    INVX1 U25180 (.I(n22411), .ZN(N38052));
    INVX1 U25181 (.I(n18523), .ZN(N38053));
    NANDX1 U25182 (.A1(n18786), .A2(N1571), .ZN(N38054));
    NOR2X1 U25183 (.A1(N4602), .A2(n21940), .ZN(N38055));
    NANDX1 U25184 (.A1(N941), .A2(n21130), .ZN(N38056));
    NOR2X1 U25185 (.A1(N4882), .A2(N8204), .ZN(N38057));
    NANDX1 U25186 (.A1(n27465), .A2(n27250), .ZN(n38058));
    NOR2X1 U25187 (.A1(n18516), .A2(n29629), .ZN(N38059));
    NANDX1 U25188 (.A1(N4789), .A2(n20717), .ZN(n38060));
    NANDX1 U25189 (.A1(N10704), .A2(n15884), .ZN(n38061));
    NOR2X1 U25190 (.A1(n19416), .A2(n20645), .ZN(N38062));
    NANDX1 U25191 (.A1(N11689), .A2(N5475), .ZN(N38063));
    INVX1 U25192 (.I(N5112), .ZN(N38064));
    NANDX1 U25193 (.A1(N10705), .A2(n14191), .ZN(N38065));
    NOR2X1 U25194 (.A1(N2508), .A2(n30068), .ZN(N38066));
    NANDX1 U25195 (.A1(N12198), .A2(n13119), .ZN(N38067));
    INVX1 U25196 (.I(n20401), .ZN(n38068));
    INVX1 U25197 (.I(n16391), .ZN(N38069));
    NANDX1 U25198 (.A1(n21080), .A2(N4769), .ZN(n38070));
    INVX1 U25199 (.I(n19947), .ZN(N38071));
    INVX1 U25200 (.I(n26281), .ZN(n38072));
    NOR2X1 U25201 (.A1(n27520), .A2(N589), .ZN(n38073));
    INVX1 U25202 (.I(n16798), .ZN(N38074));
    NANDX1 U25203 (.A1(N1910), .A2(n17047), .ZN(N38075));
    INVX1 U25204 (.I(N11044), .ZN(n38076));
    NANDX1 U25205 (.A1(n28089), .A2(N10309), .ZN(N38077));
    NOR2X1 U25206 (.A1(N3935), .A2(N1377), .ZN(N38078));
    NANDX1 U25207 (.A1(n29556), .A2(n13575), .ZN(n38079));
    NANDX1 U25208 (.A1(n29921), .A2(n22536), .ZN(N38080));
    NANDX1 U25209 (.A1(N4736), .A2(n28610), .ZN(n38081));
    NANDX1 U25210 (.A1(n28202), .A2(n22735), .ZN(N38082));
    NANDX1 U25211 (.A1(n26320), .A2(n18879), .ZN(N38083));
    NANDX1 U25212 (.A1(N12263), .A2(N8028), .ZN(N38084));
    NANDX1 U25213 (.A1(n17621), .A2(n29260), .ZN(n38085));
    INVX1 U25214 (.I(N4530), .ZN(n38086));
    NOR2X1 U25215 (.A1(n15359), .A2(n15248), .ZN(n38087));
    NOR2X1 U25216 (.A1(n25668), .A2(N10019), .ZN(N38088));
    INVX1 U25217 (.I(n27044), .ZN(n38089));
    NOR2X1 U25218 (.A1(n22954), .A2(n29179), .ZN(N38090));
    INVX1 U25219 (.I(N11298), .ZN(N38091));
    NOR2X1 U25220 (.A1(n17882), .A2(n16033), .ZN(N38092));
    NANDX1 U25221 (.A1(n25604), .A2(n14098), .ZN(N38093));
    NANDX1 U25222 (.A1(n23136), .A2(n28978), .ZN(N38094));
    NOR2X1 U25223 (.A1(n25685), .A2(n29801), .ZN(N38095));
    INVX1 U25224 (.I(n20832), .ZN(N38096));
    NOR2X1 U25225 (.A1(n15796), .A2(n25148), .ZN(N38097));
    NANDX1 U25226 (.A1(n18747), .A2(N10369), .ZN(N38098));
    NANDX1 U25227 (.A1(N8210), .A2(N5899), .ZN(N38099));
    NANDX1 U25228 (.A1(N1607), .A2(n21504), .ZN(N38100));
    INVX1 U25229 (.I(n13121), .ZN(n38101));
    INVX1 U25230 (.I(n25841), .ZN(n38102));
    NANDX1 U25231 (.A1(N546), .A2(n13585), .ZN(N38103));
    NOR2X1 U25232 (.A1(N9156), .A2(n27749), .ZN(N38104));
    INVX1 U25233 (.I(N10364), .ZN(N38105));
    INVX1 U25234 (.I(n19071), .ZN(n38106));
    NANDX1 U25235 (.A1(N4856), .A2(n18734), .ZN(n38107));
    INVX1 U25236 (.I(n14248), .ZN(N38108));
    NOR2X1 U25237 (.A1(n21342), .A2(N9258), .ZN(N38109));
    INVX1 U25238 (.I(N9951), .ZN(n38110));
    INVX1 U25239 (.I(n18995), .ZN(N38111));
    NOR2X1 U25240 (.A1(n14086), .A2(n13058), .ZN(n38112));
    NOR2X1 U25241 (.A1(n24150), .A2(N401), .ZN(N38113));
    NANDX1 U25242 (.A1(N3119), .A2(n14802), .ZN(N38114));
    NOR2X1 U25243 (.A1(n22362), .A2(n28386), .ZN(n38115));
    INVX1 U25244 (.I(n20079), .ZN(N38116));
    INVX1 U25245 (.I(N11956), .ZN(N38117));
    NANDX1 U25246 (.A1(N5169), .A2(n19588), .ZN(N38118));
    NOR2X1 U25247 (.A1(N10024), .A2(n26882), .ZN(N38119));
    INVX1 U25248 (.I(N12832), .ZN(n38120));
    NANDX1 U25249 (.A1(N4626), .A2(n22090), .ZN(N38121));
    NOR2X1 U25250 (.A1(N3137), .A2(N11579), .ZN(N38122));
    NOR2X1 U25251 (.A1(N9858), .A2(n14225), .ZN(n38123));
    INVX1 U25252 (.I(n18185), .ZN(N38124));
    NOR2X1 U25253 (.A1(n17012), .A2(n28193), .ZN(N38125));
    INVX1 U25254 (.I(n20375), .ZN(N38126));
    INVX1 U25255 (.I(N10839), .ZN(N38127));
    NANDX1 U25256 (.A1(N12769), .A2(N780), .ZN(N38128));
    NOR2X1 U25257 (.A1(n13285), .A2(N1084), .ZN(N38129));
    NANDX1 U25258 (.A1(N2735), .A2(N8959), .ZN(n38130));
    NANDX1 U25259 (.A1(n29617), .A2(n22379), .ZN(n38131));
    NOR2X1 U25260 (.A1(N9363), .A2(n15565), .ZN(N38132));
    INVX1 U25261 (.I(n24059), .ZN(N38133));
    INVX1 U25262 (.I(N280), .ZN(N38134));
    NOR2X1 U25263 (.A1(n28559), .A2(N3065), .ZN(N38135));
    NOR2X1 U25264 (.A1(N5167), .A2(n30000), .ZN(N38136));
    NOR2X1 U25265 (.A1(N3222), .A2(n29916), .ZN(N38137));
    INVX1 U25266 (.I(n24265), .ZN(n38138));
    NOR2X1 U25267 (.A1(n17080), .A2(n25594), .ZN(N38139));
    INVX1 U25268 (.I(N8685), .ZN(n38140));
    INVX1 U25269 (.I(N1042), .ZN(N38141));
    NANDX1 U25270 (.A1(N37), .A2(n28698), .ZN(N38142));
    NANDX1 U25271 (.A1(n18214), .A2(N9500), .ZN(N38143));
    INVX1 U25272 (.I(n16137), .ZN(N38144));
    NOR2X1 U25273 (.A1(n16401), .A2(N10059), .ZN(N38145));
    NOR2X1 U25274 (.A1(N5241), .A2(n26232), .ZN(N38146));
    NANDX1 U25275 (.A1(n27003), .A2(n28880), .ZN(N38147));
    INVX1 U25276 (.I(n26866), .ZN(N38148));
    NANDX1 U25277 (.A1(N8998), .A2(n15205), .ZN(N38149));
    NOR2X1 U25278 (.A1(n21824), .A2(n14383), .ZN(N38150));
    NANDX1 U25279 (.A1(N5841), .A2(n14341), .ZN(N38151));
    NOR2X1 U25280 (.A1(N3143), .A2(N3943), .ZN(N38152));
    NOR2X1 U25281 (.A1(n21878), .A2(n21201), .ZN(N38153));
    INVX1 U25282 (.I(n28652), .ZN(N38154));
    INVX1 U25283 (.I(n19396), .ZN(N38155));
    NANDX1 U25284 (.A1(n25627), .A2(n24357), .ZN(n38156));
    NOR2X1 U25285 (.A1(n27816), .A2(n18158), .ZN(N38157));
    INVX1 U25286 (.I(n16987), .ZN(n38158));
    INVX1 U25287 (.I(n26805), .ZN(N38159));
    NANDX1 U25288 (.A1(N312), .A2(N3630), .ZN(N38160));
    NANDX1 U25289 (.A1(n15517), .A2(n27747), .ZN(N38161));
    INVX1 U25290 (.I(n18460), .ZN(n38162));
    NANDX1 U25291 (.A1(N6409), .A2(n21361), .ZN(N38163));
    NANDX1 U25292 (.A1(n28250), .A2(n25303), .ZN(N38164));
    INVX1 U25293 (.I(n19990), .ZN(n38165));
    NOR2X1 U25294 (.A1(n15172), .A2(n18504), .ZN(N38166));
    INVX1 U25295 (.I(n23128), .ZN(n38167));
    NANDX1 U25296 (.A1(n19677), .A2(n17347), .ZN(N38168));
    NANDX1 U25297 (.A1(N5917), .A2(N5367), .ZN(n38169));
    NOR2X1 U25298 (.A1(n22903), .A2(N8951), .ZN(n38170));
    INVX1 U25299 (.I(N4090), .ZN(N38171));
    NOR2X1 U25300 (.A1(N10331), .A2(n12972), .ZN(n38172));
    NANDX1 U25301 (.A1(N7940), .A2(N2101), .ZN(n38173));
    NOR2X1 U25302 (.A1(n16609), .A2(N8509), .ZN(n38174));
    INVX1 U25303 (.I(n14885), .ZN(N38175));
    NANDX1 U25304 (.A1(n25447), .A2(n15482), .ZN(n38176));
    INVX1 U25305 (.I(N236), .ZN(N38177));
    NANDX1 U25306 (.A1(n22236), .A2(n24423), .ZN(N38178));
    INVX1 U25307 (.I(n13814), .ZN(N38179));
    INVX1 U25308 (.I(n18113), .ZN(n38180));
    NANDX1 U25309 (.A1(N8440), .A2(n23479), .ZN(n38181));
    NANDX1 U25310 (.A1(n19903), .A2(n20990), .ZN(N38182));
    NANDX1 U25311 (.A1(n23992), .A2(n18813), .ZN(N38183));
    INVX1 U25312 (.I(n25524), .ZN(n38184));
    NOR2X1 U25313 (.A1(N651), .A2(n27624), .ZN(n38185));
    NANDX1 U25314 (.A1(n17259), .A2(n24694), .ZN(N38186));
    NOR2X1 U25315 (.A1(n20704), .A2(n19875), .ZN(N38187));
    NOR2X1 U25316 (.A1(N6049), .A2(N4909), .ZN(N38188));
    INVX1 U25317 (.I(n25263), .ZN(N38189));
    INVX1 U25318 (.I(N12347), .ZN(N38190));
    NANDX1 U25319 (.A1(n29518), .A2(n14870), .ZN(N38191));
    INVX1 U25320 (.I(n25302), .ZN(N38192));
    NANDX1 U25321 (.A1(n26043), .A2(N982), .ZN(N38193));
    INVX1 U25322 (.I(n16895), .ZN(N38194));
    INVX1 U25323 (.I(n14188), .ZN(n38195));
    NOR2X1 U25324 (.A1(n29088), .A2(N9574), .ZN(N38196));
    INVX1 U25325 (.I(n29738), .ZN(N38197));
    INVX1 U25326 (.I(n18517), .ZN(n38198));
    NOR2X1 U25327 (.A1(n20315), .A2(N10896), .ZN(N38199));
    INVX1 U25328 (.I(N10052), .ZN(n38200));
    NANDX1 U25329 (.A1(n20733), .A2(n14960), .ZN(n38201));
    NOR2X1 U25330 (.A1(N4419), .A2(n19225), .ZN(N38202));
    INVX1 U25331 (.I(N310), .ZN(n38203));
    NANDX1 U25332 (.A1(N9543), .A2(n14312), .ZN(N38204));
    INVX1 U25333 (.I(n21412), .ZN(N38205));
    INVX1 U25334 (.I(N3313), .ZN(N38206));
    INVX1 U25335 (.I(n27112), .ZN(N38207));
    NOR2X1 U25336 (.A1(N7096), .A2(n21242), .ZN(n38208));
    NOR2X1 U25337 (.A1(N5231), .A2(n17386), .ZN(N38209));
    INVX1 U25338 (.I(N852), .ZN(N38210));
    NOR2X1 U25339 (.A1(n28042), .A2(n21166), .ZN(n38211));
    NANDX1 U25340 (.A1(N12589), .A2(N1080), .ZN(N38212));
    INVX1 U25341 (.I(N3185), .ZN(N38213));
    INVX1 U25342 (.I(N4831), .ZN(n38214));
    NANDX1 U25343 (.A1(n23825), .A2(N10943), .ZN(n38215));
    INVX1 U25344 (.I(N854), .ZN(n38216));
    INVX1 U25345 (.I(N10785), .ZN(N38217));
    NOR2X1 U25346 (.A1(N320), .A2(N9562), .ZN(N38218));
    NANDX1 U25347 (.A1(N11926), .A2(n25234), .ZN(n38219));
    INVX1 U25348 (.I(n19022), .ZN(N38220));
    NANDX1 U25349 (.A1(N4752), .A2(N12813), .ZN(N38221));
    NANDX1 U25350 (.A1(N8675), .A2(n13664), .ZN(N38222));
    INVX1 U25351 (.I(N6579), .ZN(n38223));
    NANDX1 U25352 (.A1(N10394), .A2(n19168), .ZN(N38224));
    INVX1 U25353 (.I(n21458), .ZN(N38225));
    INVX1 U25354 (.I(n17630), .ZN(N38226));
    NOR2X1 U25355 (.A1(n25774), .A2(n30016), .ZN(N38227));
    INVX1 U25356 (.I(n22247), .ZN(N38228));
    NOR2X1 U25357 (.A1(N4699), .A2(n21592), .ZN(n38229));
    NANDX1 U25358 (.A1(n23716), .A2(N1016), .ZN(N38230));
    NOR2X1 U25359 (.A1(N5504), .A2(n26250), .ZN(n38231));
    INVX1 U25360 (.I(n13086), .ZN(N38232));
    INVX1 U25361 (.I(n18672), .ZN(N38233));
    NANDX1 U25362 (.A1(n23296), .A2(n15907), .ZN(N38234));
    INVX1 U25363 (.I(N9770), .ZN(N38235));
    INVX1 U25364 (.I(N2676), .ZN(n38236));
    NOR2X1 U25365 (.A1(N77), .A2(n15706), .ZN(N38237));
    NOR2X1 U25366 (.A1(n29687), .A2(N3198), .ZN(N38238));
    NOR2X1 U25367 (.A1(n25323), .A2(n21774), .ZN(n38239));
    NOR2X1 U25368 (.A1(N5993), .A2(N11067), .ZN(N38240));
    INVX1 U25369 (.I(n27584), .ZN(n38241));
    NOR2X1 U25370 (.A1(n16080), .A2(n17161), .ZN(n38242));
    INVX1 U25371 (.I(n21583), .ZN(N38243));
    NANDX1 U25372 (.A1(N8075), .A2(n23230), .ZN(n38244));
    NANDX1 U25373 (.A1(n26746), .A2(n18990), .ZN(N38245));
    NOR2X1 U25374 (.A1(N12516), .A2(n16975), .ZN(N38246));
    NOR2X1 U25375 (.A1(n23562), .A2(N8211), .ZN(N38247));
    NANDX1 U25376 (.A1(N12199), .A2(n23916), .ZN(N38248));
    INVX1 U25377 (.I(N309), .ZN(N38249));
    INVX1 U25378 (.I(n25249), .ZN(N38250));
    INVX1 U25379 (.I(N7311), .ZN(n38251));
    NOR2X1 U25380 (.A1(n20185), .A2(n18377), .ZN(n38252));
    NOR2X1 U25381 (.A1(N6192), .A2(n29179), .ZN(n38253));
    NANDX1 U25382 (.A1(n23352), .A2(n23334), .ZN(n38254));
    INVX1 U25383 (.I(n13746), .ZN(N38255));
    NOR2X1 U25384 (.A1(n13155), .A2(n16590), .ZN(n38256));
    INVX1 U25385 (.I(n20705), .ZN(n38257));
    NANDX1 U25386 (.A1(n29093), .A2(N7542), .ZN(n38258));
    INVX1 U25387 (.I(N11078), .ZN(N38259));
    NANDX1 U25388 (.A1(n17240), .A2(n23276), .ZN(N38260));
    NANDX1 U25389 (.A1(n27597), .A2(n23584), .ZN(N38261));
    NANDX1 U25390 (.A1(N11270), .A2(N7638), .ZN(N38262));
    NANDX1 U25391 (.A1(n24184), .A2(n27822), .ZN(N38263));
    NANDX1 U25392 (.A1(n18024), .A2(N3877), .ZN(N38264));
    NANDX1 U25393 (.A1(n16503), .A2(n15789), .ZN(n38265));
    INVX1 U25394 (.I(N6428), .ZN(n38266));
    NANDX1 U25395 (.A1(n28781), .A2(N8143), .ZN(N38267));
    NOR2X1 U25396 (.A1(n15221), .A2(n28848), .ZN(N38268));
    INVX1 U25397 (.I(N2737), .ZN(n38269));
    NOR2X1 U25398 (.A1(n19885), .A2(n13814), .ZN(N38270));
    INVX1 U25399 (.I(n25685), .ZN(N38271));
    NANDX1 U25400 (.A1(n27355), .A2(N11705), .ZN(n38272));
    NOR2X1 U25401 (.A1(N10983), .A2(n22974), .ZN(n38273));
    NOR2X1 U25402 (.A1(n20620), .A2(N5582), .ZN(n38274));
    NANDX1 U25403 (.A1(n25756), .A2(n23605), .ZN(N38275));
    NOR2X1 U25404 (.A1(N11234), .A2(n28668), .ZN(N38276));
    INVX1 U25405 (.I(n27305), .ZN(N38277));
    NOR2X1 U25406 (.A1(N9162), .A2(n14509), .ZN(N38278));
    NOR2X1 U25407 (.A1(N2271), .A2(n18290), .ZN(N38279));
    NOR2X1 U25408 (.A1(n26669), .A2(n21026), .ZN(n38280));
    NOR2X1 U25409 (.A1(N4977), .A2(n23400), .ZN(N38281));
    INVX1 U25410 (.I(N524), .ZN(n38282));
    INVX1 U25411 (.I(N10225), .ZN(N38283));
    NANDX1 U25412 (.A1(n26568), .A2(N9769), .ZN(N38284));
    INVX1 U25413 (.I(N11724), .ZN(N38285));
    INVX1 U25414 (.I(n29344), .ZN(n38286));
    NANDX1 U25415 (.A1(n14567), .A2(N11372), .ZN(N38287));
    INVX1 U25416 (.I(n14362), .ZN(N38288));
    NOR2X1 U25417 (.A1(n28443), .A2(N11529), .ZN(N38289));
    NANDX1 U25418 (.A1(N7467), .A2(n26037), .ZN(N38290));
    NANDX1 U25419 (.A1(n28435), .A2(n14189), .ZN(n38291));
    NANDX1 U25420 (.A1(n24967), .A2(n23775), .ZN(n38292));
    NANDX1 U25421 (.A1(n29943), .A2(n17037), .ZN(N38293));
    NANDX1 U25422 (.A1(N330), .A2(n24509), .ZN(N38294));
    INVX1 U25423 (.I(N1119), .ZN(n38295));
    INVX1 U25424 (.I(N6581), .ZN(N38296));
    INVX1 U25425 (.I(n21223), .ZN(N38297));
    INVX1 U25426 (.I(N12649), .ZN(n38298));
    NOR2X1 U25427 (.A1(N9959), .A2(n24020), .ZN(N38299));
    NOR2X1 U25428 (.A1(n24320), .A2(N3785), .ZN(n38300));
    NANDX1 U25429 (.A1(N5711), .A2(n25904), .ZN(n38301));
    NANDX1 U25430 (.A1(n20308), .A2(n19548), .ZN(N38302));
    INVX1 U25431 (.I(N4359), .ZN(n38303));
    NANDX1 U25432 (.A1(n29183), .A2(n28133), .ZN(N38304));
    NOR2X1 U25433 (.A1(n28989), .A2(N3593), .ZN(N38305));
    NANDX1 U25434 (.A1(n17879), .A2(n28101), .ZN(n38306));
    NANDX1 U25435 (.A1(N7558), .A2(N7463), .ZN(N38307));
    NANDX1 U25436 (.A1(N2301), .A2(n28685), .ZN(N38308));
    INVX1 U25437 (.I(n14949), .ZN(N38309));
    INVX1 U25438 (.I(n19868), .ZN(n38310));
    INVX1 U25439 (.I(n14483), .ZN(n38311));
    NOR2X1 U25440 (.A1(n19875), .A2(N5676), .ZN(N38312));
    NANDX1 U25441 (.A1(n15642), .A2(N11595), .ZN(N38313));
    INVX1 U25442 (.I(n23750), .ZN(N38314));
    INVX1 U25443 (.I(N10108), .ZN(N38315));
    NOR2X1 U25444 (.A1(n14857), .A2(n26801), .ZN(N38316));
    NANDX1 U25445 (.A1(N2269), .A2(n18954), .ZN(n38317));
    INVX1 U25446 (.I(n20147), .ZN(N38318));
    INVX1 U25447 (.I(N9200), .ZN(N38319));
    NOR2X1 U25448 (.A1(n12940), .A2(n23717), .ZN(n38320));
    INVX1 U25449 (.I(N11487), .ZN(N38321));
    NANDX1 U25450 (.A1(n22075), .A2(N2944), .ZN(N38322));
    NOR2X1 U25451 (.A1(n19467), .A2(n17426), .ZN(n38323));
    NOR2X1 U25452 (.A1(N9205), .A2(N11662), .ZN(N38324));
    INVX1 U25453 (.I(n13407), .ZN(N38325));
    NOR2X1 U25454 (.A1(N5718), .A2(n25717), .ZN(N38326));
    INVX1 U25455 (.I(N4386), .ZN(n38327));
    NANDX1 U25456 (.A1(N909), .A2(N1049), .ZN(N38328));
    INVX1 U25457 (.I(N3178), .ZN(N38329));
    INVX1 U25458 (.I(n15928), .ZN(n38330));
    INVX1 U25459 (.I(n25479), .ZN(N38331));
    NOR2X1 U25460 (.A1(N9452), .A2(N8281), .ZN(N38332));
    NANDX1 U25461 (.A1(n28017), .A2(N8329), .ZN(n38333));
    INVX1 U25462 (.I(n19954), .ZN(n38334));
    INVX1 U25463 (.I(n22673), .ZN(N38335));
    INVX1 U25464 (.I(n28697), .ZN(N38336));
    INVX1 U25465 (.I(N7049), .ZN(N38337));
    INVX1 U25466 (.I(n14290), .ZN(N38338));
    NOR2X1 U25467 (.A1(n22038), .A2(N8568), .ZN(N38339));
    NANDX1 U25468 (.A1(N8090), .A2(n12954), .ZN(N38340));
    INVX1 U25469 (.I(N8999), .ZN(N38341));
    NANDX1 U25470 (.A1(n17834), .A2(N12176), .ZN(N38342));
    NOR2X1 U25471 (.A1(N3624), .A2(n24060), .ZN(n38343));
    INVX1 U25472 (.I(n17312), .ZN(n38344));
    NOR2X1 U25473 (.A1(N3309), .A2(n24579), .ZN(N38345));
    INVX1 U25474 (.I(N198), .ZN(N38346));
    NANDX1 U25475 (.A1(n28466), .A2(N11469), .ZN(n38347));
    NOR2X1 U25476 (.A1(n14871), .A2(n28726), .ZN(n38348));
    INVX1 U25477 (.I(n21919), .ZN(N38349));
    NANDX1 U25478 (.A1(N3464), .A2(n19495), .ZN(N38350));
    NOR2X1 U25479 (.A1(N12031), .A2(N12650), .ZN(N38351));
    INVX1 U25480 (.I(n13545), .ZN(n38352));
    INVX1 U25481 (.I(n25056), .ZN(N38353));
    NOR2X1 U25482 (.A1(n22211), .A2(n25792), .ZN(N38354));
    NOR2X1 U25483 (.A1(n14395), .A2(N8276), .ZN(n38355));
    NOR2X1 U25484 (.A1(n20267), .A2(N210), .ZN(n38356));
    INVX1 U25485 (.I(N3269), .ZN(n38357));
    INVX1 U25486 (.I(N2887), .ZN(n38358));
    INVX1 U25487 (.I(n25748), .ZN(N38359));
    NOR2X1 U25488 (.A1(N2017), .A2(N10481), .ZN(N38360));
    NOR2X1 U25489 (.A1(n21328), .A2(n20960), .ZN(n38361));
    NANDX1 U25490 (.A1(n13352), .A2(N10317), .ZN(N38362));
    NANDX1 U25491 (.A1(n13944), .A2(n22966), .ZN(n38363));
    NOR2X1 U25492 (.A1(n27488), .A2(n15904), .ZN(n38364));
    INVX1 U25493 (.I(N2019), .ZN(N38365));
    INVX1 U25494 (.I(N2033), .ZN(n38366));
    INVX1 U25495 (.I(N10932), .ZN(n38367));
    INVX1 U25496 (.I(n17194), .ZN(N38368));
    NANDX1 U25497 (.A1(N10518), .A2(n19883), .ZN(N38369));
    NOR2X1 U25498 (.A1(n19239), .A2(N11331), .ZN(n38370));
    NOR2X1 U25499 (.A1(N3410), .A2(n14246), .ZN(N38371));
    NOR2X1 U25500 (.A1(n13890), .A2(N4311), .ZN(N38372));
    NOR2X1 U25501 (.A1(N4712), .A2(N3184), .ZN(n38373));
    NANDX1 U25502 (.A1(N3589), .A2(N10025), .ZN(N38374));
    INVX1 U25503 (.I(n26554), .ZN(N38375));
    NANDX1 U25504 (.A1(n15028), .A2(N881), .ZN(N38376));
    NANDX1 U25505 (.A1(N5608), .A2(N8857), .ZN(n38377));
    INVX1 U25506 (.I(N11980), .ZN(N38378));
    NANDX1 U25507 (.A1(n21504), .A2(n29173), .ZN(N38379));
    NOR2X1 U25508 (.A1(n20582), .A2(N7480), .ZN(N38380));
    NOR2X1 U25509 (.A1(n28381), .A2(n18810), .ZN(N38381));
    NOR2X1 U25510 (.A1(N1653), .A2(n21616), .ZN(n38382));
    NANDX1 U25511 (.A1(N4103), .A2(n25926), .ZN(n38383));
    NOR2X1 U25512 (.A1(N8814), .A2(n29109), .ZN(N38384));
    INVX1 U25513 (.I(N12402), .ZN(N38385));
    NOR2X1 U25514 (.A1(n14642), .A2(n27516), .ZN(N38386));
    NANDX1 U25515 (.A1(n18230), .A2(n28396), .ZN(N38387));
    INVX1 U25516 (.I(N12398), .ZN(N38388));
    NOR2X1 U25517 (.A1(n16522), .A2(n24378), .ZN(N38389));
    NOR2X1 U25518 (.A1(n26587), .A2(N11974), .ZN(n38390));
    NANDX1 U25519 (.A1(n17031), .A2(N8014), .ZN(N38391));
    NANDX1 U25520 (.A1(N3836), .A2(n15384), .ZN(N38392));
    NANDX1 U25521 (.A1(n24186), .A2(N6863), .ZN(N38393));
    INVX1 U25522 (.I(n28289), .ZN(N38394));
    INVX1 U25523 (.I(n21625), .ZN(n38395));
    NANDX1 U25524 (.A1(N8882), .A2(N7150), .ZN(N38396));
    NANDX1 U25525 (.A1(N6438), .A2(N10352), .ZN(N38397));
    NANDX1 U25526 (.A1(n14039), .A2(n17143), .ZN(N38398));
    INVX1 U25527 (.I(n19365), .ZN(N38399));
    NANDX1 U25528 (.A1(n25197), .A2(N5749), .ZN(N38400));
    INVX1 U25529 (.I(n17782), .ZN(n38401));
    INVX1 U25530 (.I(n12876), .ZN(N38402));
    NOR2X1 U25531 (.A1(N7790), .A2(N9450), .ZN(N38403));
    NANDX1 U25532 (.A1(N11625), .A2(n24834), .ZN(N38404));
    INVX1 U25533 (.I(n24371), .ZN(N38405));
    NOR2X1 U25534 (.A1(n13559), .A2(n22522), .ZN(n38406));
    NOR2X1 U25535 (.A1(n23744), .A2(n29487), .ZN(N38407));
    NANDX1 U25536 (.A1(n19455), .A2(n25975), .ZN(N38408));
    NANDX1 U25537 (.A1(n18367), .A2(N8402), .ZN(N38409));
    NANDX1 U25538 (.A1(n24070), .A2(n19225), .ZN(N38410));
    INVX1 U25539 (.I(N12034), .ZN(N38411));
    NOR2X1 U25540 (.A1(n12923), .A2(n12935), .ZN(N38412));
    NOR2X1 U25541 (.A1(N3681), .A2(n14371), .ZN(N38413));
    NANDX1 U25542 (.A1(N11470), .A2(n23821), .ZN(n38414));
    INVX1 U25543 (.I(N11655), .ZN(N38415));
    NANDX1 U25544 (.A1(N6960), .A2(N5889), .ZN(N38416));
    INVX1 U25545 (.I(N9079), .ZN(n38417));
    INVX1 U25546 (.I(N8664), .ZN(N38418));
    NOR2X1 U25547 (.A1(n16320), .A2(n17574), .ZN(N38419));
    INVX1 U25548 (.I(N718), .ZN(n38420));
    INVX1 U25549 (.I(n17628), .ZN(N38421));
    INVX1 U25550 (.I(n20730), .ZN(N38422));
    INVX1 U25551 (.I(n28344), .ZN(N38423));
    NANDX1 U25552 (.A1(N12155), .A2(N1052), .ZN(N38424));
    INVX1 U25553 (.I(n25089), .ZN(n38425));
    NANDX1 U25554 (.A1(N2930), .A2(n28021), .ZN(N38426));
    NOR2X1 U25555 (.A1(n14400), .A2(n21704), .ZN(N38427));
    INVX1 U25556 (.I(n14615), .ZN(N38428));
    NOR2X1 U25557 (.A1(n26383), .A2(n20503), .ZN(N38429));
    INVX1 U25558 (.I(n24022), .ZN(N38430));
    NANDX1 U25559 (.A1(N11762), .A2(n15268), .ZN(N38431));
    NOR2X1 U25560 (.A1(n29335), .A2(N3090), .ZN(n38432));
    NANDX1 U25561 (.A1(n20679), .A2(N9279), .ZN(N38433));
    NANDX1 U25562 (.A1(n29970), .A2(N9400), .ZN(N38434));
    INVX1 U25563 (.I(n27736), .ZN(N38435));
    NANDX1 U25564 (.A1(n21312), .A2(n26985), .ZN(N38436));
    NANDX1 U25565 (.A1(N12853), .A2(n29914), .ZN(N38437));
    NANDX1 U25566 (.A1(N10479), .A2(N2737), .ZN(N38438));
    NOR2X1 U25567 (.A1(N11204), .A2(n17352), .ZN(N38439));
    NOR2X1 U25568 (.A1(n26147), .A2(n26415), .ZN(N38440));
    INVX1 U25569 (.I(n20031), .ZN(n38441));
    NOR2X1 U25570 (.A1(n26716), .A2(n23860), .ZN(n38442));
    NOR2X1 U25571 (.A1(n14474), .A2(n26949), .ZN(N38443));
    NANDX1 U25572 (.A1(n23714), .A2(n24788), .ZN(N38444));
    INVX1 U25573 (.I(n23546), .ZN(N38445));
    INVX1 U25574 (.I(n22242), .ZN(N38446));
    NANDX1 U25575 (.A1(n25603), .A2(N1977), .ZN(N38447));
    NOR2X1 U25576 (.A1(N532), .A2(n14829), .ZN(N38448));
    NANDX1 U25577 (.A1(n22178), .A2(n25308), .ZN(N38449));
    NOR2X1 U25578 (.A1(N5254), .A2(n25072), .ZN(n38450));
    NANDX1 U25579 (.A1(n17109), .A2(n21081), .ZN(n38451));
    NOR2X1 U25580 (.A1(n20624), .A2(n29672), .ZN(N38452));
    NOR2X1 U25581 (.A1(N5763), .A2(n23394), .ZN(N38453));
    NOR2X1 U25582 (.A1(N8797), .A2(N8767), .ZN(N38454));
    NANDX1 U25583 (.A1(N2373), .A2(N3417), .ZN(N38455));
    NANDX1 U25584 (.A1(n14479), .A2(N7467), .ZN(n38456));
    NOR2X1 U25585 (.A1(N12744), .A2(n21630), .ZN(n38457));
    INVX1 U25586 (.I(N7856), .ZN(N38458));
    NANDX1 U25587 (.A1(n24597), .A2(n21443), .ZN(N38459));
    NANDX1 U25588 (.A1(N8328), .A2(n26327), .ZN(N38460));
    NANDX1 U25589 (.A1(N3262), .A2(N6986), .ZN(N38461));
    NANDX1 U25590 (.A1(n12903), .A2(n25498), .ZN(N38462));
    NOR2X1 U25591 (.A1(N12438), .A2(N6048), .ZN(n38463));
    INVX1 U25592 (.I(n24392), .ZN(N38464));
    NANDX1 U25593 (.A1(N7291), .A2(N3021), .ZN(N38465));
    INVX1 U25594 (.I(N9663), .ZN(n38466));
    NANDX1 U25595 (.A1(N5863), .A2(N12703), .ZN(N38467));
    NOR2X1 U25596 (.A1(n25094), .A2(n25446), .ZN(N38468));
    INVX1 U25597 (.I(N4725), .ZN(N38469));
    NOR2X1 U25598 (.A1(N11938), .A2(n29321), .ZN(N38470));
    NANDX1 U25599 (.A1(n14700), .A2(N7512), .ZN(N38471));
    INVX1 U25600 (.I(N11276), .ZN(N38472));
    INVX1 U25601 (.I(N4903), .ZN(N38473));
    NOR2X1 U25602 (.A1(N12237), .A2(n18961), .ZN(N38474));
    NOR2X1 U25603 (.A1(n24674), .A2(n25009), .ZN(n38475));
    NOR2X1 U25604 (.A1(n18928), .A2(N8738), .ZN(N38476));
    INVX1 U25605 (.I(N10510), .ZN(n38477));
    INVX1 U25606 (.I(n21699), .ZN(N38478));
    INVX1 U25607 (.I(N12035), .ZN(N38479));
    NOR2X1 U25608 (.A1(n26670), .A2(N6991), .ZN(N38480));
    NANDX1 U25609 (.A1(n27885), .A2(N276), .ZN(n38481));
    NANDX1 U25610 (.A1(N9685), .A2(n29597), .ZN(N38482));
    INVX1 U25611 (.I(n24384), .ZN(N38483));
    NANDX1 U25612 (.A1(n21079), .A2(n24220), .ZN(n38484));
    NANDX1 U25613 (.A1(n14542), .A2(N7604), .ZN(n38485));
    NOR2X1 U25614 (.A1(N3366), .A2(n13856), .ZN(N38486));
    NOR2X1 U25615 (.A1(n28374), .A2(n18601), .ZN(N38487));
    NOR2X1 U25616 (.A1(n25672), .A2(N500), .ZN(N38488));
    NANDX1 U25617 (.A1(N1707), .A2(n22198), .ZN(N38489));
    NOR2X1 U25618 (.A1(N2303), .A2(n15022), .ZN(n38490));
    NOR2X1 U25619 (.A1(N9293), .A2(N3154), .ZN(n38491));
    NANDX1 U25620 (.A1(n28267), .A2(n13149), .ZN(n38492));
    INVX1 U25621 (.I(n27726), .ZN(N38493));
    INVX1 U25622 (.I(n26431), .ZN(N38494));
    NANDX1 U25623 (.A1(n15813), .A2(n20514), .ZN(N38495));
    INVX1 U25624 (.I(n18915), .ZN(N38496));
    NOR2X1 U25625 (.A1(n21042), .A2(N10841), .ZN(N38497));
    NOR2X1 U25626 (.A1(n29937), .A2(N9077), .ZN(N38498));
    NOR2X1 U25627 (.A1(n16184), .A2(n23310), .ZN(n38499));
    INVX1 U25628 (.I(n12940), .ZN(n38500));
    NOR2X1 U25629 (.A1(N116), .A2(n22462), .ZN(N38501));
    NANDX1 U25630 (.A1(N3698), .A2(n28516), .ZN(n38502));
    INVX1 U25631 (.I(n25550), .ZN(n38503));
    NANDX1 U25632 (.A1(N11862), .A2(N8561), .ZN(N38504));
    NANDX1 U25633 (.A1(n28148), .A2(N3294), .ZN(N38505));
    NANDX1 U25634 (.A1(N9828), .A2(N7667), .ZN(N38506));
    INVX1 U25635 (.I(N5070), .ZN(N38507));
    NANDX1 U25636 (.A1(N7574), .A2(n26111), .ZN(N38508));
    NOR2X1 U25637 (.A1(N7969), .A2(n14472), .ZN(N38509));
    NANDX1 U25638 (.A1(n15526), .A2(N518), .ZN(N38510));
    NANDX1 U25639 (.A1(n23581), .A2(N2019), .ZN(N38511));
    INVX1 U25640 (.I(n23697), .ZN(N38512));
    NANDX1 U25641 (.A1(N4672), .A2(n15955), .ZN(n38513));
    NANDX1 U25642 (.A1(n18404), .A2(N11367), .ZN(n38514));
    NOR2X1 U25643 (.A1(n18826), .A2(N8488), .ZN(N38515));
    NANDX1 U25644 (.A1(n16836), .A2(N343), .ZN(n38516));
    NOR2X1 U25645 (.A1(n26663), .A2(n26707), .ZN(N38517));
    NANDX1 U25646 (.A1(n20293), .A2(N11712), .ZN(N38518));
    INVX1 U25647 (.I(n16267), .ZN(n38519));
    INVX1 U25648 (.I(N6088), .ZN(N38520));
    NOR2X1 U25649 (.A1(N1041), .A2(N10174), .ZN(N38521));
    NANDX1 U25650 (.A1(N6394), .A2(N3617), .ZN(N38522));
    INVX1 U25651 (.I(n25323), .ZN(n38523));
    INVX1 U25652 (.I(N4738), .ZN(N38524));
    NANDX1 U25653 (.A1(N1692), .A2(n27596), .ZN(N38525));
    NOR2X1 U25654 (.A1(N1619), .A2(N11058), .ZN(n38526));
    NANDX1 U25655 (.A1(n28805), .A2(n28884), .ZN(N38527));
    NOR2X1 U25656 (.A1(n29147), .A2(n28532), .ZN(N38528));
    NANDX1 U25657 (.A1(n14277), .A2(n19077), .ZN(n38529));
    NANDX1 U25658 (.A1(n25989), .A2(n17196), .ZN(N38530));
    NANDX1 U25659 (.A1(n22107), .A2(N11844), .ZN(N38531));
    NANDX1 U25660 (.A1(N11708), .A2(n22017), .ZN(n38532));
    NOR2X1 U25661 (.A1(N6662), .A2(n25633), .ZN(N38533));
    INVX1 U25662 (.I(N1847), .ZN(n38534));
    NANDX1 U25663 (.A1(n27960), .A2(n20402), .ZN(N38535));
    NOR2X1 U25664 (.A1(n13979), .A2(n15783), .ZN(N38536));
    INVX1 U25665 (.I(n13597), .ZN(n38537));
    NANDX1 U25666 (.A1(n20605), .A2(N12343), .ZN(N38538));
    INVX1 U25667 (.I(N8175), .ZN(N38539));
    NANDX1 U25668 (.A1(n28324), .A2(N11013), .ZN(N38540));
    INVX1 U25669 (.I(N4470), .ZN(N38541));
    INVX1 U25670 (.I(N5433), .ZN(N38542));
    INVX1 U25671 (.I(n17531), .ZN(n38543));
    NOR2X1 U25672 (.A1(N8592), .A2(n29238), .ZN(N38544));
    NANDX1 U25673 (.A1(N9980), .A2(n24460), .ZN(N38545));
    NOR2X1 U25674 (.A1(n21763), .A2(n26306), .ZN(N38546));
    NANDX1 U25675 (.A1(N8146), .A2(n16570), .ZN(N38547));
    INVX1 U25676 (.I(N10685), .ZN(N38548));
    INVX1 U25677 (.I(n23959), .ZN(N38549));
    INVX1 U25678 (.I(n20766), .ZN(N38550));
    NANDX1 U25679 (.A1(n25184), .A2(n21522), .ZN(N38551));
    NOR2X1 U25680 (.A1(n24482), .A2(n19708), .ZN(N38552));
    NOR2X1 U25681 (.A1(N12719), .A2(N12738), .ZN(N38553));
    INVX1 U25682 (.I(n18151), .ZN(n38554));
    INVX1 U25683 (.I(N4991), .ZN(N38555));
    INVX1 U25684 (.I(N6771), .ZN(N38556));
    NOR2X1 U25685 (.A1(n21702), .A2(N5312), .ZN(N38557));
    INVX1 U25686 (.I(N3473), .ZN(N38558));
    NOR2X1 U25687 (.A1(N1840), .A2(n15312), .ZN(N38559));
    INVX1 U25688 (.I(N6971), .ZN(n38560));
    INVX1 U25689 (.I(N4328), .ZN(N38561));
    NOR2X1 U25690 (.A1(N11153), .A2(n17170), .ZN(N38562));
    NANDX1 U25691 (.A1(n14140), .A2(N12216), .ZN(N38563));
    NANDX1 U25692 (.A1(n13862), .A2(n25258), .ZN(n38564));
    INVX1 U25693 (.I(N5898), .ZN(n38565));
    INVX1 U25694 (.I(N765), .ZN(n38566));
    NOR2X1 U25695 (.A1(n14550), .A2(n29082), .ZN(N38567));
    NOR2X1 U25696 (.A1(N8399), .A2(N5715), .ZN(n38568));
    NANDX1 U25697 (.A1(n18661), .A2(N11026), .ZN(N38569));
    NOR2X1 U25698 (.A1(N10695), .A2(n26661), .ZN(N38570));
    NANDX1 U25699 (.A1(n14567), .A2(N8865), .ZN(N38571));
    INVX1 U25700 (.I(N1761), .ZN(N38572));
    INVX1 U25701 (.I(n17743), .ZN(N38573));
    INVX1 U25702 (.I(N224), .ZN(N38574));
    NANDX1 U25703 (.A1(n15614), .A2(N1001), .ZN(N38575));
    NANDX1 U25704 (.A1(n29475), .A2(n14819), .ZN(N38576));
    NANDX1 U25705 (.A1(n23933), .A2(N11219), .ZN(N38577));
    NOR2X1 U25706 (.A1(N5851), .A2(n25768), .ZN(n38578));
    NANDX1 U25707 (.A1(N11457), .A2(n22728), .ZN(N38579));
    NANDX1 U25708 (.A1(n28412), .A2(n29949), .ZN(N38580));
    NANDX1 U25709 (.A1(n20901), .A2(N10506), .ZN(n38581));
    NOR2X1 U25710 (.A1(n15229), .A2(n25072), .ZN(N38582));
    INVX1 U25711 (.I(n16528), .ZN(N38583));
    NANDX1 U25712 (.A1(N12009), .A2(N4133), .ZN(n38584));
    NANDX1 U25713 (.A1(N793), .A2(n28948), .ZN(N38585));
    INVX1 U25714 (.I(n20491), .ZN(N38586));
    INVX1 U25715 (.I(n20379), .ZN(N38587));
    INVX1 U25716 (.I(n14682), .ZN(N38588));
    NOR2X1 U25717 (.A1(n16391), .A2(n26744), .ZN(N38589));
    NANDX1 U25718 (.A1(N582), .A2(n26312), .ZN(n38590));
    INVX1 U25719 (.I(n23309), .ZN(N38591));
    NOR2X1 U25720 (.A1(n18315), .A2(N11682), .ZN(n38592));
    NANDX1 U25721 (.A1(N9078), .A2(n22187), .ZN(n38593));
    NANDX1 U25722 (.A1(n24306), .A2(N5683), .ZN(n38594));
    NANDX1 U25723 (.A1(n29394), .A2(n21076), .ZN(n38595));
    INVX1 U25724 (.I(n22088), .ZN(N38596));
    NANDX1 U25725 (.A1(n15154), .A2(n20898), .ZN(N38597));
    NOR2X1 U25726 (.A1(N5507), .A2(N12842), .ZN(N38598));
    NANDX1 U25727 (.A1(n29377), .A2(n27523), .ZN(N38599));
    NANDX1 U25728 (.A1(n15630), .A2(N12690), .ZN(n38600));
    INVX1 U25729 (.I(n16212), .ZN(n38601));
    NOR2X1 U25730 (.A1(N8870), .A2(n28081), .ZN(N38602));
    NOR2X1 U25731 (.A1(n27184), .A2(N9625), .ZN(n38603));
    NANDX1 U25732 (.A1(n24822), .A2(n20373), .ZN(N38604));
    NOR2X1 U25733 (.A1(n18990), .A2(n14616), .ZN(n38605));
    INVX1 U25734 (.I(N6808), .ZN(n38606));
    NOR2X1 U25735 (.A1(n25455), .A2(n28895), .ZN(n38607));
    INVX1 U25736 (.I(n29169), .ZN(N38608));
    NOR2X1 U25737 (.A1(N7888), .A2(n23236), .ZN(N38609));
    NOR2X1 U25738 (.A1(N4097), .A2(n22476), .ZN(n38610));
    NANDX1 U25739 (.A1(n14479), .A2(N7968), .ZN(n38611));
    NANDX1 U25740 (.A1(N3308), .A2(N12740), .ZN(n38612));
    NOR2X1 U25741 (.A1(N12177), .A2(n29382), .ZN(n38613));
    NANDX1 U25742 (.A1(n27921), .A2(n27567), .ZN(N38614));
    NOR2X1 U25743 (.A1(n22605), .A2(N6363), .ZN(N38615));
    NOR2X1 U25744 (.A1(N18), .A2(n20978), .ZN(N38616));
    NANDX1 U25745 (.A1(N6825), .A2(n15092), .ZN(n38617));
    INVX1 U25746 (.I(n24280), .ZN(N38618));
    NOR2X1 U25747 (.A1(N4147), .A2(N2358), .ZN(N38619));
    NANDX1 U25748 (.A1(n27382), .A2(n23414), .ZN(N38620));
    NOR2X1 U25749 (.A1(n19720), .A2(N279), .ZN(n38621));
    NOR2X1 U25750 (.A1(n16249), .A2(N8532), .ZN(N38622));
    NANDX1 U25751 (.A1(n17549), .A2(n14209), .ZN(N38623));
    NANDX1 U25752 (.A1(N5354), .A2(n26025), .ZN(n38624));
    NANDX1 U25753 (.A1(N2784), .A2(n20169), .ZN(n38625));
    INVX1 U25754 (.I(N9146), .ZN(n38626));
    INVX1 U25755 (.I(N10726), .ZN(N38627));
    NOR2X1 U25756 (.A1(N2714), .A2(N6111), .ZN(N38628));
    INVX1 U25757 (.I(N7829), .ZN(N38629));
    NANDX1 U25758 (.A1(n16470), .A2(N536), .ZN(N38630));
    INVX1 U25759 (.I(n18489), .ZN(N38631));
    INVX1 U25760 (.I(n14586), .ZN(N38632));
    INVX1 U25761 (.I(N6061), .ZN(N38633));
    NOR2X1 U25762 (.A1(n22320), .A2(n22309), .ZN(N38634));
    NOR2X1 U25763 (.A1(n23343), .A2(n28419), .ZN(n38635));
    NANDX1 U25764 (.A1(N6404), .A2(N3635), .ZN(N38636));
    NOR2X1 U25765 (.A1(N5947), .A2(N6418), .ZN(N38637));
    INVX1 U25766 (.I(n16654), .ZN(N38638));
    NOR2X1 U25767 (.A1(N12257), .A2(n27379), .ZN(N38639));
    NANDX1 U25768 (.A1(N3532), .A2(n22051), .ZN(n38640));
    NOR2X1 U25769 (.A1(N11360), .A2(n22304), .ZN(n38641));
    INVX1 U25770 (.I(N11896), .ZN(n38642));
    INVX1 U25771 (.I(N8390), .ZN(N38643));
    NOR2X1 U25772 (.A1(n28060), .A2(N10116), .ZN(n38644));
    NANDX1 U25773 (.A1(N1348), .A2(n20996), .ZN(n38645));
    INVX1 U25774 (.I(n13303), .ZN(N38646));
    NANDX1 U25775 (.A1(N2009), .A2(n16589), .ZN(n38647));
    INVX1 U25776 (.I(N5643), .ZN(N38648));
    NOR2X1 U25777 (.A1(N3673), .A2(N622), .ZN(n38649));
    NOR2X1 U25778 (.A1(N8887), .A2(n23444), .ZN(N38650));
    INVX1 U25779 (.I(n24827), .ZN(n38651));
    NOR2X1 U25780 (.A1(N2055), .A2(n16740), .ZN(N38652));
    NOR2X1 U25781 (.A1(N1976), .A2(N8906), .ZN(N38653));
    NANDX1 U25782 (.A1(N2432), .A2(N10941), .ZN(N38654));
    NOR2X1 U25783 (.A1(N668), .A2(n27562), .ZN(N38655));
    NOR2X1 U25784 (.A1(n23662), .A2(n28909), .ZN(N38656));
    NANDX1 U25785 (.A1(n27389), .A2(N635), .ZN(N38657));
    NANDX1 U25786 (.A1(n29397), .A2(N5784), .ZN(N38658));
    NOR2X1 U25787 (.A1(n23601), .A2(N2847), .ZN(N38659));
    INVX1 U25788 (.I(N12783), .ZN(N38660));
    NOR2X1 U25789 (.A1(n27812), .A2(N6089), .ZN(n38661));
    INVX1 U25790 (.I(n22501), .ZN(N38662));
    INVX1 U25791 (.I(N8390), .ZN(N38663));
    NOR2X1 U25792 (.A1(N7568), .A2(N10365), .ZN(N38664));
    INVX1 U25793 (.I(N5712), .ZN(N38665));
    NANDX1 U25794 (.A1(n17510), .A2(N12245), .ZN(n38666));
    INVX1 U25795 (.I(N3495), .ZN(N38667));
    INVX1 U25796 (.I(N2808), .ZN(N38668));
    NOR2X1 U25797 (.A1(N2083), .A2(N59), .ZN(N38669));
    NOR2X1 U25798 (.A1(N912), .A2(n18017), .ZN(N38670));
    INVX1 U25799 (.I(n27604), .ZN(N38671));
    NOR2X1 U25800 (.A1(n18789), .A2(n16392), .ZN(N38672));
    INVX1 U25801 (.I(N7903), .ZN(n38673));
    NANDX1 U25802 (.A1(n18911), .A2(n14238), .ZN(N38674));
    INVX1 U25803 (.I(n18235), .ZN(N38675));
    NOR2X1 U25804 (.A1(N4093), .A2(n25802), .ZN(N38676));
    NANDX1 U25805 (.A1(N10662), .A2(N1377), .ZN(n38677));
    INVX1 U25806 (.I(n16732), .ZN(n38678));
    NOR2X1 U25807 (.A1(N2055), .A2(n20226), .ZN(N38679));
    INVX1 U25808 (.I(N4862), .ZN(N38680));
    INVX1 U25809 (.I(n28977), .ZN(n38681));
    NANDX1 U25810 (.A1(n21210), .A2(n29888), .ZN(N38682));
    INVX1 U25811 (.I(N7015), .ZN(n38683));
    INVX1 U25812 (.I(N98), .ZN(N38684));
    INVX1 U25813 (.I(n20867), .ZN(n38685));
    NOR2X1 U25814 (.A1(N10828), .A2(N4795), .ZN(N38686));
    NANDX1 U25815 (.A1(n25065), .A2(n29922), .ZN(N38687));
    INVX1 U25816 (.I(N6115), .ZN(N38688));
    NANDX1 U25817 (.A1(n22851), .A2(n16228), .ZN(N38689));
    INVX1 U25818 (.I(N12788), .ZN(n38690));
    INVX1 U25819 (.I(n19831), .ZN(n38691));
    INVX1 U25820 (.I(n18313), .ZN(n38692));
    INVX1 U25821 (.I(N11726), .ZN(n38693));
    NOR2X1 U25822 (.A1(N9531), .A2(N10565), .ZN(n38694));
    NANDX1 U25823 (.A1(n19301), .A2(n29013), .ZN(N38695));
    NOR2X1 U25824 (.A1(n14877), .A2(N3351), .ZN(N38696));
    NANDX1 U25825 (.A1(n29241), .A2(n24217), .ZN(N38697));
    NOR2X1 U25826 (.A1(n28629), .A2(n17573), .ZN(n38698));
    INVX1 U25827 (.I(n23556), .ZN(N38699));
    NANDX1 U25828 (.A1(N12851), .A2(n18231), .ZN(N38700));
    INVX1 U25829 (.I(N5564), .ZN(n38701));
    NOR2X1 U25830 (.A1(N1455), .A2(N6912), .ZN(n38702));
    NOR2X1 U25831 (.A1(N9846), .A2(N10441), .ZN(n38703));
    NANDX1 U25832 (.A1(N8325), .A2(N10728), .ZN(N38704));
    INVX1 U25833 (.I(N6416), .ZN(N38705));
    NANDX1 U25834 (.A1(N10084), .A2(n14278), .ZN(n38706));
    INVX1 U25835 (.I(N3917), .ZN(N38707));
    NANDX1 U25836 (.A1(N640), .A2(n16546), .ZN(N38708));
    INVX1 U25837 (.I(n24857), .ZN(n38709));
    INVX1 U25838 (.I(n15309), .ZN(N38710));
    NOR2X1 U25839 (.A1(n27758), .A2(n27425), .ZN(n38711));
    NANDX1 U25840 (.A1(n29169), .A2(n15518), .ZN(N38712));
    INVX1 U25841 (.I(N4595), .ZN(N38713));
    NANDX1 U25842 (.A1(n18019), .A2(N67), .ZN(N38714));
    INVX1 U25843 (.I(n27865), .ZN(N38715));
    NANDX1 U25844 (.A1(n22114), .A2(N6052), .ZN(n38716));
    NANDX1 U25845 (.A1(N8285), .A2(N1029), .ZN(N38717));
    NOR2X1 U25846 (.A1(n18369), .A2(n15306), .ZN(N38718));
    INVX1 U25847 (.I(N10846), .ZN(N38719));
    NANDX1 U25848 (.A1(n29016), .A2(n27391), .ZN(N38720));
    NANDX1 U25849 (.A1(n23735), .A2(N9210), .ZN(N38721));
    INVX1 U25850 (.I(n24587), .ZN(N38722));
    NANDX1 U25851 (.A1(n20856), .A2(N12658), .ZN(N38723));
    NANDX1 U25852 (.A1(N6236), .A2(n29222), .ZN(n38724));
    INVX1 U25853 (.I(n21895), .ZN(N38725));
    INVX1 U25854 (.I(n17782), .ZN(N38726));
    NANDX1 U25855 (.A1(N3392), .A2(n28289), .ZN(n38727));
    NANDX1 U25856 (.A1(n28141), .A2(N7947), .ZN(N38728));
    NANDX1 U25857 (.A1(n29169), .A2(n27595), .ZN(n38729));
    NANDX1 U25858 (.A1(N2898), .A2(n25833), .ZN(N38730));
    INVX1 U25859 (.I(N5780), .ZN(N38731));
    NOR2X1 U25860 (.A1(n20406), .A2(n25479), .ZN(n38732));
    NOR2X1 U25861 (.A1(n18177), .A2(n18910), .ZN(N38733));
    NANDX1 U25862 (.A1(n13568), .A2(N9628), .ZN(N38734));
    INVX1 U25863 (.I(n26688), .ZN(n38735));
    NANDX1 U25864 (.A1(N8880), .A2(n14266), .ZN(N38736));
    NOR2X1 U25865 (.A1(n14544), .A2(n20609), .ZN(N38737));
    NANDX1 U25866 (.A1(N6496), .A2(n18760), .ZN(n38738));
    INVX1 U25867 (.I(N4500), .ZN(N38739));
    NOR2X1 U25868 (.A1(n15208), .A2(n22229), .ZN(N38740));
    NOR2X1 U25869 (.A1(n27514), .A2(n25127), .ZN(N38741));
    NOR2X1 U25870 (.A1(n20529), .A2(n19467), .ZN(n38742));
    INVX1 U25871 (.I(n29496), .ZN(n38743));
    NANDX1 U25872 (.A1(N5682), .A2(n17535), .ZN(N38744));
    NOR2X1 U25873 (.A1(n25698), .A2(n19663), .ZN(n38745));
    NOR2X1 U25874 (.A1(N5356), .A2(n16213), .ZN(N38746));
    NANDX1 U25875 (.A1(n14235), .A2(n19040), .ZN(N38747));
    INVX1 U25876 (.I(n28779), .ZN(n38748));
    INVX1 U25877 (.I(N10931), .ZN(N38749));
    INVX1 U25878 (.I(n16831), .ZN(N38750));
    INVX1 U25879 (.I(n28334), .ZN(N38751));
    NANDX1 U25880 (.A1(N5831), .A2(n20426), .ZN(n38752));
    NANDX1 U25881 (.A1(n21905), .A2(N3976), .ZN(N38753));
    NOR2X1 U25882 (.A1(N12297), .A2(N12003), .ZN(n38754));
    NOR2X1 U25883 (.A1(N216), .A2(n15372), .ZN(N38755));
    NANDX1 U25884 (.A1(N6311), .A2(n26212), .ZN(N38756));
    NOR2X1 U25885 (.A1(n14534), .A2(n16542), .ZN(N38757));
    NANDX1 U25886 (.A1(n19307), .A2(n29994), .ZN(N38758));
    INVX1 U25887 (.I(N8209), .ZN(N38759));
    INVX1 U25888 (.I(n18512), .ZN(n38760));
    NANDX1 U25889 (.A1(N8981), .A2(N12209), .ZN(N38761));
    NANDX1 U25890 (.A1(n18302), .A2(n29104), .ZN(N38762));
    INVX1 U25891 (.I(n24132), .ZN(n38763));
    NOR2X1 U25892 (.A1(n16878), .A2(n15900), .ZN(N38764));
    INVX1 U25893 (.I(n17104), .ZN(N38765));
    NOR2X1 U25894 (.A1(N12491), .A2(n27582), .ZN(N38766));
    INVX1 U25895 (.I(n27863), .ZN(N38767));
    NOR2X1 U25896 (.A1(N11843), .A2(n23937), .ZN(N38768));
    INVX1 U25897 (.I(n14937), .ZN(N38769));
    INVX1 U25898 (.I(N8081), .ZN(N38770));
    NANDX1 U25899 (.A1(n17456), .A2(n27951), .ZN(N38771));
    NOR2X1 U25900 (.A1(n15506), .A2(N4886), .ZN(N38772));
    INVX1 U25901 (.I(n13047), .ZN(n38773));
    NANDX1 U25902 (.A1(N128), .A2(N1212), .ZN(n38774));
    NOR2X1 U25903 (.A1(n13760), .A2(n13904), .ZN(N38775));
    NANDX1 U25904 (.A1(n19198), .A2(n29803), .ZN(N38776));
    NANDX1 U25905 (.A1(n24862), .A2(N4983), .ZN(n38777));
    NANDX1 U25906 (.A1(N10867), .A2(N10515), .ZN(N38778));
    NANDX1 U25907 (.A1(n13031), .A2(N10918), .ZN(N38779));
    INVX1 U25908 (.I(n15476), .ZN(N38780));
    NANDX1 U25909 (.A1(n23236), .A2(n23557), .ZN(N38781));
    INVX1 U25910 (.I(N10554), .ZN(N38782));
    NOR2X1 U25911 (.A1(N698), .A2(n14620), .ZN(n38783));
    NOR2X1 U25912 (.A1(N7852), .A2(n16228), .ZN(N38784));
    NANDX1 U25913 (.A1(n26678), .A2(N6000), .ZN(N38785));
    INVX1 U25914 (.I(N10300), .ZN(N38786));
    INVX1 U25915 (.I(n14788), .ZN(n38787));
    INVX1 U25916 (.I(N8130), .ZN(N38788));
    INVX1 U25917 (.I(N12782), .ZN(n38789));
    NOR2X1 U25918 (.A1(N11824), .A2(n23648), .ZN(n38790));
    NANDX1 U25919 (.A1(n23662), .A2(N6541), .ZN(N38791));
    INVX1 U25920 (.I(n17859), .ZN(N38792));
    NOR2X1 U25921 (.A1(n26081), .A2(n29656), .ZN(N38793));
    NOR2X1 U25922 (.A1(n14464), .A2(n28770), .ZN(N38794));
    NANDX1 U25923 (.A1(n15161), .A2(N1814), .ZN(N38795));
    NANDX1 U25924 (.A1(N11573), .A2(n18041), .ZN(N38796));
    INVX1 U25925 (.I(N8113), .ZN(n38797));
    NANDX1 U25926 (.A1(n17111), .A2(N6973), .ZN(N38798));
    NANDX1 U25927 (.A1(N1761), .A2(n25030), .ZN(n38799));
    NANDX1 U25928 (.A1(n18170), .A2(N7674), .ZN(n38800));
    NOR2X1 U25929 (.A1(n18555), .A2(n19882), .ZN(N38801));
    INVX1 U25930 (.I(N12079), .ZN(N38802));
    INVX1 U25931 (.I(n13142), .ZN(N38803));
    NANDX1 U25932 (.A1(n25561), .A2(N9085), .ZN(n38804));
    NOR2X1 U25933 (.A1(n18118), .A2(n23548), .ZN(N38805));
    NANDX1 U25934 (.A1(N9166), .A2(n27269), .ZN(N38806));
    INVX1 U25935 (.I(N3592), .ZN(n38807));
    NOR2X1 U25936 (.A1(n13624), .A2(N7049), .ZN(N38808));
    NOR2X1 U25937 (.A1(n26224), .A2(N12721), .ZN(n38809));
    NOR2X1 U25938 (.A1(n17150), .A2(N3042), .ZN(n38810));
    NOR2X1 U25939 (.A1(n16206), .A2(n21212), .ZN(n38811));
    NANDX1 U25940 (.A1(n16934), .A2(N9629), .ZN(N38812));
    INVX1 U25941 (.I(n18410), .ZN(N38813));
    NOR2X1 U25942 (.A1(N8205), .A2(N1414), .ZN(n38814));
    NANDX1 U25943 (.A1(n22326), .A2(n29197), .ZN(N38815));
    NANDX1 U25944 (.A1(N10306), .A2(N11168), .ZN(n38816));
    INVX1 U25945 (.I(N8033), .ZN(N38817));
    NANDX1 U25946 (.A1(n13256), .A2(N11624), .ZN(n38818));
    NANDX1 U25947 (.A1(n15440), .A2(n18672), .ZN(N38819));
    INVX1 U25948 (.I(N87), .ZN(n38820));
    INVX1 U25949 (.I(N11853), .ZN(N38821));
    NANDX1 U25950 (.A1(n22995), .A2(N7657), .ZN(n38822));
    NOR2X1 U25951 (.A1(n14069), .A2(n29832), .ZN(N38823));
    NOR2X1 U25952 (.A1(N12258), .A2(N11614), .ZN(n38824));
    NANDX1 U25953 (.A1(n22525), .A2(N8380), .ZN(n38825));
    NOR2X1 U25954 (.A1(n28411), .A2(N568), .ZN(N38826));
    NANDX1 U25955 (.A1(n22176), .A2(N10874), .ZN(N38827));
    INVX1 U25956 (.I(n28409), .ZN(n38828));
    INVX1 U25957 (.I(N12829), .ZN(N38829));
    INVX1 U25958 (.I(n19090), .ZN(N38830));
    INVX1 U25959 (.I(n15527), .ZN(n38831));
    NOR2X1 U25960 (.A1(n29335), .A2(N4174), .ZN(N38832));
    INVX1 U25961 (.I(N11050), .ZN(n38833));
    NANDX1 U25962 (.A1(N8995), .A2(N7267), .ZN(N38834));
    INVX1 U25963 (.I(N11624), .ZN(N38835));
    NANDX1 U25964 (.A1(n29331), .A2(n23881), .ZN(N38836));
    NANDX1 U25965 (.A1(N3522), .A2(N4829), .ZN(n38837));
    NOR2X1 U25966 (.A1(N9264), .A2(N3102), .ZN(N38838));
    NANDX1 U25967 (.A1(n14065), .A2(n13839), .ZN(n38839));
    NOR2X1 U25968 (.A1(n18595), .A2(N12110), .ZN(N38840));
    INVX1 U25969 (.I(N1286), .ZN(N38841));
    INVX1 U25970 (.I(n23373), .ZN(N38842));
    INVX1 U25971 (.I(N4846), .ZN(n38843));
    INVX1 U25972 (.I(N7437), .ZN(N38844));
    INVX1 U25973 (.I(n24256), .ZN(N38845));
    INVX1 U25974 (.I(N7551), .ZN(n38846));
    NANDX1 U25975 (.A1(N2875), .A2(n28083), .ZN(n38847));
    NOR2X1 U25976 (.A1(N9835), .A2(n27276), .ZN(n38848));
    INVX1 U25977 (.I(n28409), .ZN(N38849));
    INVX1 U25978 (.I(N1868), .ZN(N38850));
    INVX1 U25979 (.I(n28622), .ZN(N38851));
    NANDX1 U25980 (.A1(N11170), .A2(N1111), .ZN(n38852));
    NANDX1 U25981 (.A1(N7987), .A2(n19705), .ZN(N38853));
    NANDX1 U25982 (.A1(N832), .A2(N9551), .ZN(n38854));
    NANDX1 U25983 (.A1(N12765), .A2(n17790), .ZN(n38855));
    NANDX1 U25984 (.A1(n20883), .A2(n13787), .ZN(N38856));
    NOR2X1 U25985 (.A1(n15001), .A2(N9395), .ZN(N38857));
    NANDX1 U25986 (.A1(N6674), .A2(N12269), .ZN(N38858));
    NOR2X1 U25987 (.A1(n21409), .A2(n22103), .ZN(N38859));
    NANDX1 U25988 (.A1(n18448), .A2(N8936), .ZN(n38860));
    NANDX1 U25989 (.A1(N8876), .A2(n22721), .ZN(n38861));
    NANDX1 U25990 (.A1(n13845), .A2(N3753), .ZN(N38862));
    NOR2X1 U25991 (.A1(n21212), .A2(N301), .ZN(n38863));
    INVX1 U25992 (.I(n17811), .ZN(n38864));
    NOR2X1 U25993 (.A1(N9048), .A2(n26607), .ZN(N38865));
    NOR2X1 U25994 (.A1(n15399), .A2(N10112), .ZN(n38866));
    INVX1 U25995 (.I(n29185), .ZN(N38867));
    NOR2X1 U25996 (.A1(N8203), .A2(n27140), .ZN(N38868));
    NOR2X1 U25997 (.A1(n14877), .A2(N9271), .ZN(N38869));
    NANDX1 U25998 (.A1(n24846), .A2(n19935), .ZN(N38870));
    NOR2X1 U25999 (.A1(N1718), .A2(n28870), .ZN(n38871));
    NANDX1 U26000 (.A1(N10593), .A2(n21453), .ZN(n38872));
    INVX1 U26001 (.I(n12998), .ZN(n38873));
    INVX1 U26002 (.I(n28050), .ZN(N38874));
    NANDX1 U26003 (.A1(N2628), .A2(n27547), .ZN(n38875));
    NANDX1 U26004 (.A1(n22457), .A2(n25155), .ZN(N38876));
    NANDX1 U26005 (.A1(n13474), .A2(n29114), .ZN(N38877));
    NANDX1 U26006 (.A1(N6676), .A2(n28162), .ZN(n38878));
    NANDX1 U26007 (.A1(N3440), .A2(n25164), .ZN(n38879));
    INVX1 U26008 (.I(N6877), .ZN(N38880));
    NANDX1 U26009 (.A1(n17813), .A2(n20283), .ZN(n38881));
    INVX1 U26010 (.I(N5338), .ZN(N38882));
    INVX1 U26011 (.I(N86), .ZN(N38883));
    NANDX1 U26012 (.A1(n21154), .A2(N10099), .ZN(N38884));
    NOR2X1 U26013 (.A1(n22712), .A2(n23865), .ZN(N38885));
    NOR2X1 U26014 (.A1(n15345), .A2(n15053), .ZN(N38886));
    INVX1 U26015 (.I(n14350), .ZN(N38887));
    NOR2X1 U26016 (.A1(N7475), .A2(N9824), .ZN(N38888));
    NANDX1 U26017 (.A1(N6452), .A2(N3970), .ZN(N38889));
    NOR2X1 U26018 (.A1(n23174), .A2(N8009), .ZN(N38890));
    NOR2X1 U26019 (.A1(N6761), .A2(N10577), .ZN(N38891));
    NANDX1 U26020 (.A1(n29756), .A2(n28389), .ZN(N38892));
    INVX1 U26021 (.I(N972), .ZN(N38893));
    NOR2X1 U26022 (.A1(n27103), .A2(N1057), .ZN(n38894));
    NANDX1 U26023 (.A1(N6680), .A2(N11156), .ZN(N38895));
    INVX1 U26024 (.I(n29392), .ZN(n38896));
    NANDX1 U26025 (.A1(n20272), .A2(N3160), .ZN(N38897));
    NOR2X1 U26026 (.A1(N2592), .A2(N6070), .ZN(N38898));
    NOR2X1 U26027 (.A1(N10067), .A2(N4454), .ZN(n38899));
    INVX1 U26028 (.I(n16518), .ZN(n38900));
    NOR2X1 U26029 (.A1(N7039), .A2(n28252), .ZN(N38901));
    NOR2X1 U26030 (.A1(n15120), .A2(N4875), .ZN(n38902));
    NOR2X1 U26031 (.A1(n30078), .A2(N4494), .ZN(N38903));
    NOR2X1 U26032 (.A1(N5044), .A2(n24163), .ZN(N38904));
    NOR2X1 U26033 (.A1(n20707), .A2(n25220), .ZN(N38905));
    NANDX1 U26034 (.A1(n27387), .A2(n24936), .ZN(N38906));
    INVX1 U26035 (.I(n15202), .ZN(N38907));
    INVX1 U26036 (.I(n18451), .ZN(n38908));
    NANDX1 U26037 (.A1(n15436), .A2(n21043), .ZN(n38909));
    NOR2X1 U26038 (.A1(N8426), .A2(N972), .ZN(N38910));
    NOR2X1 U26039 (.A1(n29519), .A2(N6050), .ZN(N38911));
    INVX1 U26040 (.I(N6420), .ZN(n38912));
    INVX1 U26041 (.I(n19421), .ZN(N38913));
    NANDX1 U26042 (.A1(n27736), .A2(n23550), .ZN(N38914));
    NANDX1 U26043 (.A1(n20790), .A2(n25930), .ZN(N38915));
    NANDX1 U26044 (.A1(n14816), .A2(N9021), .ZN(N38916));
    INVX1 U26045 (.I(n28596), .ZN(N38917));
    NANDX1 U26046 (.A1(N2902), .A2(n23394), .ZN(N38918));
    NANDX1 U26047 (.A1(n18103), .A2(N196), .ZN(N38919));
    NOR2X1 U26048 (.A1(n25025), .A2(N4193), .ZN(N38920));
    INVX1 U26049 (.I(N7879), .ZN(N38921));
    INVX1 U26050 (.I(N3223), .ZN(N38922));
    INVX1 U26051 (.I(N560), .ZN(N38923));
    NOR2X1 U26052 (.A1(n28312), .A2(N6980), .ZN(N38924));
    INVX1 U26053 (.I(N6156), .ZN(N38925));
    INVX1 U26054 (.I(n18293), .ZN(N38926));
    NOR2X1 U26055 (.A1(N8422), .A2(N8945), .ZN(n38927));
    NOR2X1 U26056 (.A1(n23505), .A2(N12321), .ZN(N38928));
    NANDX1 U26057 (.A1(n29157), .A2(N10779), .ZN(n38929));
    NOR2X1 U26058 (.A1(n20620), .A2(N4035), .ZN(n38930));
    NANDX1 U26059 (.A1(n27283), .A2(n22929), .ZN(N38931));
    NANDX1 U26060 (.A1(n22170), .A2(n27121), .ZN(N38932));
    NANDX1 U26061 (.A1(n18609), .A2(n28299), .ZN(N38933));
    INVX1 U26062 (.I(N2356), .ZN(N38934));
    NANDX1 U26063 (.A1(N2467), .A2(n19228), .ZN(n38935));
    INVX1 U26064 (.I(N11722), .ZN(n38936));
    NOR2X1 U26065 (.A1(N11340), .A2(n18575), .ZN(N38937));
    NOR2X1 U26066 (.A1(N8322), .A2(n16080), .ZN(N38938));
    NOR2X1 U26067 (.A1(n20387), .A2(n28401), .ZN(N38939));
    NANDX1 U26068 (.A1(N7968), .A2(N9042), .ZN(N38940));
    INVX1 U26069 (.I(n28587), .ZN(N38941));
    INVX1 U26070 (.I(n21941), .ZN(n38942));
    INVX1 U26071 (.I(n13127), .ZN(n38943));
    NANDX1 U26072 (.A1(N6326), .A2(N10110), .ZN(N38944));
    INVX1 U26073 (.I(n24934), .ZN(n38945));
    INVX1 U26074 (.I(N1189), .ZN(N38946));
    INVX1 U26075 (.I(n14250), .ZN(N38947));
    INVX1 U26076 (.I(n23639), .ZN(n38948));
    INVX1 U26077 (.I(n22636), .ZN(N38949));
    INVX1 U26078 (.I(N8411), .ZN(N38950));
    NOR2X1 U26079 (.A1(n20957), .A2(N5294), .ZN(N38951));
    NANDX1 U26080 (.A1(N6951), .A2(n25680), .ZN(N38952));
    INVX1 U26081 (.I(n23282), .ZN(N38953));
    NANDX1 U26082 (.A1(N11579), .A2(n15832), .ZN(N38954));
    NOR2X1 U26083 (.A1(N1777), .A2(N7635), .ZN(n38955));
    INVX1 U26084 (.I(n14903), .ZN(N38956));
    NANDX1 U26085 (.A1(N11138), .A2(n13573), .ZN(N38957));
    INVX1 U26086 (.I(N5934), .ZN(n38958));
    NANDX1 U26087 (.A1(n15039), .A2(N10345), .ZN(n38959));
    INVX1 U26088 (.I(N7255), .ZN(N38960));
    INVX1 U26089 (.I(n21724), .ZN(N38961));
    INVX1 U26090 (.I(n29989), .ZN(N38962));
    INVX1 U26091 (.I(n29523), .ZN(n38963));
    INVX1 U26092 (.I(n23989), .ZN(N38964));
    NOR2X1 U26093 (.A1(n16319), .A2(N8092), .ZN(n38965));
    NOR2X1 U26094 (.A1(n28161), .A2(N163), .ZN(N38966));
    NANDX1 U26095 (.A1(n13856), .A2(n20819), .ZN(N38967));
    NANDX1 U26096 (.A1(n21490), .A2(n25631), .ZN(N38968));
    NOR2X1 U26097 (.A1(N1390), .A2(N6631), .ZN(n38969));
    INVX1 U26098 (.I(n26679), .ZN(N38970));
    INVX1 U26099 (.I(N5412), .ZN(N38971));
    NOR2X1 U26100 (.A1(N31), .A2(n30065), .ZN(N38972));
    NOR2X1 U26101 (.A1(n22574), .A2(n21651), .ZN(n38973));
    INVX1 U26102 (.I(n22425), .ZN(N38974));
    NOR2X1 U26103 (.A1(N2354), .A2(N1656), .ZN(n38975));
    INVX1 U26104 (.I(N6013), .ZN(N38976));
    NANDX1 U26105 (.A1(N713), .A2(n23647), .ZN(N38977));
    INVX1 U26106 (.I(n19573), .ZN(n38978));
    NOR2X1 U26107 (.A1(N6975), .A2(N10254), .ZN(n38979));
    INVX1 U26108 (.I(n17026), .ZN(N38980));
    INVX1 U26109 (.I(n19529), .ZN(n38981));
    NOR2X1 U26110 (.A1(N939), .A2(n14537), .ZN(n38982));
    NOR2X1 U26111 (.A1(n20762), .A2(n19949), .ZN(n38983));
    NANDX1 U26112 (.A1(n20792), .A2(N8437), .ZN(N38984));
    NANDX1 U26113 (.A1(N1789), .A2(n30087), .ZN(n38985));
    NOR2X1 U26114 (.A1(n24213), .A2(n28857), .ZN(N38986));
    NANDX1 U26115 (.A1(n14430), .A2(n21477), .ZN(N38987));
    NANDX1 U26116 (.A1(N9526), .A2(N10750), .ZN(n38988));
    NANDX1 U26117 (.A1(N2645), .A2(N185), .ZN(n38989));
    INVX1 U26118 (.I(n28318), .ZN(N38990));
    INVX1 U26119 (.I(n19513), .ZN(n38991));
    NANDX1 U26120 (.A1(n23445), .A2(N8904), .ZN(n38992));
    NANDX1 U26121 (.A1(n12944), .A2(n23440), .ZN(N38993));
    INVX1 U26122 (.I(N3569), .ZN(N38994));
    NOR2X1 U26123 (.A1(n17914), .A2(n12921), .ZN(n38995));
    NOR2X1 U26124 (.A1(N6088), .A2(n14710), .ZN(n38996));
    NOR2X1 U26125 (.A1(N8668), .A2(n27483), .ZN(n38997));
    NANDX1 U26126 (.A1(n13601), .A2(N336), .ZN(n38998));
    NANDX1 U26127 (.A1(n24546), .A2(N9861), .ZN(N38999));
    NANDX1 U26128 (.A1(n17561), .A2(N1067), .ZN(N39000));
    NANDX1 U26129 (.A1(n29119), .A2(n29384), .ZN(N39001));
    NOR2X1 U26130 (.A1(n18494), .A2(N3013), .ZN(N39002));
    INVX1 U26131 (.I(n15958), .ZN(N39003));
    INVX1 U26132 (.I(n19519), .ZN(n39004));
    INVX1 U26133 (.I(N9313), .ZN(N39005));
    INVX1 U26134 (.I(N11072), .ZN(n39006));
    NANDX1 U26135 (.A1(n13129), .A2(N9880), .ZN(N39007));
    INVX1 U26136 (.I(n27838), .ZN(N39008));
    NOR2X1 U26137 (.A1(N404), .A2(n13745), .ZN(n39009));
    INVX1 U26138 (.I(N2565), .ZN(N39010));
    NANDX1 U26139 (.A1(N2191), .A2(n27110), .ZN(N39011));
    NANDX1 U26140 (.A1(N9016), .A2(N3095), .ZN(n39012));
    NANDX1 U26141 (.A1(N4586), .A2(n20774), .ZN(n39013));
    NOR2X1 U26142 (.A1(n17854), .A2(N9130), .ZN(N39014));
    NANDX1 U26143 (.A1(n24428), .A2(n25087), .ZN(n39015));
    NOR2X1 U26144 (.A1(N2370), .A2(n22907), .ZN(N39016));
    INVX1 U26145 (.I(N2578), .ZN(N39017));
    NANDX1 U26146 (.A1(n13101), .A2(n15707), .ZN(n39018));
    NOR2X1 U26147 (.A1(n23536), .A2(N1968), .ZN(N39019));
    NANDX1 U26148 (.A1(N12500), .A2(n15712), .ZN(N39020));
    INVX1 U26149 (.I(n15065), .ZN(N39021));
    NANDX1 U26150 (.A1(N7785), .A2(N598), .ZN(n39022));
    NOR2X1 U26151 (.A1(N5361), .A2(n22390), .ZN(N39023));
    NANDX1 U26152 (.A1(n28644), .A2(n13026), .ZN(N39024));
    INVX1 U26153 (.I(n16360), .ZN(N39025));
    NOR2X1 U26154 (.A1(n20044), .A2(N10651), .ZN(N39026));
    NOR2X1 U26155 (.A1(N8046), .A2(n13020), .ZN(n39027));
    INVX1 U26156 (.I(N5360), .ZN(N39028));
    INVX1 U26157 (.I(N9534), .ZN(N39029));
    INVX1 U26158 (.I(n19865), .ZN(N39030));
    NANDX1 U26159 (.A1(N419), .A2(n21832), .ZN(N39031));
    INVX1 U26160 (.I(N1480), .ZN(n39032));
    NANDX1 U26161 (.A1(n28328), .A2(n16544), .ZN(N39033));
    NOR2X1 U26162 (.A1(n24673), .A2(N5702), .ZN(N39034));
    NOR2X1 U26163 (.A1(n30033), .A2(n28092), .ZN(N39035));
    INVX1 U26164 (.I(n17100), .ZN(N39036));
    INVX1 U26165 (.I(N321), .ZN(N39037));
    INVX1 U26166 (.I(n21696), .ZN(N39038));
    INVX1 U26167 (.I(n13973), .ZN(n39039));
    NANDX1 U26168 (.A1(n16970), .A2(n15553), .ZN(n39040));
    NOR2X1 U26169 (.A1(N10890), .A2(n19711), .ZN(N39041));
    NOR2X1 U26170 (.A1(n17910), .A2(n28136), .ZN(N39042));
    NANDX1 U26171 (.A1(N6890), .A2(n19831), .ZN(N39043));
    NANDX1 U26172 (.A1(N8369), .A2(n27237), .ZN(N39044));
    NOR2X1 U26173 (.A1(n13473), .A2(n22858), .ZN(N39045));
    NANDX1 U26174 (.A1(N7735), .A2(N11936), .ZN(N39046));
    NOR2X1 U26175 (.A1(N5689), .A2(n15297), .ZN(N39047));
    NANDX1 U26176 (.A1(N5230), .A2(N4178), .ZN(N39048));
    NANDX1 U26177 (.A1(n15486), .A2(n24541), .ZN(N39049));
    NOR2X1 U26178 (.A1(n19967), .A2(n30071), .ZN(N39050));
    INVX1 U26179 (.I(n22883), .ZN(N39051));
    NANDX1 U26180 (.A1(n29201), .A2(n23893), .ZN(n39052));
    INVX1 U26181 (.I(n27199), .ZN(N39053));
    NOR2X1 U26182 (.A1(n24182), .A2(N5453), .ZN(N39054));
    NOR2X1 U26183 (.A1(n21111), .A2(N2552), .ZN(N39055));
    NOR2X1 U26184 (.A1(n23144), .A2(n13970), .ZN(n39056));
    NANDX1 U26185 (.A1(N742), .A2(n14466), .ZN(N39057));
    INVX1 U26186 (.I(N6430), .ZN(n39058));
    NANDX1 U26187 (.A1(n21656), .A2(N220), .ZN(N39059));
    NANDX1 U26188 (.A1(n24499), .A2(N4266), .ZN(N39060));
    NOR2X1 U26189 (.A1(N11177), .A2(n24233), .ZN(N39061));
    NOR2X1 U26190 (.A1(n20667), .A2(n16978), .ZN(N39062));
    INVX1 U26191 (.I(n19730), .ZN(N39063));
    NOR2X1 U26192 (.A1(n14814), .A2(n16791), .ZN(N39064));
    NANDX1 U26193 (.A1(n27556), .A2(N10805), .ZN(N39065));
    NANDX1 U26194 (.A1(N7091), .A2(n13356), .ZN(N39066));
    NANDX1 U26195 (.A1(N97), .A2(n15887), .ZN(n39067));
    NOR2X1 U26196 (.A1(N838), .A2(N215), .ZN(N39068));
    NOR2X1 U26197 (.A1(n25966), .A2(n29977), .ZN(N39069));
    NOR2X1 U26198 (.A1(n14746), .A2(n22339), .ZN(N39070));
    NOR2X1 U26199 (.A1(n19012), .A2(n27803), .ZN(N39071));
    NOR2X1 U26200 (.A1(n13107), .A2(n14501), .ZN(n39072));
    INVX1 U26201 (.I(n18645), .ZN(N39073));
    NANDX1 U26202 (.A1(n18393), .A2(n17938), .ZN(N39074));
    INVX1 U26203 (.I(n23744), .ZN(n39075));
    NANDX1 U26204 (.A1(n20073), .A2(N4411), .ZN(N39076));
    INVX1 U26205 (.I(n27163), .ZN(N39077));
    NANDX1 U26206 (.A1(n13791), .A2(n15821), .ZN(N39078));
    NOR2X1 U26207 (.A1(N6914), .A2(N5219), .ZN(N39079));
    INVX1 U26208 (.I(n29430), .ZN(n39080));
    NOR2X1 U26209 (.A1(N10828), .A2(n13328), .ZN(N39081));
    NOR2X1 U26210 (.A1(N3030), .A2(n21725), .ZN(N39082));
    INVX1 U26211 (.I(n19393), .ZN(n39083));
    NOR2X1 U26212 (.A1(n13593), .A2(N3756), .ZN(N39084));
    INVX1 U26213 (.I(N2100), .ZN(n39085));
    INVX1 U26214 (.I(n16777), .ZN(N39086));
    INVX1 U26215 (.I(n15553), .ZN(n39087));
    NANDX1 U26216 (.A1(N9529), .A2(n24187), .ZN(n39088));
    NOR2X1 U26217 (.A1(n16894), .A2(N9773), .ZN(N39089));
    INVX1 U26218 (.I(n19245), .ZN(N39090));
    NANDX1 U26219 (.A1(N1758), .A2(n14719), .ZN(N39091));
    NOR2X1 U26220 (.A1(n24185), .A2(n14012), .ZN(N39092));
    NOR2X1 U26221 (.A1(n23574), .A2(n15900), .ZN(N39093));
    NOR2X1 U26222 (.A1(n15164), .A2(n26185), .ZN(n39094));
    NOR2X1 U26223 (.A1(N4419), .A2(n14467), .ZN(n39095));
    NOR2X1 U26224 (.A1(n26872), .A2(N12851), .ZN(n39096));
    INVX1 U26225 (.I(n19771), .ZN(N39097));
    INVX1 U26226 (.I(n15229), .ZN(N39098));
    NOR2X1 U26227 (.A1(n17132), .A2(n24758), .ZN(n39099));
    INVX1 U26228 (.I(n20486), .ZN(n39100));
    NANDX1 U26229 (.A1(n16267), .A2(N30), .ZN(N39101));
    INVX1 U26230 (.I(N11722), .ZN(N39102));
    NOR2X1 U26231 (.A1(N3901), .A2(N957), .ZN(N39103));
    NOR2X1 U26232 (.A1(N6473), .A2(n28635), .ZN(N39104));
    NANDX1 U26233 (.A1(n22373), .A2(N391), .ZN(N39105));
    NOR2X1 U26234 (.A1(N6981), .A2(n14210), .ZN(N39106));
    NOR2X1 U26235 (.A1(n21448), .A2(N44), .ZN(N39107));
    NOR2X1 U26236 (.A1(n22859), .A2(n18115), .ZN(N39108));
    INVX1 U26237 (.I(N10910), .ZN(N39109));
    INVX1 U26238 (.I(N3483), .ZN(N39110));
    NOR2X1 U26239 (.A1(n16524), .A2(N9977), .ZN(N39111));
    NOR2X1 U26240 (.A1(n16599), .A2(n26243), .ZN(N39112));
    NANDX1 U26241 (.A1(N5781), .A2(n26525), .ZN(n39113));
    NANDX1 U26242 (.A1(n28379), .A2(n27482), .ZN(n39114));
    INVX1 U26243 (.I(N4715), .ZN(n39115));
    NANDX1 U26244 (.A1(n15645), .A2(n15648), .ZN(n39116));
    NOR2X1 U26245 (.A1(n27336), .A2(N11189), .ZN(N39117));
    NANDX1 U26246 (.A1(N1870), .A2(N2499), .ZN(n39118));
    INVX1 U26247 (.I(n14714), .ZN(N39119));
    INVX1 U26248 (.I(N5721), .ZN(n39120));
    NOR2X1 U26249 (.A1(N6130), .A2(n27624), .ZN(n39121));
    NOR2X1 U26250 (.A1(n22731), .A2(n14011), .ZN(N39122));
    INVX1 U26251 (.I(n29680), .ZN(N39123));
    NOR2X1 U26252 (.A1(N3876), .A2(n25219), .ZN(N39124));
    NANDX1 U26253 (.A1(N264), .A2(N11105), .ZN(N39125));
    NOR2X1 U26254 (.A1(n16306), .A2(N83), .ZN(N39126));
    NOR2X1 U26255 (.A1(N708), .A2(N4288), .ZN(n39127));
    NANDX1 U26256 (.A1(n15637), .A2(n20185), .ZN(N39128));
    INVX1 U26257 (.I(N3200), .ZN(N39129));
    INVX1 U26258 (.I(N4224), .ZN(n39130));
    NANDX1 U26259 (.A1(n25328), .A2(n18142), .ZN(N39131));
    NOR2X1 U26260 (.A1(n19640), .A2(N12832), .ZN(N39132));
    INVX1 U26261 (.I(N5995), .ZN(N39133));
    NANDX1 U26262 (.A1(n26720), .A2(n13766), .ZN(N39134));
    INVX1 U26263 (.I(n15752), .ZN(N39135));
    NANDX1 U26264 (.A1(N7307), .A2(N10564), .ZN(N39136));
    NANDX1 U26265 (.A1(N6972), .A2(n22316), .ZN(N39137));
    INVX1 U26266 (.I(n25753), .ZN(n39138));
    INVX1 U26267 (.I(N599), .ZN(N39139));
    NANDX1 U26268 (.A1(n29318), .A2(n16236), .ZN(n39140));
    NOR2X1 U26269 (.A1(n19604), .A2(N7996), .ZN(n39141));
    INVX1 U26270 (.I(n23827), .ZN(N39142));
    NANDX1 U26271 (.A1(n25891), .A2(N393), .ZN(N39143));
    NANDX1 U26272 (.A1(N3954), .A2(n13224), .ZN(N39144));
    NOR2X1 U26273 (.A1(N9949), .A2(N7210), .ZN(n39145));
    NOR2X1 U26274 (.A1(N12275), .A2(N737), .ZN(n39146));
    NOR2X1 U26275 (.A1(n18476), .A2(n26742), .ZN(n39147));
    INVX1 U26276 (.I(n13502), .ZN(N39148));
    NANDX1 U26277 (.A1(N11672), .A2(n13393), .ZN(N39149));
    NANDX1 U26278 (.A1(N8876), .A2(n13992), .ZN(n39150));
    INVX1 U26279 (.I(n26754), .ZN(N39151));
    INVX1 U26280 (.I(N7741), .ZN(n39152));
    NOR2X1 U26281 (.A1(n26783), .A2(N8305), .ZN(N39153));
    NANDX1 U26282 (.A1(n25583), .A2(n22756), .ZN(N39154));
    INVX1 U26283 (.I(N9469), .ZN(N39155));
    NANDX1 U26284 (.A1(N12086), .A2(n17503), .ZN(N39156));
    NANDX1 U26285 (.A1(n19295), .A2(N10681), .ZN(N39157));
    NOR2X1 U26286 (.A1(n20032), .A2(n19611), .ZN(n39158));
    INVX1 U26287 (.I(n16636), .ZN(n39159));
    NANDX1 U26288 (.A1(n27893), .A2(N8772), .ZN(N39160));
    NOR2X1 U26289 (.A1(n29847), .A2(N7963), .ZN(N39161));
    NOR2X1 U26290 (.A1(n13701), .A2(N7056), .ZN(n39162));
    NOR2X1 U26291 (.A1(n21049), .A2(N3357), .ZN(N39163));
    NANDX1 U26292 (.A1(N6255), .A2(N222), .ZN(N39164));
    INVX1 U26293 (.I(N1700), .ZN(N39165));
    NANDX1 U26294 (.A1(n28242), .A2(N11168), .ZN(N39166));
    NOR2X1 U26295 (.A1(n28889), .A2(n17231), .ZN(n39167));
    NANDX1 U26296 (.A1(n18046), .A2(n27912), .ZN(N39168));
    INVX1 U26297 (.I(n26638), .ZN(N39169));
    NOR2X1 U26298 (.A1(n20758), .A2(N1697), .ZN(N39170));
    INVX1 U26299 (.I(N7075), .ZN(N39171));
    NOR2X1 U26300 (.A1(N12671), .A2(N6784), .ZN(N39172));
    INVX1 U26301 (.I(n19305), .ZN(N39173));
    NANDX1 U26302 (.A1(n14047), .A2(n22556), .ZN(n39174));
    NANDX1 U26303 (.A1(N5964), .A2(N11890), .ZN(N39175));
    NANDX1 U26304 (.A1(N6186), .A2(n29830), .ZN(N39176));
    INVX1 U26305 (.I(n17724), .ZN(N39177));
    NOR2X1 U26306 (.A1(n26335), .A2(N2956), .ZN(N39178));
    NANDX1 U26307 (.A1(n13428), .A2(n13406), .ZN(n39179));
    NOR2X1 U26308 (.A1(n29900), .A2(N8333), .ZN(n39180));
    NANDX1 U26309 (.A1(N5708), .A2(n29090), .ZN(N39181));
    INVX1 U26310 (.I(N9180), .ZN(N39182));
    NANDX1 U26311 (.A1(n19079), .A2(n21850), .ZN(n39183));
    NANDX1 U26312 (.A1(N7372), .A2(n29716), .ZN(N39184));
    INVX1 U26313 (.I(N9979), .ZN(N39185));
    INVX1 U26314 (.I(N6190), .ZN(N39186));
    INVX1 U26315 (.I(N11145), .ZN(N39187));
    NOR2X1 U26316 (.A1(n22128), .A2(n29536), .ZN(N39188));
    INVX1 U26317 (.I(n28412), .ZN(n39189));
    INVX1 U26318 (.I(N885), .ZN(N39190));
    INVX1 U26319 (.I(N8262), .ZN(n39191));
    NOR2X1 U26320 (.A1(n14635), .A2(n30114), .ZN(n39192));
    NOR2X1 U26321 (.A1(n22967), .A2(N6891), .ZN(n39193));
    NOR2X1 U26322 (.A1(N10480), .A2(n26941), .ZN(N39194));
    NOR2X1 U26323 (.A1(n23766), .A2(n15882), .ZN(N39195));
    NANDX1 U26324 (.A1(n13697), .A2(N11815), .ZN(N39196));
    INVX1 U26325 (.I(N1234), .ZN(N39197));
    NOR2X1 U26326 (.A1(n26767), .A2(N7423), .ZN(n39198));
    NOR2X1 U26327 (.A1(n26473), .A2(n27081), .ZN(n39199));
    NANDX1 U26328 (.A1(n25871), .A2(n13070), .ZN(N39200));
    NOR2X1 U26329 (.A1(n18886), .A2(n13955), .ZN(N39201));
    INVX1 U26330 (.I(n27147), .ZN(n39202));
    NANDX1 U26331 (.A1(N9545), .A2(n27123), .ZN(N39203));
    NANDX1 U26332 (.A1(n21072), .A2(n22575), .ZN(N39204));
    INVX1 U26333 (.I(n20113), .ZN(n39205));
    INVX1 U26334 (.I(n22451), .ZN(N39206));
    NOR2X1 U26335 (.A1(n23820), .A2(N8808), .ZN(n39207));
    NANDX1 U26336 (.A1(n24195), .A2(n24880), .ZN(N39208));
    INVX1 U26337 (.I(n15851), .ZN(N39209));
    NANDX1 U26338 (.A1(n13215), .A2(N12009), .ZN(n39210));
    NOR2X1 U26339 (.A1(n28856), .A2(n18856), .ZN(N39211));
    NOR2X1 U26340 (.A1(N11788), .A2(n23976), .ZN(n39212));
    INVX1 U26341 (.I(n14303), .ZN(N39213));
    NOR2X1 U26342 (.A1(n25291), .A2(n19691), .ZN(N39214));
    NANDX1 U26343 (.A1(n22277), .A2(n27715), .ZN(n39215));
    NOR2X1 U26344 (.A1(n14714), .A2(N2505), .ZN(N39216));
    NANDX1 U26345 (.A1(n22652), .A2(n24955), .ZN(N39217));
    NANDX1 U26346 (.A1(N4895), .A2(n22323), .ZN(N39218));
    NOR2X1 U26347 (.A1(n29090), .A2(N5626), .ZN(N39219));
    INVX1 U26348 (.I(N3364), .ZN(N39220));
    NOR2X1 U26349 (.A1(n16508), .A2(N3933), .ZN(n39221));
    NANDX1 U26350 (.A1(n15226), .A2(N11349), .ZN(N39222));
    NOR2X1 U26351 (.A1(n15574), .A2(N5188), .ZN(N39223));
    INVX1 U26352 (.I(n18438), .ZN(N39224));
    NANDX1 U26353 (.A1(n13356), .A2(n26689), .ZN(N39225));
    INVX1 U26354 (.I(n24193), .ZN(n39226));
    NOR2X1 U26355 (.A1(N156), .A2(n27467), .ZN(N39227));
    INVX1 U26356 (.I(n28194), .ZN(N39228));
    NOR2X1 U26357 (.A1(n28847), .A2(N9698), .ZN(N39229));
    NOR2X1 U26358 (.A1(n21033), .A2(N7200), .ZN(N39230));
    NOR2X1 U26359 (.A1(n26658), .A2(N10493), .ZN(n39231));
    INVX1 U26360 (.I(N777), .ZN(n39232));
    INVX1 U26361 (.I(n26943), .ZN(N39233));
    NOR2X1 U26362 (.A1(N649), .A2(N8154), .ZN(N39234));
    NANDX1 U26363 (.A1(N4783), .A2(N1902), .ZN(n39235));
    NOR2X1 U26364 (.A1(n23220), .A2(n14536), .ZN(N39236));
    INVX1 U26365 (.I(n19772), .ZN(n39237));
    INVX1 U26366 (.I(N4091), .ZN(N39238));
    NOR2X1 U26367 (.A1(n25619), .A2(N1420), .ZN(n39239));
    NOR2X1 U26368 (.A1(N12237), .A2(N9961), .ZN(n39240));
    INVX1 U26369 (.I(n21934), .ZN(N39241));
    NOR2X1 U26370 (.A1(N3217), .A2(n29133), .ZN(N39242));
    NANDX1 U26371 (.A1(n18435), .A2(N9488), .ZN(N39243));
    INVX1 U26372 (.I(N7773), .ZN(N39244));
    NANDX1 U26373 (.A1(N2584), .A2(N7771), .ZN(n39245));
    INVX1 U26374 (.I(n29435), .ZN(n39246));
    NOR2X1 U26375 (.A1(N342), .A2(n19898), .ZN(N39247));
    NANDX1 U26376 (.A1(N12122), .A2(N4296), .ZN(N39248));
    NOR2X1 U26377 (.A1(n20454), .A2(n29759), .ZN(N39249));
    NOR2X1 U26378 (.A1(N11476), .A2(n13802), .ZN(N39250));
    NOR2X1 U26379 (.A1(N6389), .A2(n26038), .ZN(N39251));
    NANDX1 U26380 (.A1(N12), .A2(n17834), .ZN(N39252));
    INVX1 U26381 (.I(n21926), .ZN(N39253));
    NOR2X1 U26382 (.A1(n29119), .A2(N10224), .ZN(n39254));
    INVX1 U26383 (.I(N4760), .ZN(N39255));
    NOR2X1 U26384 (.A1(n28487), .A2(n26041), .ZN(n39256));
    INVX1 U26385 (.I(N12606), .ZN(N39257));
    NOR2X1 U26386 (.A1(N576), .A2(N1508), .ZN(N39258));
    NOR2X1 U26387 (.A1(n13642), .A2(n13630), .ZN(n39259));
    NOR2X1 U26388 (.A1(n25305), .A2(N3946), .ZN(N39260));
    NOR2X1 U26389 (.A1(N10922), .A2(N3982), .ZN(N39261));
    INVX1 U26390 (.I(n28095), .ZN(N39262));
    NOR2X1 U26391 (.A1(n24536), .A2(N2213), .ZN(n39263));
    NOR2X1 U26392 (.A1(N794), .A2(n29865), .ZN(n39264));
    INVX1 U26393 (.I(n24882), .ZN(n39265));
    NOR2X1 U26394 (.A1(n19653), .A2(n28320), .ZN(n39266));
    INVX1 U26395 (.I(n26209), .ZN(N39267));
    NANDX1 U26396 (.A1(N6630), .A2(N10398), .ZN(N39268));
    NOR2X1 U26397 (.A1(n20528), .A2(N10973), .ZN(n39269));
    NOR2X1 U26398 (.A1(n24187), .A2(n13175), .ZN(N39270));
    INVX1 U26399 (.I(n20702), .ZN(N39271));
    INVX1 U26400 (.I(n24040), .ZN(N39272));
    INVX1 U26401 (.I(n19264), .ZN(N39273));
    INVX1 U26402 (.I(N3898), .ZN(N39274));
    INVX1 U26403 (.I(n26952), .ZN(n39275));
    NANDX1 U26404 (.A1(N7994), .A2(n25895), .ZN(n39276));
    INVX1 U26405 (.I(n26419), .ZN(N39277));
    NANDX1 U26406 (.A1(N1092), .A2(n13688), .ZN(N39278));
    NANDX1 U26407 (.A1(n29412), .A2(n24414), .ZN(n39279));
    INVX1 U26408 (.I(n14504), .ZN(n39280));
    INVX1 U26409 (.I(N8429), .ZN(N39281));
    NANDX1 U26410 (.A1(n21434), .A2(N7962), .ZN(n39282));
    NANDX1 U26411 (.A1(N4044), .A2(n21136), .ZN(N39283));
    NANDX1 U26412 (.A1(n13306), .A2(n18039), .ZN(N39284));
    NOR2X1 U26413 (.A1(n18704), .A2(N7165), .ZN(N39285));
    NANDX1 U26414 (.A1(N11162), .A2(N1507), .ZN(N39286));
    NANDX1 U26415 (.A1(n28156), .A2(n28199), .ZN(N39287));
    NOR2X1 U26416 (.A1(N4366), .A2(n24480), .ZN(n39288));
    NANDX1 U26417 (.A1(n24156), .A2(n26729), .ZN(N39289));
    INVX1 U26418 (.I(n23430), .ZN(N39290));
    INVX1 U26419 (.I(n28294), .ZN(N39291));
    INVX1 U26420 (.I(n21911), .ZN(n39292));
    NANDX1 U26421 (.A1(n27257), .A2(N1768), .ZN(N39293));
    INVX1 U26422 (.I(n15786), .ZN(N39294));
    NOR2X1 U26423 (.A1(N12804), .A2(n17149), .ZN(N39295));
    INVX1 U26424 (.I(N705), .ZN(n39296));
    INVX1 U26425 (.I(n26380), .ZN(N39297));
    INVX1 U26426 (.I(N1384), .ZN(N39298));
    NANDX1 U26427 (.A1(n16635), .A2(n28743), .ZN(N39299));
    INVX1 U26428 (.I(n14696), .ZN(n39300));
    NOR2X1 U26429 (.A1(N5608), .A2(N9039), .ZN(N39301));
    INVX1 U26430 (.I(n29763), .ZN(n39302));
    NOR2X1 U26431 (.A1(N4395), .A2(N11616), .ZN(N39303));
    NOR2X1 U26432 (.A1(N2551), .A2(N7973), .ZN(N39304));
    INVX1 U26433 (.I(n16395), .ZN(N39305));
    INVX1 U26434 (.I(N8735), .ZN(N39306));
    NOR2X1 U26435 (.A1(N9438), .A2(N3106), .ZN(n39307));
    INVX1 U26436 (.I(n15147), .ZN(N39308));
    INVX1 U26437 (.I(n21570), .ZN(n39309));
    NOR2X1 U26438 (.A1(n25723), .A2(N6561), .ZN(N39310));
    NANDX1 U26439 (.A1(N10249), .A2(n23195), .ZN(N39311));
    NANDX1 U26440 (.A1(n22930), .A2(N7754), .ZN(n39312));
    INVX1 U26441 (.I(n28537), .ZN(n39313));
    NOR2X1 U26442 (.A1(n19223), .A2(n16724), .ZN(n39314));
    NANDX1 U26443 (.A1(n23617), .A2(n28339), .ZN(n39315));
    INVX1 U26444 (.I(n14729), .ZN(N39316));
    NOR2X1 U26445 (.A1(N10266), .A2(N986), .ZN(n39317));
    NOR2X1 U26446 (.A1(n19000), .A2(N9047), .ZN(N39318));
    NANDX1 U26447 (.A1(N10667), .A2(n29912), .ZN(n39319));
    NANDX1 U26448 (.A1(n21448), .A2(n21344), .ZN(N39320));
    INVX1 U26449 (.I(N5594), .ZN(N39321));
    NOR2X1 U26450 (.A1(n19539), .A2(n15842), .ZN(N39322));
    NANDX1 U26451 (.A1(N12771), .A2(N8634), .ZN(n39323));
    INVX1 U26452 (.I(n16286), .ZN(N39324));
    NOR2X1 U26453 (.A1(n22627), .A2(N5371), .ZN(N39325));
    NANDX1 U26454 (.A1(n22169), .A2(n17549), .ZN(n39326));
    INVX1 U26455 (.I(N6769), .ZN(N39327));
    NOR2X1 U26456 (.A1(n23952), .A2(n17034), .ZN(N39328));
    NOR2X1 U26457 (.A1(N899), .A2(n24594), .ZN(N39329));
    NOR2X1 U26458 (.A1(N5982), .A2(N5123), .ZN(N39330));
    NANDX1 U26459 (.A1(n26211), .A2(n15132), .ZN(N39331));
    NOR2X1 U26460 (.A1(n20985), .A2(n20725), .ZN(N39332));
    NOR2X1 U26461 (.A1(n29084), .A2(n25128), .ZN(n39333));
    NOR2X1 U26462 (.A1(N11717), .A2(N3624), .ZN(N39334));
    NOR2X1 U26463 (.A1(n16563), .A2(n17916), .ZN(N39335));
    NOR2X1 U26464 (.A1(N10495), .A2(N96), .ZN(N39336));
    NOR2X1 U26465 (.A1(n28043), .A2(n17874), .ZN(N39337));
    NANDX1 U26466 (.A1(N45), .A2(N249), .ZN(N39338));
    NOR2X1 U26467 (.A1(n21867), .A2(n19845), .ZN(N39339));
    NANDX1 U26468 (.A1(n22598), .A2(n25826), .ZN(N39340));
    NOR2X1 U26469 (.A1(n23104), .A2(N10460), .ZN(n39341));
    NANDX1 U26470 (.A1(N3376), .A2(N1308), .ZN(N39342));
    NOR2X1 U26471 (.A1(N11552), .A2(n18952), .ZN(n39343));
    NOR2X1 U26472 (.A1(n17810), .A2(n19230), .ZN(n39344));
    INVX1 U26473 (.I(n22644), .ZN(N39345));
    NANDX1 U26474 (.A1(n26624), .A2(N8529), .ZN(n39346));
    NOR2X1 U26475 (.A1(n15280), .A2(n16583), .ZN(N39347));
    NANDX1 U26476 (.A1(N3016), .A2(N1267), .ZN(N39348));
    NOR2X1 U26477 (.A1(N3264), .A2(N10244), .ZN(n39349));
    INVX1 U26478 (.I(N11670), .ZN(n39350));
    NOR2X1 U26479 (.A1(N12806), .A2(N7358), .ZN(N39351));
    NOR2X1 U26480 (.A1(N5772), .A2(n17818), .ZN(N39352));
    NOR2X1 U26481 (.A1(n27845), .A2(N7686), .ZN(N39353));
    NANDX1 U26482 (.A1(n27957), .A2(n15198), .ZN(N39354));
    INVX1 U26483 (.I(n15629), .ZN(n39355));
    NANDX1 U26484 (.A1(n16789), .A2(N8136), .ZN(n39356));
    NANDX1 U26485 (.A1(n13275), .A2(N5225), .ZN(N39357));
    INVX1 U26486 (.I(n28555), .ZN(N39358));
    NOR2X1 U26487 (.A1(n13089), .A2(n20131), .ZN(N39359));
    NANDX1 U26488 (.A1(n23006), .A2(N11956), .ZN(N39360));
    NOR2X1 U26489 (.A1(n13214), .A2(n23625), .ZN(N39361));
    NOR2X1 U26490 (.A1(n26019), .A2(N845), .ZN(n39362));
    NANDX1 U26491 (.A1(n20351), .A2(N7223), .ZN(n39363));
    NANDX1 U26492 (.A1(N6619), .A2(N3469), .ZN(n39364));
    NOR2X1 U26493 (.A1(N4439), .A2(n18667), .ZN(n39365));
    INVX1 U26494 (.I(n20067), .ZN(N39366));
    NOR2X1 U26495 (.A1(N2662), .A2(n16763), .ZN(n39367));
    INVX1 U26496 (.I(N4497), .ZN(N39368));
    INVX1 U26497 (.I(n13237), .ZN(N39369));
    NOR2X1 U26498 (.A1(n13657), .A2(n26325), .ZN(n39370));
    NOR2X1 U26499 (.A1(n25291), .A2(n19193), .ZN(n39371));
    INVX1 U26500 (.I(N5592), .ZN(N39372));
    NOR2X1 U26501 (.A1(n17048), .A2(n29706), .ZN(N39373));
    NANDX1 U26502 (.A1(n17892), .A2(n23037), .ZN(n39374));
    NANDX1 U26503 (.A1(n13676), .A2(n27968), .ZN(N39375));
    NOR2X1 U26504 (.A1(n17144), .A2(n24458), .ZN(N39376));
    INVX1 U26505 (.I(N5673), .ZN(n39377));
    NANDX1 U26506 (.A1(n15306), .A2(n17190), .ZN(N39378));
    NANDX1 U26507 (.A1(n20630), .A2(N8513), .ZN(N39379));
    NANDX1 U26508 (.A1(N12480), .A2(n21749), .ZN(N39380));
    NANDX1 U26509 (.A1(n26136), .A2(N6497), .ZN(n39381));
    INVX1 U26510 (.I(N9851), .ZN(n39382));
    NANDX1 U26511 (.A1(N2551), .A2(N4003), .ZN(N39383));
    INVX1 U26512 (.I(n19598), .ZN(N39384));
    NANDX1 U26513 (.A1(N10489), .A2(n26051), .ZN(n39385));
    NANDX1 U26514 (.A1(n24808), .A2(n28287), .ZN(n39386));
    NOR2X1 U26515 (.A1(N4170), .A2(n15293), .ZN(n39387));
    INVX1 U26516 (.I(n29546), .ZN(N39388));
    INVX1 U26517 (.I(n13469), .ZN(N39389));
    NOR2X1 U26518 (.A1(n26716), .A2(n15020), .ZN(N39390));
    INVX1 U26519 (.I(n23789), .ZN(N39391));
    INVX1 U26520 (.I(N6247), .ZN(n39392));
    NOR2X1 U26521 (.A1(n25850), .A2(n20943), .ZN(N39393));
    INVX1 U26522 (.I(N4840), .ZN(N39394));
    NOR2X1 U26523 (.A1(n24708), .A2(n26089), .ZN(N39395));
    INVX1 U26524 (.I(n29788), .ZN(N39396));
    NOR2X1 U26525 (.A1(N4050), .A2(n28837), .ZN(n39397));
    INVX1 U26526 (.I(N7779), .ZN(N39398));
    INVX1 U26527 (.I(n28309), .ZN(n39399));
    NOR2X1 U26528 (.A1(n16238), .A2(N2026), .ZN(n39400));
    INVX1 U26529 (.I(N4207), .ZN(N39401));
    NOR2X1 U26530 (.A1(n25945), .A2(n26180), .ZN(n39402));
    NOR2X1 U26531 (.A1(n29525), .A2(n19947), .ZN(N39403));
    NANDX1 U26532 (.A1(n27715), .A2(n14754), .ZN(N39404));
    INVX1 U26533 (.I(n23427), .ZN(n39405));
    NOR2X1 U26534 (.A1(N4761), .A2(n16827), .ZN(N39406));
    NOR2X1 U26535 (.A1(n29468), .A2(N12778), .ZN(N39407));
    NOR2X1 U26536 (.A1(n17679), .A2(n16888), .ZN(n39408));
    NOR2X1 U26537 (.A1(n16378), .A2(n16910), .ZN(N39409));
    NOR2X1 U26538 (.A1(n17007), .A2(N3643), .ZN(N39410));
    NOR2X1 U26539 (.A1(N3107), .A2(N5668), .ZN(N39411));
    INVX1 U26540 (.I(n26011), .ZN(n39412));
    INVX1 U26541 (.I(N9083), .ZN(N39413));
    NANDX1 U26542 (.A1(N2470), .A2(n27168), .ZN(N39414));
    NANDX1 U26543 (.A1(N11509), .A2(n24745), .ZN(n39415));
    NANDX1 U26544 (.A1(N5812), .A2(N6595), .ZN(n39416));
    INVX1 U26545 (.I(n29270), .ZN(N39417));
    NANDX1 U26546 (.A1(n30030), .A2(n17161), .ZN(N39418));
    NOR2X1 U26547 (.A1(n13845), .A2(N4703), .ZN(N39419));
    NANDX1 U26548 (.A1(N1708), .A2(N9641), .ZN(N39420));
    NOR2X1 U26549 (.A1(n16048), .A2(n26647), .ZN(N39421));
    NANDX1 U26550 (.A1(N9588), .A2(n18314), .ZN(N39422));
    NOR2X1 U26551 (.A1(N4165), .A2(n14188), .ZN(N39423));
    NOR2X1 U26552 (.A1(n13247), .A2(n24802), .ZN(n39424));
    NOR2X1 U26553 (.A1(n28975), .A2(n25225), .ZN(N39425));
    NANDX1 U26554 (.A1(n23583), .A2(n28963), .ZN(n39426));
    INVX1 U26555 (.I(N40), .ZN(n39427));
    INVX1 U26556 (.I(N5233), .ZN(n39428));
    NANDX1 U26557 (.A1(n15275), .A2(n22394), .ZN(N39429));
    NOR2X1 U26558 (.A1(n17680), .A2(n27096), .ZN(n39430));
    NANDX1 U26559 (.A1(N7948), .A2(n25297), .ZN(N39431));
    NANDX1 U26560 (.A1(n23995), .A2(N10368), .ZN(N39432));
    NOR2X1 U26561 (.A1(n22143), .A2(n28681), .ZN(N39433));
    NOR2X1 U26562 (.A1(n26307), .A2(N1292), .ZN(n39434));
    NOR2X1 U26563 (.A1(n28114), .A2(n26093), .ZN(n39435));
    NANDX1 U26564 (.A1(n26952), .A2(n21181), .ZN(N39436));
    NANDX1 U26565 (.A1(N8958), .A2(N8567), .ZN(N39437));
    NANDX1 U26566 (.A1(n27695), .A2(n23949), .ZN(N39438));
    NANDX1 U26567 (.A1(N9580), .A2(n27784), .ZN(N39439));
    NOR2X1 U26568 (.A1(n27663), .A2(N3887), .ZN(N39440));
    NOR2X1 U26569 (.A1(n15679), .A2(N11834), .ZN(N39441));
    INVX1 U26570 (.I(N1978), .ZN(N39442));
    NANDX1 U26571 (.A1(n26105), .A2(n27596), .ZN(N39443));
    NOR2X1 U26572 (.A1(n13210), .A2(N7791), .ZN(N39444));
    NANDX1 U26573 (.A1(n14501), .A2(n15873), .ZN(N39445));
    INVX1 U26574 (.I(N10457), .ZN(n39446));
    NOR2X1 U26575 (.A1(N3175), .A2(n20198), .ZN(n39447));
    INVX1 U26576 (.I(N12132), .ZN(n39448));
    INVX1 U26577 (.I(n25683), .ZN(n39449));
    INVX1 U26578 (.I(N11136), .ZN(N39450));
    INVX1 U26579 (.I(n19269), .ZN(N39451));
    NOR2X1 U26580 (.A1(n13134), .A2(N5355), .ZN(N39452));
    NOR2X1 U26581 (.A1(N3575), .A2(n21033), .ZN(N39453));
    NOR2X1 U26582 (.A1(n19313), .A2(N11571), .ZN(n39454));
    INVX1 U26583 (.I(N3841), .ZN(n39455));
    NANDX1 U26584 (.A1(N12270), .A2(n17050), .ZN(N39456));
    NANDX1 U26585 (.A1(n13395), .A2(N1414), .ZN(n39457));
    INVX1 U26586 (.I(n19756), .ZN(n39458));
    NANDX1 U26587 (.A1(n26730), .A2(n22930), .ZN(N39459));
    NOR2X1 U26588 (.A1(N3403), .A2(N4925), .ZN(n39460));
    NOR2X1 U26589 (.A1(n17647), .A2(N3175), .ZN(N39461));
    INVX1 U26590 (.I(n14419), .ZN(n39462));
    NOR2X1 U26591 (.A1(N4854), .A2(n27553), .ZN(N39463));
    NANDX1 U26592 (.A1(n24781), .A2(n19688), .ZN(n39464));
    NOR2X1 U26593 (.A1(n26404), .A2(n27561), .ZN(N39465));
    NOR2X1 U26594 (.A1(n22279), .A2(N1265), .ZN(n39466));
    INVX1 U26595 (.I(n23109), .ZN(N39467));
    INVX1 U26596 (.I(N10355), .ZN(N39468));
    NANDX1 U26597 (.A1(N8288), .A2(n20168), .ZN(n39469));
    INVX1 U26598 (.I(n27416), .ZN(n39470));
    NANDX1 U26599 (.A1(N7475), .A2(N6467), .ZN(n39471));
    NANDX1 U26600 (.A1(N960), .A2(N2843), .ZN(N39472));
    NANDX1 U26601 (.A1(N4134), .A2(n29052), .ZN(N39473));
    NOR2X1 U26602 (.A1(n15137), .A2(n22466), .ZN(n39474));
    NANDX1 U26603 (.A1(N1357), .A2(n17109), .ZN(N39475));
    INVX1 U26604 (.I(n27308), .ZN(n39476));
    INVX1 U26605 (.I(n20998), .ZN(N39477));
    NOR2X1 U26606 (.A1(N12775), .A2(N10823), .ZN(n39478));
    INVX1 U26607 (.I(N5747), .ZN(n39479));
    NANDX1 U26608 (.A1(N8444), .A2(n19372), .ZN(N39480));
    INVX1 U26609 (.I(n28611), .ZN(n39481));
    NOR2X1 U26610 (.A1(N11824), .A2(n22493), .ZN(N39482));
    NANDX1 U26611 (.A1(n18291), .A2(n19778), .ZN(n39483));
    INVX1 U26612 (.I(n21133), .ZN(N39484));
    NOR2X1 U26613 (.A1(n23743), .A2(N8608), .ZN(N39485));
    NOR2X1 U26614 (.A1(N8743), .A2(N936), .ZN(N39486));
    INVX1 U26615 (.I(n28797), .ZN(N39487));
    INVX1 U26616 (.I(n15624), .ZN(N39488));
    NANDX1 U26617 (.A1(N8541), .A2(n25182), .ZN(N39489));
    NANDX1 U26618 (.A1(N9877), .A2(N5867), .ZN(N39490));
    NANDX1 U26619 (.A1(N4184), .A2(N12124), .ZN(N39491));
    NANDX1 U26620 (.A1(n23555), .A2(n26669), .ZN(n39492));
    INVX1 U26621 (.I(n16032), .ZN(n39493));
    NANDX1 U26622 (.A1(n16443), .A2(n15983), .ZN(N39494));
    NOR2X1 U26623 (.A1(N6083), .A2(N5455), .ZN(n39495));
    INVX1 U26624 (.I(n17913), .ZN(N39496));
    NANDX1 U26625 (.A1(n14809), .A2(n17515), .ZN(N39497));
    INVX1 U26626 (.I(N4305), .ZN(n39498));
    NOR2X1 U26627 (.A1(n25160), .A2(n29608), .ZN(N39499));
    NANDX1 U26628 (.A1(n20990), .A2(N8012), .ZN(N39500));
    INVX1 U26629 (.I(N9934), .ZN(N39501));
    NOR2X1 U26630 (.A1(n14659), .A2(n27105), .ZN(N39502));
    NOR2X1 U26631 (.A1(n26782), .A2(n22581), .ZN(N39503));
    NANDX1 U26632 (.A1(n23314), .A2(n16531), .ZN(n39504));
    INVX1 U26633 (.I(n20230), .ZN(n39505));
    INVX1 U26634 (.I(n24623), .ZN(N39506));
    NOR2X1 U26635 (.A1(n27617), .A2(n18639), .ZN(N39507));
    INVX1 U26636 (.I(n15392), .ZN(N39508));
    INVX1 U26637 (.I(n14869), .ZN(N39509));
    NANDX1 U26638 (.A1(N2623), .A2(n19173), .ZN(n39510));
    NANDX1 U26639 (.A1(n27782), .A2(N7205), .ZN(N39511));
    NOR2X1 U26640 (.A1(N7195), .A2(n15216), .ZN(N39512));
    INVX1 U26641 (.I(N5690), .ZN(n39513));
    NANDX1 U26642 (.A1(n26654), .A2(n21355), .ZN(n39514));
    INVX1 U26643 (.I(N11859), .ZN(n39515));
    NANDX1 U26644 (.A1(n24904), .A2(N5035), .ZN(N39516));
    NOR2X1 U26645 (.A1(N3407), .A2(n25264), .ZN(N39517));
    INVX1 U26646 (.I(n16590), .ZN(n39518));
    NANDX1 U26647 (.A1(n19205), .A2(N5091), .ZN(N39519));
    NANDX1 U26648 (.A1(n23158), .A2(n30048), .ZN(n39520));
    NANDX1 U26649 (.A1(N3049), .A2(N2533), .ZN(N39521));
    NOR2X1 U26650 (.A1(n22641), .A2(n18876), .ZN(N39522));
    NANDX1 U26651 (.A1(N7146), .A2(n14631), .ZN(n39523));
    INVX1 U26652 (.I(n19141), .ZN(N39524));
    INVX1 U26653 (.I(n14154), .ZN(n39525));
    INVX1 U26654 (.I(N98), .ZN(N39526));
    NANDX1 U26655 (.A1(n27515), .A2(N2457), .ZN(N39527));
    NOR2X1 U26656 (.A1(n21111), .A2(N2648), .ZN(N39528));
    NOR2X1 U26657 (.A1(N4798), .A2(n24373), .ZN(n39529));
    INVX1 U26658 (.I(n23921), .ZN(N39530));
    NOR2X1 U26659 (.A1(N1846), .A2(n24405), .ZN(N39531));
    NOR2X1 U26660 (.A1(n20454), .A2(N9621), .ZN(n39532));
    INVX1 U26661 (.I(n22987), .ZN(N39533));
    NOR2X1 U26662 (.A1(N9270), .A2(N286), .ZN(N39534));
    INVX1 U26663 (.I(N4976), .ZN(N39535));
    NOR2X1 U26664 (.A1(N6652), .A2(N12677), .ZN(N39536));
    INVX1 U26665 (.I(N9366), .ZN(N39537));
    NOR2X1 U26666 (.A1(N1016), .A2(n14237), .ZN(n39538));
    NANDX1 U26667 (.A1(N3472), .A2(N2435), .ZN(N39539));
    NANDX1 U26668 (.A1(N6119), .A2(N12737), .ZN(N39540));
    NANDX1 U26669 (.A1(n19052), .A2(N9491), .ZN(n39541));
    INVX1 U26670 (.I(N9614), .ZN(n39542));
    NOR2X1 U26671 (.A1(N5352), .A2(n23332), .ZN(N39543));
    NOR2X1 U26672 (.A1(N3533), .A2(N9962), .ZN(N39544));
    INVX1 U26673 (.I(N6102), .ZN(N39545));
    NOR2X1 U26674 (.A1(N2046), .A2(n27522), .ZN(n39546));
    NOR2X1 U26675 (.A1(N5522), .A2(n22734), .ZN(N39547));
    INVX1 U26676 (.I(n17879), .ZN(N39548));
    INVX1 U26677 (.I(n19460), .ZN(n39549));
    NANDX1 U26678 (.A1(N4759), .A2(n22292), .ZN(n39550));
    NOR2X1 U26679 (.A1(N7193), .A2(N4658), .ZN(N39551));
    INVX1 U26680 (.I(n19929), .ZN(N39552));
    NOR2X1 U26681 (.A1(n24658), .A2(n29419), .ZN(N39553));
    NANDX1 U26682 (.A1(N4134), .A2(n29316), .ZN(N39554));
    INVX1 U26683 (.I(n16027), .ZN(N39555));
    INVX1 U26684 (.I(n19047), .ZN(N39556));
    NANDX1 U26685 (.A1(n21289), .A2(n25148), .ZN(N39557));
    NANDX1 U26686 (.A1(n23334), .A2(N11093), .ZN(N39558));
    INVX1 U26687 (.I(n17416), .ZN(n39559));
    NOR2X1 U26688 (.A1(n14795), .A2(N5158), .ZN(N39560));
    INVX1 U26689 (.I(N4117), .ZN(N39561));
    INVX1 U26690 (.I(n29106), .ZN(n39562));
    INVX1 U26691 (.I(n23539), .ZN(N39563));
    INVX1 U26692 (.I(n19626), .ZN(N39564));
    INVX1 U26693 (.I(N3211), .ZN(N39565));
    INVX1 U26694 (.I(N12227), .ZN(N39566));
    NANDX1 U26695 (.A1(N2911), .A2(N4921), .ZN(N39567));
    NOR2X1 U26696 (.A1(n18425), .A2(n20947), .ZN(N39568));
    INVX1 U26697 (.I(N7334), .ZN(N39569));
    NOR2X1 U26698 (.A1(N8169), .A2(n21042), .ZN(N39570));
    NANDX1 U26699 (.A1(N1365), .A2(N1997), .ZN(N39571));
    NOR2X1 U26700 (.A1(N7342), .A2(n24383), .ZN(N39572));
    NANDX1 U26701 (.A1(N1060), .A2(n18593), .ZN(N39573));
    NOR2X1 U26702 (.A1(n13672), .A2(N6122), .ZN(N39574));
    NOR2X1 U26703 (.A1(n25771), .A2(N843), .ZN(N39575));
    INVX1 U26704 (.I(n13340), .ZN(N39576));
    INVX1 U26705 (.I(n28982), .ZN(n39577));
    NOR2X1 U26706 (.A1(n25243), .A2(N1755), .ZN(N39578));
    NOR2X1 U26707 (.A1(N4034), .A2(N8741), .ZN(N39579));
    NOR2X1 U26708 (.A1(N2354), .A2(N4635), .ZN(n39580));
    NANDX1 U26709 (.A1(N10522), .A2(n25677), .ZN(N39581));
    INVX1 U26710 (.I(N448), .ZN(N39582));
    NANDX1 U26711 (.A1(N6944), .A2(n26487), .ZN(n39583));
    NANDX1 U26712 (.A1(n27346), .A2(n27546), .ZN(N39584));
    NANDX1 U26713 (.A1(N10289), .A2(N11080), .ZN(n39585));
    INVX1 U26714 (.I(N8199), .ZN(N39586));
    INVX1 U26715 (.I(n13158), .ZN(N39587));
    NANDX1 U26716 (.A1(N8613), .A2(N5772), .ZN(N39588));
    NANDX1 U26717 (.A1(n22739), .A2(N877), .ZN(N39589));
    NOR2X1 U26718 (.A1(N11649), .A2(n23608), .ZN(n39590));
    INVX1 U26719 (.I(n21505), .ZN(N39591));
    NANDX1 U26720 (.A1(n28269), .A2(N6581), .ZN(N39592));
    NOR2X1 U26721 (.A1(N12369), .A2(n15175), .ZN(N39593));
    NANDX1 U26722 (.A1(n28602), .A2(N10679), .ZN(n39594));
    INVX1 U26723 (.I(n27642), .ZN(N39595));
    NANDX1 U26724 (.A1(N7809), .A2(n15138), .ZN(N39596));
    NOR2X1 U26725 (.A1(N7449), .A2(n27453), .ZN(n39597));
    INVX1 U26726 (.I(n21420), .ZN(N39598));
    NOR2X1 U26727 (.A1(N10532), .A2(n18594), .ZN(n39599));
    INVX1 U26728 (.I(N4973), .ZN(n39600));
    NANDX1 U26729 (.A1(n24379), .A2(n19866), .ZN(n39601));
    INVX1 U26730 (.I(n17850), .ZN(N39602));
    INVX1 U26731 (.I(n14210), .ZN(N39603));
    INVX1 U26732 (.I(N55), .ZN(n39604));
    NOR2X1 U26733 (.A1(n15838), .A2(N12423), .ZN(n39605));
    NANDX1 U26734 (.A1(n18450), .A2(N10887), .ZN(N39606));
    INVX1 U26735 (.I(n17411), .ZN(n39607));
    NANDX1 U26736 (.A1(n20212), .A2(n13780), .ZN(N39608));
    NOR2X1 U26737 (.A1(n26948), .A2(N9789), .ZN(N39609));
    NOR2X1 U26738 (.A1(N11745), .A2(N1072), .ZN(N39610));
    NANDX1 U26739 (.A1(n22276), .A2(n19665), .ZN(N39611));
    INVX1 U26740 (.I(n15809), .ZN(n39612));
    NOR2X1 U26741 (.A1(n14743), .A2(N5537), .ZN(N39613));
    INVX1 U26742 (.I(n21153), .ZN(n39614));
    NOR2X1 U26743 (.A1(n14896), .A2(N11948), .ZN(N39615));
    INVX1 U26744 (.I(N12808), .ZN(N39616));
    NANDX1 U26745 (.A1(n19936), .A2(n25894), .ZN(N39617));
    NOR2X1 U26746 (.A1(n19384), .A2(n19521), .ZN(N39618));
    NOR2X1 U26747 (.A1(N4897), .A2(n28294), .ZN(n39619));
    NOR2X1 U26748 (.A1(n16986), .A2(n25104), .ZN(n39620));
    NANDX1 U26749 (.A1(N3512), .A2(n25409), .ZN(N39621));
    NOR2X1 U26750 (.A1(n19208), .A2(N6108), .ZN(N39622));
    INVX1 U26751 (.I(n28270), .ZN(N39623));
    NANDX1 U26752 (.A1(N2640), .A2(N1437), .ZN(N39624));
    INVX1 U26753 (.I(N3326), .ZN(N39625));
    INVX1 U26754 (.I(n23473), .ZN(N39626));
    NANDX1 U26755 (.A1(N4399), .A2(N849), .ZN(N39627));
    NANDX1 U26756 (.A1(n20745), .A2(N9346), .ZN(N39628));
    NANDX1 U26757 (.A1(n25403), .A2(n17290), .ZN(N39629));
    INVX1 U26758 (.I(N5895), .ZN(n39630));
    INVX1 U26759 (.I(N10145), .ZN(N39631));
    INVX1 U26760 (.I(n27732), .ZN(n39632));
    NOR2X1 U26761 (.A1(n15667), .A2(n19804), .ZN(N39633));
    INVX1 U26762 (.I(N9359), .ZN(N39634));
    NOR2X1 U26763 (.A1(n13748), .A2(n22716), .ZN(N39635));
    INVX1 U26764 (.I(n24224), .ZN(N39636));
    INVX1 U26765 (.I(n27141), .ZN(N39637));
    NOR2X1 U26766 (.A1(n17241), .A2(n19592), .ZN(N39638));
    INVX1 U26767 (.I(n24022), .ZN(n39639));
    NANDX1 U26768 (.A1(n22981), .A2(n13474), .ZN(n39640));
    INVX1 U26769 (.I(n20887), .ZN(n39641));
    NANDX1 U26770 (.A1(N5683), .A2(n26737), .ZN(N39642));
    NOR2X1 U26771 (.A1(N11577), .A2(N7346), .ZN(N39643));
    NANDX1 U26772 (.A1(N11744), .A2(n23638), .ZN(n39644));
    NANDX1 U26773 (.A1(n15971), .A2(n13304), .ZN(N39645));
    NOR2X1 U26774 (.A1(n25329), .A2(N10738), .ZN(N39646));
    NOR2X1 U26775 (.A1(N6468), .A2(N6305), .ZN(N39647));
    NOR2X1 U26776 (.A1(n20383), .A2(N3308), .ZN(n39648));
    NANDX1 U26777 (.A1(N7486), .A2(N11461), .ZN(N39649));
    NOR2X1 U26778 (.A1(N1371), .A2(N12573), .ZN(n39650));
    NANDX1 U26779 (.A1(N3405), .A2(N4292), .ZN(n39651));
    INVX1 U26780 (.I(N9346), .ZN(n39652));
    INVX1 U26781 (.I(n26761), .ZN(N39653));
    INVX1 U26782 (.I(n21550), .ZN(N39654));
    NANDX1 U26783 (.A1(N6513), .A2(n21854), .ZN(n39655));
    NOR2X1 U26784 (.A1(n28257), .A2(N7687), .ZN(N39656));
    INVX1 U26785 (.I(N8806), .ZN(n39657));
    INVX1 U26786 (.I(n28768), .ZN(N39658));
    INVX1 U26787 (.I(n16605), .ZN(n39659));
    INVX1 U26788 (.I(n28880), .ZN(n39660));
    NANDX1 U26789 (.A1(n15502), .A2(n15922), .ZN(N39661));
    INVX1 U26790 (.I(n26962), .ZN(N39662));
    NANDX1 U26791 (.A1(N4267), .A2(n28095), .ZN(N39663));
    NOR2X1 U26792 (.A1(n26370), .A2(N2249), .ZN(N39664));
    INVX1 U26793 (.I(N5578), .ZN(n39665));
    INVX1 U26794 (.I(N8139), .ZN(N39666));
    NOR2X1 U26795 (.A1(n22333), .A2(N668), .ZN(n39667));
    NOR2X1 U26796 (.A1(n14049), .A2(N5395), .ZN(n39668));
    NANDX1 U26797 (.A1(N10297), .A2(n23425), .ZN(N39669));
    NOR2X1 U26798 (.A1(N1736), .A2(n22055), .ZN(n39670));
    INVX1 U26799 (.I(n18340), .ZN(n39671));
    INVX1 U26800 (.I(n13817), .ZN(N39672));
    NOR2X1 U26801 (.A1(n19614), .A2(n18299), .ZN(n39673));
    INVX1 U26802 (.I(N4999), .ZN(N39674));
    NOR2X1 U26803 (.A1(n20914), .A2(N2957), .ZN(n39675));
    NOR2X1 U26804 (.A1(N5707), .A2(n23903), .ZN(n39676));
    INVX1 U26805 (.I(n29983), .ZN(n39677));
    NOR2X1 U26806 (.A1(n14263), .A2(n21259), .ZN(n39678));
    NOR2X1 U26807 (.A1(n14930), .A2(n19047), .ZN(N39679));
    NANDX1 U26808 (.A1(n20324), .A2(N3516), .ZN(N39680));
    NANDX1 U26809 (.A1(N2172), .A2(n26928), .ZN(N39681));
    NOR2X1 U26810 (.A1(N12788), .A2(N11865), .ZN(N39682));
    INVX1 U26811 (.I(n16899), .ZN(n39683));
    NOR2X1 U26812 (.A1(N3337), .A2(n25073), .ZN(n39684));
    NANDX1 U26813 (.A1(n19984), .A2(n18633), .ZN(N39685));
    NANDX1 U26814 (.A1(n29459), .A2(N10150), .ZN(N39686));
    NOR2X1 U26815 (.A1(N5028), .A2(N3915), .ZN(N39687));
    NOR2X1 U26816 (.A1(N4873), .A2(N9902), .ZN(n39688));
    INVX1 U26817 (.I(n14692), .ZN(n39689));
    NOR2X1 U26818 (.A1(n18527), .A2(N3602), .ZN(n39690));
    NANDX1 U26819 (.A1(N8714), .A2(N7117), .ZN(n39691));
    INVX1 U26820 (.I(n29583), .ZN(N39692));
    NOR2X1 U26821 (.A1(n28606), .A2(N12233), .ZN(n39693));
    NOR2X1 U26822 (.A1(n18192), .A2(n29132), .ZN(n39694));
    NOR2X1 U26823 (.A1(N10089), .A2(N12628), .ZN(N39695));
    NANDX1 U26824 (.A1(n18634), .A2(N1123), .ZN(n39696));
    INVX1 U26825 (.I(N6516), .ZN(N39697));
    INVX1 U26826 (.I(n27104), .ZN(N39698));
    NANDX1 U26827 (.A1(n15187), .A2(n27878), .ZN(N39699));
    NANDX1 U26828 (.A1(n13649), .A2(N12777), .ZN(N39700));
    NOR2X1 U26829 (.A1(N10294), .A2(N1166), .ZN(N39701));
    INVX1 U26830 (.I(n26428), .ZN(N39702));
    NANDX1 U26831 (.A1(N7508), .A2(n23512), .ZN(N39703));
    INVX1 U26832 (.I(n30112), .ZN(N39704));
    INVX1 U26833 (.I(N10118), .ZN(n39705));
    NOR2X1 U26834 (.A1(n28732), .A2(n27810), .ZN(N39706));
    NOR2X1 U26835 (.A1(n27382), .A2(n28999), .ZN(N39707));
    INVX1 U26836 (.I(N4439), .ZN(N39708));
    NANDX1 U26837 (.A1(N11856), .A2(N10954), .ZN(N39709));
    INVX1 U26838 (.I(n27521), .ZN(n39710));
    INVX1 U26839 (.I(n15003), .ZN(N39711));
    NANDX1 U26840 (.A1(N4594), .A2(n17212), .ZN(n39712));
    NOR2X1 U26841 (.A1(N12823), .A2(n16066), .ZN(N39713));
    NOR2X1 U26842 (.A1(n13213), .A2(N12356), .ZN(N39714));
    NOR2X1 U26843 (.A1(n20720), .A2(n24429), .ZN(N39715));
    INVX1 U26844 (.I(n20695), .ZN(n39716));
    NOR2X1 U26845 (.A1(N11327), .A2(n25001), .ZN(N39717));
    NOR2X1 U26846 (.A1(n27698), .A2(n25002), .ZN(N39718));
    NOR2X1 U26847 (.A1(n26559), .A2(N4403), .ZN(n39719));
    INVX1 U26848 (.I(n15103), .ZN(N39720));
    NOR2X1 U26849 (.A1(n23321), .A2(n14919), .ZN(N39721));
    NANDX1 U26850 (.A1(n22938), .A2(n18482), .ZN(N39722));
    INVX1 U26851 (.I(n27532), .ZN(n39723));
    NANDX1 U26852 (.A1(N12483), .A2(N10217), .ZN(N39724));
    INVX1 U26853 (.I(n28807), .ZN(N39725));
    NOR2X1 U26854 (.A1(n22539), .A2(N1994), .ZN(N39726));
    NOR2X1 U26855 (.A1(N5391), .A2(N3203), .ZN(N39727));
    NANDX1 U26856 (.A1(N10222), .A2(n14529), .ZN(n39728));
    INVX1 U26857 (.I(N2209), .ZN(N39729));
    NOR2X1 U26858 (.A1(N1555), .A2(N10138), .ZN(N39730));
    NOR2X1 U26859 (.A1(N5957), .A2(n22505), .ZN(N39731));
    NANDX1 U26860 (.A1(N10775), .A2(N4249), .ZN(n39732));
    INVX1 U26861 (.I(n12977), .ZN(N39733));
    INVX1 U26862 (.I(N11257), .ZN(N39734));
    INVX1 U26863 (.I(n24581), .ZN(n39735));
    INVX1 U26864 (.I(n18604), .ZN(N39736));
    NANDX1 U26865 (.A1(n26995), .A2(n17273), .ZN(N39737));
    INVX1 U26866 (.I(n19396), .ZN(n39738));
    NANDX1 U26867 (.A1(N7782), .A2(n13347), .ZN(n39739));
    NANDX1 U26868 (.A1(n19609), .A2(n23569), .ZN(N39740));
    NANDX1 U26869 (.A1(n26299), .A2(n25777), .ZN(N39741));
    NOR2X1 U26870 (.A1(n16414), .A2(n24476), .ZN(n39742));
    NANDX1 U26871 (.A1(n22370), .A2(n16843), .ZN(N39743));
    INVX1 U26872 (.I(n21706), .ZN(n39744));
    INVX1 U26873 (.I(N12606), .ZN(N39745));
    NOR2X1 U26874 (.A1(n18141), .A2(n23862), .ZN(n39746));
    NOR2X1 U26875 (.A1(N1145), .A2(n29235), .ZN(n39747));
    INVX1 U26876 (.I(n24502), .ZN(N39748));
    INVX1 U26877 (.I(N4964), .ZN(n39749));
    NOR2X1 U26878 (.A1(N3912), .A2(N12790), .ZN(n39750));
    INVX1 U26879 (.I(n17258), .ZN(N39751));
    INVX1 U26880 (.I(N4086), .ZN(n39752));
    NOR2X1 U26881 (.A1(n19238), .A2(n18946), .ZN(n39753));
    NOR2X1 U26882 (.A1(n22566), .A2(N5222), .ZN(N39754));
    INVX1 U26883 (.I(N11525), .ZN(N39755));
    INVX1 U26884 (.I(n13329), .ZN(N39756));
    INVX1 U26885 (.I(N7721), .ZN(N39757));
    INVX1 U26886 (.I(N2385), .ZN(N39758));
    NANDX1 U26887 (.A1(N10984), .A2(n14807), .ZN(N39759));
    NANDX1 U26888 (.A1(N689), .A2(n13904), .ZN(N39760));
    INVX1 U26889 (.I(n13751), .ZN(N39761));
    NANDX1 U26890 (.A1(n22843), .A2(N1886), .ZN(n39762));
    NOR2X1 U26891 (.A1(n24194), .A2(N5061), .ZN(N39763));
    NOR2X1 U26892 (.A1(n17874), .A2(N9146), .ZN(n39764));
    NANDX1 U26893 (.A1(n25672), .A2(n28091), .ZN(N39765));
    INVX1 U26894 (.I(n18100), .ZN(N39766));
    NANDX1 U26895 (.A1(n17471), .A2(n29625), .ZN(n39767));
    NANDX1 U26896 (.A1(N663), .A2(n19404), .ZN(N39768));
    NANDX1 U26897 (.A1(n23643), .A2(N10349), .ZN(n39769));
    NOR2X1 U26898 (.A1(N4490), .A2(n25155), .ZN(N39770));
    NANDX1 U26899 (.A1(n23876), .A2(n27619), .ZN(N39771));
    NANDX1 U26900 (.A1(N7490), .A2(n26037), .ZN(n39772));
    NOR2X1 U26901 (.A1(N9375), .A2(n16928), .ZN(N39773));
    NANDX1 U26902 (.A1(n14435), .A2(n13637), .ZN(n39774));
    INVX1 U26903 (.I(N12141), .ZN(n39775));
    NOR2X1 U26904 (.A1(n18914), .A2(n28793), .ZN(N39776));
    NANDX1 U26905 (.A1(N6876), .A2(n20529), .ZN(n39777));
    INVX1 U26906 (.I(n25061), .ZN(N39778));
    NOR2X1 U26907 (.A1(N7136), .A2(N2888), .ZN(N39779));
    INVX1 U26908 (.I(N642), .ZN(n39780));
    NANDX1 U26909 (.A1(n14702), .A2(n23829), .ZN(N39781));
    NOR2X1 U26910 (.A1(n27005), .A2(n17567), .ZN(N39782));
    NOR2X1 U26911 (.A1(N8353), .A2(n25056), .ZN(N39783));
    INVX1 U26912 (.I(n19802), .ZN(n39784));
    INVX1 U26913 (.I(N7122), .ZN(n39785));
    NOR2X1 U26914 (.A1(n25986), .A2(n20758), .ZN(N39786));
    INVX1 U26915 (.I(n26688), .ZN(N39787));
    NOR2X1 U26916 (.A1(N7324), .A2(n13904), .ZN(N39788));
    NANDX1 U26917 (.A1(n14200), .A2(n22993), .ZN(N39789));
    NOR2X1 U26918 (.A1(n27821), .A2(N9833), .ZN(N39790));
    NANDX1 U26919 (.A1(N572), .A2(n19540), .ZN(N39791));
    NOR2X1 U26920 (.A1(n13807), .A2(N4104), .ZN(N39792));
    NOR2X1 U26921 (.A1(N10621), .A2(N971), .ZN(N39793));
    INVX1 U26922 (.I(N4915), .ZN(N39794));
    NOR2X1 U26923 (.A1(N5464), .A2(n13807), .ZN(N39795));
    INVX1 U26924 (.I(n17016), .ZN(n39796));
    NOR2X1 U26925 (.A1(N12854), .A2(N1425), .ZN(N39797));
    NOR2X1 U26926 (.A1(N1265), .A2(n28112), .ZN(N39798));
    INVX1 U26927 (.I(N8588), .ZN(n39799));
    INVX1 U26928 (.I(N8239), .ZN(N39800));
    NANDX1 U26929 (.A1(N4733), .A2(N3930), .ZN(N39801));
    NOR2X1 U26930 (.A1(N3126), .A2(n25455), .ZN(n39802));
    NANDX1 U26931 (.A1(n22665), .A2(n17483), .ZN(N39803));
    NOR2X1 U26932 (.A1(n15329), .A2(n21901), .ZN(N39804));
    INVX1 U26933 (.I(N4861), .ZN(N39805));
    NANDX1 U26934 (.A1(n16066), .A2(n21442), .ZN(N39806));
    NOR2X1 U26935 (.A1(n29872), .A2(n27688), .ZN(n39807));
    INVX1 U26936 (.I(N9224), .ZN(N39808));
    NANDX1 U26937 (.A1(n14773), .A2(N9332), .ZN(N39809));
    INVX1 U26938 (.I(N1308), .ZN(N39810));
    NANDX1 U26939 (.A1(n27515), .A2(n13186), .ZN(N39811));
    INVX1 U26940 (.I(n27423), .ZN(n39812));
    NOR2X1 U26941 (.A1(n17643), .A2(n25015), .ZN(N39813));
    INVX1 U26942 (.I(n12960), .ZN(N39814));
    NANDX1 U26943 (.A1(n20830), .A2(n19004), .ZN(N39815));
    NANDX1 U26944 (.A1(n24720), .A2(n29465), .ZN(N39816));
    NOR2X1 U26945 (.A1(n29580), .A2(N1636), .ZN(N39817));
    NOR2X1 U26946 (.A1(N9445), .A2(n28105), .ZN(N39818));
    NANDX1 U26947 (.A1(N6995), .A2(N11316), .ZN(n39819));
    NOR2X1 U26948 (.A1(N5960), .A2(n14649), .ZN(N39820));
    INVX1 U26949 (.I(n24886), .ZN(N39821));
    INVX1 U26950 (.I(N2975), .ZN(N39822));
    NOR2X1 U26951 (.A1(n17702), .A2(n16688), .ZN(N39823));
    NOR2X1 U26952 (.A1(N12742), .A2(N4193), .ZN(n39824));
    NOR2X1 U26953 (.A1(N10907), .A2(N5714), .ZN(N39825));
    NANDX1 U26954 (.A1(n20297), .A2(n13278), .ZN(n39826));
    INVX1 U26955 (.I(n14879), .ZN(N39827));
    NANDX1 U26956 (.A1(n13018), .A2(N2882), .ZN(N39828));
    INVX1 U26957 (.I(N3668), .ZN(n39829));
    INVX1 U26958 (.I(n19466), .ZN(N39830));
    NANDX1 U26959 (.A1(n19321), .A2(n19342), .ZN(N39831));
    NANDX1 U26960 (.A1(n13841), .A2(N3853), .ZN(n39832));
    NANDX1 U26961 (.A1(N8590), .A2(N8370), .ZN(N39833));
    NANDX1 U26962 (.A1(n19413), .A2(n26071), .ZN(N39834));
    NANDX1 U26963 (.A1(n16083), .A2(N8675), .ZN(n39835));
    INVX1 U26964 (.I(N7631), .ZN(n39836));
    NOR2X1 U26965 (.A1(N12365), .A2(n22356), .ZN(N39837));
    INVX1 U26966 (.I(n25642), .ZN(N39838));
    NOR2X1 U26967 (.A1(N1741), .A2(n26807), .ZN(N39839));
    NOR2X1 U26968 (.A1(N4623), .A2(n29607), .ZN(n39840));
    INVX1 U26969 (.I(N5510), .ZN(N39841));
    NOR2X1 U26970 (.A1(N7070), .A2(n13391), .ZN(N39842));
    NOR2X1 U26971 (.A1(n26685), .A2(n27232), .ZN(N39843));
    INVX1 U26972 (.I(n20922), .ZN(n39844));
    INVX1 U26973 (.I(n27620), .ZN(n39845));
    INVX1 U26974 (.I(n13657), .ZN(N39846));
    NANDX1 U26975 (.A1(N1893), .A2(n29740), .ZN(N39847));
    NANDX1 U26976 (.A1(N8544), .A2(n25931), .ZN(N39848));
    NANDX1 U26977 (.A1(n20908), .A2(N6710), .ZN(N39849));
    NANDX1 U26978 (.A1(n16412), .A2(n25922), .ZN(N39850));
    NANDX1 U26979 (.A1(N1642), .A2(n28014), .ZN(N39851));
    NOR2X1 U26980 (.A1(n19809), .A2(N10896), .ZN(N39852));
    NOR2X1 U26981 (.A1(n27304), .A2(n17965), .ZN(N39853));
    NOR2X1 U26982 (.A1(n24004), .A2(N3074), .ZN(N39854));
    NANDX1 U26983 (.A1(N1679), .A2(n23995), .ZN(N39855));
    NANDX1 U26984 (.A1(n29298), .A2(N11989), .ZN(N39856));
    NOR2X1 U26985 (.A1(n29973), .A2(N2442), .ZN(n39857));
    NANDX1 U26986 (.A1(N9186), .A2(N10985), .ZN(n39858));
    INVX1 U26987 (.I(n26677), .ZN(n39859));
    NOR2X1 U26988 (.A1(N9656), .A2(N893), .ZN(N39860));
    NOR2X1 U26989 (.A1(N5440), .A2(N6986), .ZN(n39861));
    NANDX1 U26990 (.A1(n22015), .A2(N6263), .ZN(N39862));
    INVX1 U26991 (.I(N2773), .ZN(N39863));
    INVX1 U26992 (.I(n13904), .ZN(N39864));
    INVX1 U26993 (.I(N6346), .ZN(N39865));
    INVX1 U26994 (.I(N932), .ZN(N39866));
    NANDX1 U26995 (.A1(n28146), .A2(n24926), .ZN(N39867));
    NOR2X1 U26996 (.A1(n15868), .A2(n25476), .ZN(N39868));
    NOR2X1 U26997 (.A1(n15703), .A2(n16478), .ZN(n39869));
    INVX1 U26998 (.I(n24888), .ZN(N39870));
    NANDX1 U26999 (.A1(N3026), .A2(N9988), .ZN(N39871));
    INVX1 U27000 (.I(N12681), .ZN(N39872));
    NANDX1 U27001 (.A1(n13066), .A2(N6682), .ZN(n39873));
    NOR2X1 U27002 (.A1(n28692), .A2(n17257), .ZN(n39874));
    INVX1 U27003 (.I(n15292), .ZN(N39875));
    NANDX1 U27004 (.A1(n23736), .A2(n17756), .ZN(N39876));
    NOR2X1 U27005 (.A1(n30082), .A2(n14086), .ZN(N39877));
    NANDX1 U27006 (.A1(n17380), .A2(N656), .ZN(n39878));
    NOR2X1 U27007 (.A1(N2754), .A2(N5084), .ZN(N39879));
    INVX1 U27008 (.I(n25816), .ZN(N39880));
    INVX1 U27009 (.I(n21243), .ZN(n39881));
    NOR2X1 U27010 (.A1(N4098), .A2(n18568), .ZN(N39882));
    NANDX1 U27011 (.A1(n14085), .A2(n24906), .ZN(N39883));
    INVX1 U27012 (.I(n24965), .ZN(N39884));
    INVX1 U27013 (.I(N6705), .ZN(N39885));
    NANDX1 U27014 (.A1(n13648), .A2(N12522), .ZN(N39886));
    NOR2X1 U27015 (.A1(n28939), .A2(n21111), .ZN(n39887));
    NANDX1 U27016 (.A1(n16557), .A2(n27558), .ZN(n39888));
    INVX1 U27017 (.I(n19203), .ZN(N39889));
    NOR2X1 U27018 (.A1(n13425), .A2(N8419), .ZN(N39890));
    NOR2X1 U27019 (.A1(N4739), .A2(n13502), .ZN(n39891));
    INVX1 U27020 (.I(N417), .ZN(N39892));
    NANDX1 U27021 (.A1(n21535), .A2(n14871), .ZN(n39893));
    NOR2X1 U27022 (.A1(n28663), .A2(n13653), .ZN(N39894));
    NANDX1 U27023 (.A1(N11993), .A2(n13676), .ZN(N39895));
    INVX1 U27024 (.I(n27085), .ZN(N39896));
    NOR2X1 U27025 (.A1(N2793), .A2(N10595), .ZN(N39897));
    NANDX1 U27026 (.A1(n16734), .A2(n28094), .ZN(n39898));
    INVX1 U27027 (.I(N12835), .ZN(N39899));
    INVX1 U27028 (.I(n17114), .ZN(n39900));
    NANDX1 U27029 (.A1(n22277), .A2(N10475), .ZN(N39901));
    NANDX1 U27030 (.A1(N558), .A2(n24701), .ZN(N39902));
    NOR2X1 U27031 (.A1(N2621), .A2(n13554), .ZN(n39903));
    NOR2X1 U27032 (.A1(n25469), .A2(n23650), .ZN(N39904));
    NOR2X1 U27033 (.A1(N10838), .A2(n22175), .ZN(N39905));
    NANDX1 U27034 (.A1(n28989), .A2(n22728), .ZN(N39906));
    INVX1 U27035 (.I(N392), .ZN(N39907));
    INVX1 U27036 (.I(N9961), .ZN(n39908));
    NOR2X1 U27037 (.A1(N7392), .A2(n19983), .ZN(n39909));
    NOR2X1 U27038 (.A1(N5349), .A2(n20978), .ZN(N39910));
    NOR2X1 U27039 (.A1(N8422), .A2(n26652), .ZN(n39911));
    NANDX1 U27040 (.A1(n19259), .A2(N6989), .ZN(N39912));
    INVX1 U27041 (.I(N8378), .ZN(N39913));
    NANDX1 U27042 (.A1(n29598), .A2(N10998), .ZN(N39914));
    NANDX1 U27043 (.A1(n22738), .A2(n25027), .ZN(N39915));
    NANDX1 U27044 (.A1(n19309), .A2(n24425), .ZN(n39916));
    NANDX1 U27045 (.A1(n29532), .A2(N11837), .ZN(N39917));
    NOR2X1 U27046 (.A1(N415), .A2(N12228), .ZN(N39918));
    INVX1 U27047 (.I(N10375), .ZN(n39919));
    NOR2X1 U27048 (.A1(N4693), .A2(N220), .ZN(N39920));
    NANDX1 U27049 (.A1(N10041), .A2(N9758), .ZN(N39921));
    NANDX1 U27050 (.A1(N7024), .A2(N6272), .ZN(N39922));
    NOR2X1 U27051 (.A1(n14843), .A2(n13261), .ZN(N39923));
    NOR2X1 U27052 (.A1(n23220), .A2(N3373), .ZN(N39924));
    INVX1 U27053 (.I(n22778), .ZN(N39925));
    NOR2X1 U27054 (.A1(n28434), .A2(N6228), .ZN(N39926));
    INVX1 U27055 (.I(n17605), .ZN(N39927));
    NOR2X1 U27056 (.A1(N12131), .A2(N5560), .ZN(N39928));
    INVX1 U27057 (.I(N1196), .ZN(N39929));
    NOR2X1 U27058 (.A1(n13140), .A2(n28634), .ZN(N39930));
    NOR2X1 U27059 (.A1(n17112), .A2(n21887), .ZN(N39931));
    NOR2X1 U27060 (.A1(N10864), .A2(n20489), .ZN(n39932));
    NANDX1 U27061 (.A1(N3050), .A2(n27512), .ZN(N39933));
    NANDX1 U27062 (.A1(n13988), .A2(N778), .ZN(n39934));
    NANDX1 U27063 (.A1(n20223), .A2(n23998), .ZN(N39935));
    NANDX1 U27064 (.A1(n25919), .A2(N5199), .ZN(N39936));
    NANDX1 U27065 (.A1(n24215), .A2(N11427), .ZN(n39937));
    NOR2X1 U27066 (.A1(N243), .A2(N502), .ZN(n39938));
    NOR2X1 U27067 (.A1(n24500), .A2(N1414), .ZN(N39939));
    NOR2X1 U27068 (.A1(N336), .A2(N3115), .ZN(N39940));
    NOR2X1 U27069 (.A1(N5244), .A2(n20226), .ZN(n39941));
    NOR2X1 U27070 (.A1(n29069), .A2(N953), .ZN(N39942));
    INVX1 U27071 (.I(n13816), .ZN(n39943));
    NOR2X1 U27072 (.A1(n20540), .A2(n23533), .ZN(N39944));
    NANDX1 U27073 (.A1(n21318), .A2(n16372), .ZN(n39945));
    NANDX1 U27074 (.A1(N3739), .A2(n19843), .ZN(N39946));
    NOR2X1 U27075 (.A1(N8937), .A2(N216), .ZN(n39947));
    NANDX1 U27076 (.A1(N8924), .A2(N3503), .ZN(N39948));
    NOR2X1 U27077 (.A1(n28124), .A2(n18920), .ZN(n39949));
    NANDX1 U27078 (.A1(n18098), .A2(N12654), .ZN(N39950));
    NANDX1 U27079 (.A1(n21212), .A2(N4884), .ZN(N39951));
    NOR2X1 U27080 (.A1(N11301), .A2(n19000), .ZN(N39952));
    NOR2X1 U27081 (.A1(N814), .A2(N12029), .ZN(n39953));
    INVX1 U27082 (.I(n23513), .ZN(N39954));
    INVX1 U27083 (.I(N7339), .ZN(N39955));
    NANDX1 U27084 (.A1(N12309), .A2(N12271), .ZN(N39956));
    INVX1 U27085 (.I(n16047), .ZN(N39957));
    INVX1 U27086 (.I(n26373), .ZN(n39958));
    INVX1 U27087 (.I(N2192), .ZN(N39959));
    NANDX1 U27088 (.A1(N3770), .A2(N5694), .ZN(N39960));
    NANDX1 U27089 (.A1(n20454), .A2(n13174), .ZN(N39961));
    NOR2X1 U27090 (.A1(N8415), .A2(n14388), .ZN(N39962));
    NANDX1 U27091 (.A1(n29626), .A2(n19271), .ZN(N39963));
    NANDX1 U27092 (.A1(N10789), .A2(n26831), .ZN(n39964));
    NANDX1 U27093 (.A1(N11602), .A2(n27420), .ZN(N39965));
    NANDX1 U27094 (.A1(n23676), .A2(n29851), .ZN(N39966));
    NOR2X1 U27095 (.A1(n23601), .A2(N12022), .ZN(n39967));
    NOR2X1 U27096 (.A1(n27420), .A2(n28069), .ZN(N39968));
    NOR2X1 U27097 (.A1(N12216), .A2(N11476), .ZN(N39969));
    NOR2X1 U27098 (.A1(n20903), .A2(N3806), .ZN(n39970));
    NANDX1 U27099 (.A1(N4887), .A2(n24260), .ZN(n39971));
    NOR2X1 U27100 (.A1(n26064), .A2(N2537), .ZN(N39972));
    NANDX1 U27101 (.A1(N5797), .A2(N2025), .ZN(N39973));
    NANDX1 U27102 (.A1(N5425), .A2(N1375), .ZN(N39974));
    NOR2X1 U27103 (.A1(n16619), .A2(N1537), .ZN(N39975));
    INVX1 U27104 (.I(N180), .ZN(N39976));
    NANDX1 U27105 (.A1(N3613), .A2(N9777), .ZN(N39977));
    INVX1 U27106 (.I(N4196), .ZN(N39978));
    INVX1 U27107 (.I(n23216), .ZN(n39979));
    NOR2X1 U27108 (.A1(n13912), .A2(N5295), .ZN(N39980));
    INVX1 U27109 (.I(n17068), .ZN(n39981));
    INVX1 U27110 (.I(n24666), .ZN(N39982));
    NANDX1 U27111 (.A1(n19644), .A2(N7349), .ZN(n39983));
    NANDX1 U27112 (.A1(N4131), .A2(N9885), .ZN(N39984));
    NANDX1 U27113 (.A1(n28625), .A2(N471), .ZN(N39985));
    NOR2X1 U27114 (.A1(N3912), .A2(n20543), .ZN(n39986));
    NOR2X1 U27115 (.A1(N9091), .A2(n22079), .ZN(N39987));
    NANDX1 U27116 (.A1(N9270), .A2(n17154), .ZN(N39988));
    NANDX1 U27117 (.A1(n19046), .A2(n12950), .ZN(n39989));
    NANDX1 U27118 (.A1(N9114), .A2(N6029), .ZN(N39990));
    INVX1 U27119 (.I(n23025), .ZN(N39991));
    NANDX1 U27120 (.A1(n18114), .A2(n28653), .ZN(N39992));
    NANDX1 U27121 (.A1(N1204), .A2(n12994), .ZN(N39993));
    NANDX1 U27122 (.A1(N8552), .A2(n26617), .ZN(N39994));
    INVX1 U27123 (.I(N6998), .ZN(N39995));
    INVX1 U27124 (.I(n25462), .ZN(N39996));
    NANDX1 U27125 (.A1(N11876), .A2(n29374), .ZN(n39997));
    NOR2X1 U27126 (.A1(N6736), .A2(N8327), .ZN(n39998));
    NANDX1 U27127 (.A1(n16934), .A2(N6158), .ZN(N39999));
    INVX1 U27128 (.I(N607), .ZN(n40000));
    NOR2X1 U27129 (.A1(n27176), .A2(N7174), .ZN(N40001));
    NANDX1 U27130 (.A1(n21765), .A2(n23125), .ZN(n40002));
    NOR2X1 U27131 (.A1(n21648), .A2(n29800), .ZN(N40003));
    INVX1 U27132 (.I(N6151), .ZN(n40004));
    NOR2X1 U27133 (.A1(N4395), .A2(n28995), .ZN(N40005));
    NANDX1 U27134 (.A1(n19572), .A2(n25832), .ZN(N40006));
    INVX1 U27135 (.I(N1629), .ZN(N40007));
    NOR2X1 U27136 (.A1(N1003), .A2(N2066), .ZN(N40008));
    NOR2X1 U27137 (.A1(n17573), .A2(N8801), .ZN(N40009));
    NANDX1 U27138 (.A1(n14646), .A2(n25734), .ZN(n40010));
    INVX1 U27139 (.I(n17432), .ZN(N40011));
    NANDX1 U27140 (.A1(n14322), .A2(N3031), .ZN(n40012));
    INVX1 U27141 (.I(n25760), .ZN(N40013));
    INVX1 U27142 (.I(N3623), .ZN(N40014));
    NOR2X1 U27143 (.A1(n16305), .A2(N3285), .ZN(n40015));
    NOR2X1 U27144 (.A1(n22455), .A2(N4150), .ZN(N40016));
    NANDX1 U27145 (.A1(N9873), .A2(N2127), .ZN(N40017));
    NOR2X1 U27146 (.A1(N5567), .A2(N7102), .ZN(n40018));
    NANDX1 U27147 (.A1(n15284), .A2(n26802), .ZN(N40019));
    NOR2X1 U27148 (.A1(N12797), .A2(n14238), .ZN(n40020));
    INVX1 U27149 (.I(N7198), .ZN(n40021));
    NANDX1 U27150 (.A1(N7785), .A2(N7756), .ZN(n40022));
    NOR2X1 U27151 (.A1(n22685), .A2(n22078), .ZN(N40023));
    NOR2X1 U27152 (.A1(N3183), .A2(N6261), .ZN(N40024));
    NOR2X1 U27153 (.A1(n25503), .A2(n24905), .ZN(n40025));
    NOR2X1 U27154 (.A1(n28787), .A2(N4814), .ZN(n40026));
    NOR2X1 U27155 (.A1(n21497), .A2(N7815), .ZN(N40027));
    NOR2X1 U27156 (.A1(n23623), .A2(n18948), .ZN(N40028));
    NANDX1 U27157 (.A1(n19285), .A2(n20271), .ZN(n40029));
    NANDX1 U27158 (.A1(n15950), .A2(n23659), .ZN(n40030));
    NANDX1 U27159 (.A1(n18748), .A2(n24408), .ZN(N40031));
    INVX1 U27160 (.I(N6054), .ZN(N40032));
    NOR2X1 U27161 (.A1(n23764), .A2(N10791), .ZN(n40033));
    NOR2X1 U27162 (.A1(N4265), .A2(n18559), .ZN(n40034));
    INVX1 U27163 (.I(N10525), .ZN(n40035));
    INVX1 U27164 (.I(N409), .ZN(N40036));
    NOR2X1 U27165 (.A1(n16837), .A2(n17756), .ZN(N40037));
    INVX1 U27166 (.I(n16445), .ZN(N40038));
    NANDX1 U27167 (.A1(n25178), .A2(n14487), .ZN(N40039));
    INVX1 U27168 (.I(N2550), .ZN(n40040));
    NOR2X1 U27169 (.A1(n29144), .A2(n22820), .ZN(n40041));
    INVX1 U27170 (.I(n14956), .ZN(n40042));
    INVX1 U27171 (.I(n22919), .ZN(n40043));
    NANDX1 U27172 (.A1(n29310), .A2(N8790), .ZN(N40044));
    NOR2X1 U27173 (.A1(n19926), .A2(n21114), .ZN(n40045));
    NOR2X1 U27174 (.A1(n21787), .A2(n13939), .ZN(N40046));
    INVX1 U27175 (.I(n15391), .ZN(N40047));
    NANDX1 U27176 (.A1(n25635), .A2(N4360), .ZN(N40048));
    NANDX1 U27177 (.A1(N12334), .A2(n22115), .ZN(n40049));
    INVX1 U27178 (.I(n17339), .ZN(n40050));
    INVX1 U27179 (.I(N582), .ZN(N40051));
    NANDX1 U27180 (.A1(N10950), .A2(N3131), .ZN(N40052));
    NANDX1 U27181 (.A1(N9956), .A2(n14512), .ZN(N40053));
    NANDX1 U27182 (.A1(n13472), .A2(n19414), .ZN(N40054));
    NOR2X1 U27183 (.A1(N5598), .A2(N7147), .ZN(N40055));
    INVX1 U27184 (.I(n22475), .ZN(N40056));
    NOR2X1 U27185 (.A1(n18079), .A2(n20006), .ZN(N40057));
    INVX1 U27186 (.I(N1880), .ZN(N40058));
    NANDX1 U27187 (.A1(n22672), .A2(n14903), .ZN(n40059));
    NOR2X1 U27188 (.A1(n27031), .A2(N3080), .ZN(n40060));
    INVX1 U27189 (.I(N7569), .ZN(N40061));
    NANDX1 U27190 (.A1(n26946), .A2(n27358), .ZN(N40062));
    NANDX1 U27191 (.A1(n17195), .A2(n26869), .ZN(N40063));
    NOR2X1 U27192 (.A1(N2661), .A2(n25385), .ZN(N40064));
    NOR2X1 U27193 (.A1(n20934), .A2(N8720), .ZN(n40065));
    NOR2X1 U27194 (.A1(n20549), .A2(N2878), .ZN(N40066));
    NOR2X1 U27195 (.A1(n17514), .A2(n25353), .ZN(n40067));
    NOR2X1 U27196 (.A1(N5455), .A2(n15221), .ZN(N40068));
    NANDX1 U27197 (.A1(N7334), .A2(N9739), .ZN(N40069));
    NOR2X1 U27198 (.A1(n22236), .A2(n29891), .ZN(N40070));
    NANDX1 U27199 (.A1(n13876), .A2(N9361), .ZN(N40071));
    INVX1 U27200 (.I(N11058), .ZN(n40072));
    INVX1 U27201 (.I(n20599), .ZN(N40073));
    INVX1 U27202 (.I(N11925), .ZN(N40074));
    NOR2X1 U27203 (.A1(n16973), .A2(N3146), .ZN(n40075));
    NOR2X1 U27204 (.A1(n28198), .A2(N12640), .ZN(N40076));
    INVX1 U27205 (.I(n28698), .ZN(N40077));
    INVX1 U27206 (.I(N12735), .ZN(N40078));
    NOR2X1 U27207 (.A1(n20564), .A2(n26648), .ZN(n40079));
    NOR2X1 U27208 (.A1(n14579), .A2(N292), .ZN(N40080));
    INVX1 U27209 (.I(n21912), .ZN(N40081));
    NOR2X1 U27210 (.A1(N7251), .A2(N2571), .ZN(N40082));
    NANDX1 U27211 (.A1(N4362), .A2(N5008), .ZN(N40083));
    INVX1 U27212 (.I(n27740), .ZN(N40084));
    NANDX1 U27213 (.A1(n13872), .A2(N6762), .ZN(N40085));
    NOR2X1 U27214 (.A1(n25796), .A2(n24091), .ZN(n40086));
    NOR2X1 U27215 (.A1(n28942), .A2(n25228), .ZN(n40087));
    NOR2X1 U27216 (.A1(N11444), .A2(N4948), .ZN(N40088));
    NOR2X1 U27217 (.A1(N3056), .A2(N6243), .ZN(N40089));
    NANDX1 U27218 (.A1(N12180), .A2(N2753), .ZN(N40090));
    NANDX1 U27219 (.A1(n26759), .A2(N3044), .ZN(N40091));
    NOR2X1 U27220 (.A1(N7094), .A2(N1634), .ZN(N40092));
    INVX1 U27221 (.I(N9665), .ZN(n40093));
    NOR2X1 U27222 (.A1(N1305), .A2(n14672), .ZN(N40094));
    NOR2X1 U27223 (.A1(n17605), .A2(n19297), .ZN(n40095));
    NOR2X1 U27224 (.A1(n24366), .A2(n21303), .ZN(N40096));
    NOR2X1 U27225 (.A1(n18319), .A2(n17403), .ZN(n40097));
    NANDX1 U27226 (.A1(N1971), .A2(n23003), .ZN(n40098));
    INVX1 U27227 (.I(N6918), .ZN(N40099));
    INVX1 U27228 (.I(n26332), .ZN(n40100));
    NOR2X1 U27229 (.A1(N3213), .A2(N8375), .ZN(N40101));
    NANDX1 U27230 (.A1(N8751), .A2(n23694), .ZN(N40102));
    NOR2X1 U27231 (.A1(N9882), .A2(N650), .ZN(N40103));
    NANDX1 U27232 (.A1(N6825), .A2(n29012), .ZN(N40104));
    INVX1 U27233 (.I(N8130), .ZN(n40105));
    INVX1 U27234 (.I(n24063), .ZN(N40106));
    NANDX1 U27235 (.A1(n21403), .A2(N4037), .ZN(N40107));
    NANDX1 U27236 (.A1(N1129), .A2(N9807), .ZN(N40108));
    NOR2X1 U27237 (.A1(n18532), .A2(n21640), .ZN(N40109));
    INVX1 U27238 (.I(n30095), .ZN(n40110));
    NANDX1 U27239 (.A1(N12851), .A2(n15681), .ZN(N40111));
    NANDX1 U27240 (.A1(n14571), .A2(n18893), .ZN(N40112));
    NOR2X1 U27241 (.A1(N7604), .A2(n16204), .ZN(n40113));
    NOR2X1 U27242 (.A1(n22378), .A2(n26086), .ZN(N40114));
    NANDX1 U27243 (.A1(N8648), .A2(n21471), .ZN(N40115));
    NOR2X1 U27244 (.A1(n25031), .A2(n29600), .ZN(N40116));
    NANDX1 U27245 (.A1(N7517), .A2(n13758), .ZN(n40117));
    NANDX1 U27246 (.A1(N11554), .A2(n22281), .ZN(N40118));
    NOR2X1 U27247 (.A1(N9921), .A2(N7546), .ZN(N40119));
    NANDX1 U27248 (.A1(N1424), .A2(n24919), .ZN(N40120));
    INVX1 U27249 (.I(n16203), .ZN(N40121));
    NANDX1 U27250 (.A1(n25478), .A2(n15737), .ZN(n40122));
    NOR2X1 U27251 (.A1(N2794), .A2(N12207), .ZN(n40123));
    NOR2X1 U27252 (.A1(n18998), .A2(N2232), .ZN(N40124));
    INVX1 U27253 (.I(N3507), .ZN(N40125));
    NOR2X1 U27254 (.A1(n19255), .A2(n24977), .ZN(N40126));
    INVX1 U27255 (.I(N2710), .ZN(N40127));
    NANDX1 U27256 (.A1(n22948), .A2(N10226), .ZN(N40128));
    NOR2X1 U27257 (.A1(n24567), .A2(n21779), .ZN(N40129));
    INVX1 U27258 (.I(n15876), .ZN(n40130));
    NOR2X1 U27259 (.A1(n15007), .A2(n25716), .ZN(n40131));
    INVX1 U27260 (.I(n28486), .ZN(n40132));
    INVX1 U27261 (.I(N7749), .ZN(N40133));
    NOR2X1 U27262 (.A1(n19414), .A2(N12046), .ZN(N40134));
    NANDX1 U27263 (.A1(n22208), .A2(n24252), .ZN(n40135));
    INVX1 U27264 (.I(n29766), .ZN(N40136));
    INVX1 U27265 (.I(n22839), .ZN(N40137));
    INVX1 U27266 (.I(N7951), .ZN(N40138));
    NANDX1 U27267 (.A1(n16672), .A2(n27803), .ZN(N40139));
    NOR2X1 U27268 (.A1(n29672), .A2(N9174), .ZN(n40140));
    NOR2X1 U27269 (.A1(n14853), .A2(N3604), .ZN(n40141));
    NANDX1 U27270 (.A1(n22314), .A2(N8040), .ZN(N40142));
    INVX1 U27271 (.I(n25882), .ZN(N40143));
    INVX1 U27272 (.I(n24159), .ZN(N40144));
    NOR2X1 U27273 (.A1(n27692), .A2(n20468), .ZN(N40145));
    NANDX1 U27274 (.A1(n16969), .A2(N2376), .ZN(n40146));
    NOR2X1 U27275 (.A1(n27737), .A2(n15189), .ZN(N40147));
    NANDX1 U27276 (.A1(n15926), .A2(N96), .ZN(N40148));
    INVX1 U27277 (.I(n19060), .ZN(n40149));
    INVX1 U27278 (.I(N6647), .ZN(n40150));
    NOR2X1 U27279 (.A1(n24410), .A2(n28571), .ZN(n40151));
    INVX1 U27280 (.I(N3446), .ZN(N40152));
    NANDX1 U27281 (.A1(n27240), .A2(n25747), .ZN(N40153));
    NOR2X1 U27282 (.A1(n19417), .A2(N3650), .ZN(N40154));
    INVX1 U27283 (.I(N3722), .ZN(N40155));
    NANDX1 U27284 (.A1(n27993), .A2(n16512), .ZN(N40156));
    NOR2X1 U27285 (.A1(n18323), .A2(N12405), .ZN(N40157));
    NOR2X1 U27286 (.A1(N9259), .A2(n25040), .ZN(N40158));
    NOR2X1 U27287 (.A1(n24447), .A2(N8331), .ZN(N40159));
    NANDX1 U27288 (.A1(n24542), .A2(n14461), .ZN(N40160));
    NANDX1 U27289 (.A1(n21149), .A2(N9668), .ZN(N40161));
    NANDX1 U27290 (.A1(N3982), .A2(N8102), .ZN(n40162));
    NOR2X1 U27291 (.A1(N7427), .A2(N8548), .ZN(n40163));
    INVX1 U27292 (.I(n21735), .ZN(N40164));
    NOR2X1 U27293 (.A1(n20238), .A2(n25384), .ZN(n40165));
    NOR2X1 U27294 (.A1(N12520), .A2(n21212), .ZN(N40166));
    INVX1 U27295 (.I(n29032), .ZN(n40167));
    NOR2X1 U27296 (.A1(N7040), .A2(n29997), .ZN(N40168));
    NOR2X1 U27297 (.A1(n16298), .A2(n13460), .ZN(N40169));
    NOR2X1 U27298 (.A1(N10608), .A2(n21791), .ZN(N40170));
    NANDX1 U27299 (.A1(n23710), .A2(n24812), .ZN(N40171));
    INVX1 U27300 (.I(n14721), .ZN(N40172));
    NOR2X1 U27301 (.A1(n25479), .A2(N7263), .ZN(N40173));
    INVX1 U27302 (.I(N10500), .ZN(N40174));
    INVX1 U27303 (.I(N9551), .ZN(n40175));
    INVX1 U27304 (.I(n24985), .ZN(N40176));
    INVX1 U27305 (.I(n20120), .ZN(N40177));
    INVX1 U27306 (.I(N10319), .ZN(N40178));
    NOR2X1 U27307 (.A1(n30003), .A2(N10475), .ZN(N40179));
    NOR2X1 U27308 (.A1(n21718), .A2(n17514), .ZN(N40180));
    INVX1 U27309 (.I(n23784), .ZN(N40181));
    NOR2X1 U27310 (.A1(N3276), .A2(n18181), .ZN(n40182));
    INVX1 U27311 (.I(n13627), .ZN(n40183));
    NANDX1 U27312 (.A1(n26552), .A2(N8301), .ZN(n40184));
    NOR2X1 U27313 (.A1(n29834), .A2(N1204), .ZN(n40185));
    NOR2X1 U27314 (.A1(N6959), .A2(N2207), .ZN(n40186));
    NANDX1 U27315 (.A1(n21648), .A2(N11758), .ZN(n40187));
    NOR2X1 U27316 (.A1(N5056), .A2(N8336), .ZN(N40188));
    NANDX1 U27317 (.A1(n25286), .A2(n18655), .ZN(n40189));
    NANDX1 U27318 (.A1(n13712), .A2(n29129), .ZN(n40190));
    NANDX1 U27319 (.A1(N5293), .A2(n16506), .ZN(N40191));
    NOR2X1 U27320 (.A1(n17637), .A2(N8741), .ZN(N40192));
    NOR2X1 U27321 (.A1(N5680), .A2(N11583), .ZN(n40193));
    NOR2X1 U27322 (.A1(n19253), .A2(N7997), .ZN(n40194));
    NOR2X1 U27323 (.A1(N6699), .A2(N7693), .ZN(n40195));
    INVX1 U27324 (.I(N8184), .ZN(N40196));
    NOR2X1 U27325 (.A1(N4377), .A2(N8729), .ZN(n40197));
    NOR2X1 U27326 (.A1(N4695), .A2(n20596), .ZN(n40198));
    NOR2X1 U27327 (.A1(n13030), .A2(N11006), .ZN(N40199));
    NOR2X1 U27328 (.A1(N1547), .A2(n22616), .ZN(N40200));
    NANDX1 U27329 (.A1(N539), .A2(n24183), .ZN(N40201));
    NOR2X1 U27330 (.A1(N5605), .A2(n22825), .ZN(N40202));
    INVX1 U27331 (.I(n14345), .ZN(n40203));
    INVX1 U27332 (.I(N2930), .ZN(N40204));
    INVX1 U27333 (.I(n28847), .ZN(N40205));
    INVX1 U27334 (.I(N3786), .ZN(N40206));
    NANDX1 U27335 (.A1(n17441), .A2(N40), .ZN(N40207));
    NANDX1 U27336 (.A1(n25624), .A2(N3252), .ZN(N40208));
    INVX1 U27337 (.I(N4216), .ZN(N40209));
    NANDX1 U27338 (.A1(N10916), .A2(n13372), .ZN(N40210));
    NANDX1 U27339 (.A1(n23946), .A2(n24377), .ZN(N40211));
    NANDX1 U27340 (.A1(n25492), .A2(n16855), .ZN(N40212));
    NOR2X1 U27341 (.A1(n14591), .A2(n29598), .ZN(N40213));
    NOR2X1 U27342 (.A1(n20195), .A2(n22285), .ZN(N40214));
    INVX1 U27343 (.I(N4402), .ZN(n40215));
    INVX1 U27344 (.I(n14324), .ZN(N40216));
    INVX1 U27345 (.I(N4160), .ZN(N40217));
    NOR2X1 U27346 (.A1(n22675), .A2(N3836), .ZN(N40218));
    INVX1 U27347 (.I(N11275), .ZN(n40219));
    NANDX1 U27348 (.A1(n26555), .A2(n14526), .ZN(N40220));
    NOR2X1 U27349 (.A1(n19331), .A2(n19758), .ZN(N40221));
    NOR2X1 U27350 (.A1(N2565), .A2(n24769), .ZN(N40222));
    NOR2X1 U27351 (.A1(n15502), .A2(n13267), .ZN(N40223));
    INVX1 U27352 (.I(n20917), .ZN(n40224));
    INVX1 U27353 (.I(N10952), .ZN(N40225));
    NANDX1 U27354 (.A1(n20368), .A2(n19708), .ZN(n40226));
    NANDX1 U27355 (.A1(n20323), .A2(n24109), .ZN(N40227));
    NANDX1 U27356 (.A1(n23208), .A2(N12861), .ZN(n40228));
    NOR2X1 U27357 (.A1(n18137), .A2(n24096), .ZN(N40229));
    NOR2X1 U27358 (.A1(n19067), .A2(n23931), .ZN(N40230));
    NANDX1 U27359 (.A1(n15484), .A2(N8319), .ZN(N40231));
    NANDX1 U27360 (.A1(N4677), .A2(n28076), .ZN(N40232));
    INVX1 U27361 (.I(N7241), .ZN(N40233));
    NANDX1 U27362 (.A1(n17438), .A2(N11303), .ZN(N40234));
    NANDX1 U27363 (.A1(n13799), .A2(N2082), .ZN(n40235));
    NOR2X1 U27364 (.A1(n24750), .A2(n22458), .ZN(N40236));
    NOR2X1 U27365 (.A1(n14320), .A2(N12103), .ZN(N40237));
    INVX1 U27366 (.I(n26990), .ZN(N40238));
    NANDX1 U27367 (.A1(N11501), .A2(n28411), .ZN(N40239));
    NANDX1 U27368 (.A1(n29637), .A2(n22369), .ZN(N40240));
    NOR2X1 U27369 (.A1(N7127), .A2(n16162), .ZN(n40241));
    NANDX1 U27370 (.A1(n22611), .A2(n13041), .ZN(N40242));
    NOR2X1 U27371 (.A1(n27287), .A2(n29677), .ZN(n40243));
    INVX1 U27372 (.I(n23089), .ZN(N40244));
    NANDX1 U27373 (.A1(N4213), .A2(N4254), .ZN(N40245));
    INVX1 U27374 (.I(N6572), .ZN(n40246));
    INVX1 U27375 (.I(n13082), .ZN(N40247));
    NOR2X1 U27376 (.A1(n17354), .A2(n29887), .ZN(N40248));
    NOR2X1 U27377 (.A1(n29457), .A2(n18180), .ZN(N40249));
    NANDX1 U27378 (.A1(N6517), .A2(n18241), .ZN(N40250));
    INVX1 U27379 (.I(n12967), .ZN(n40251));
    INVX1 U27380 (.I(n28817), .ZN(N40252));
    NANDX1 U27381 (.A1(n24867), .A2(N3402), .ZN(N40253));
    NOR2X1 U27382 (.A1(N5901), .A2(N5003), .ZN(N40254));
    NANDX1 U27383 (.A1(n21748), .A2(N4543), .ZN(n40255));
    INVX1 U27384 (.I(N3260), .ZN(n40256));
    NANDX1 U27385 (.A1(n28104), .A2(n26212), .ZN(n40257));
    NOR2X1 U27386 (.A1(N4539), .A2(n21108), .ZN(N40258));
    INVX1 U27387 (.I(n24421), .ZN(N40259));
    NANDX1 U27388 (.A1(n17765), .A2(n17046), .ZN(N40260));
    INVX1 U27389 (.I(N5807), .ZN(N40261));
    NANDX1 U27390 (.A1(n21418), .A2(n24048), .ZN(n40262));
    NOR2X1 U27391 (.A1(N4248), .A2(N211), .ZN(N40263));
    NOR2X1 U27392 (.A1(n26753), .A2(n13638), .ZN(n40264));
    NANDX1 U27393 (.A1(n14552), .A2(N8099), .ZN(n40265));
    NANDX1 U27394 (.A1(N2832), .A2(n29847), .ZN(n40266));
    NANDX1 U27395 (.A1(n26723), .A2(N2969), .ZN(N40267));
    INVX1 U27396 (.I(n24690), .ZN(N40268));
    NANDX1 U27397 (.A1(N10563), .A2(n29228), .ZN(n40269));
    NANDX1 U27398 (.A1(n28578), .A2(n23511), .ZN(N40270));
    NANDX1 U27399 (.A1(n16205), .A2(n29117), .ZN(n40271));
    NANDX1 U27400 (.A1(N10572), .A2(N5503), .ZN(N40272));
    INVX1 U27401 (.I(n23180), .ZN(n40273));
    INVX1 U27402 (.I(n27464), .ZN(N40274));
    NANDX1 U27403 (.A1(N7248), .A2(N12640), .ZN(N40275));
    NANDX1 U27404 (.A1(N10861), .A2(n27191), .ZN(N40276));
    NANDX1 U27405 (.A1(N8038), .A2(n18584), .ZN(n40277));
    INVX1 U27406 (.I(N9757), .ZN(N40278));
    NOR2X1 U27407 (.A1(n13487), .A2(N3947), .ZN(N40279));
    NANDX1 U27408 (.A1(N1091), .A2(N3071), .ZN(N40280));
    NANDX1 U27409 (.A1(N9801), .A2(N1511), .ZN(N40281));
    INVX1 U27410 (.I(n15396), .ZN(N40282));
    NANDX1 U27411 (.A1(N8423), .A2(N5756), .ZN(n40283));
    NANDX1 U27412 (.A1(N2486), .A2(n17533), .ZN(N40284));
    INVX1 U27413 (.I(n28219), .ZN(n40285));
    INVX1 U27414 (.I(n21841), .ZN(n40286));
    INVX1 U27415 (.I(n16059), .ZN(N40287));
    INVX1 U27416 (.I(N4751), .ZN(N40288));
    INVX1 U27417 (.I(n28101), .ZN(N40289));
    INVX1 U27418 (.I(n20257), .ZN(n40290));
    NOR2X1 U27419 (.A1(n22545), .A2(n23986), .ZN(N40291));
    NOR2X1 U27420 (.A1(n15052), .A2(n22268), .ZN(n40292));
    NANDX1 U27421 (.A1(n18122), .A2(n19639), .ZN(n40293));
    INVX1 U27422 (.I(n19632), .ZN(N40294));
    NOR2X1 U27423 (.A1(N6679), .A2(n14468), .ZN(n40295));
    NOR2X1 U27424 (.A1(N995), .A2(n19876), .ZN(N40296));
    NANDX1 U27425 (.A1(n18527), .A2(n18326), .ZN(n40297));
    NOR2X1 U27426 (.A1(n21946), .A2(n28727), .ZN(n40298));
    INVX1 U27427 (.I(n26565), .ZN(N40299));
    INVX1 U27428 (.I(n25271), .ZN(N40300));
    INVX1 U27429 (.I(n21104), .ZN(N40301));
    NANDX1 U27430 (.A1(N6918), .A2(N10887), .ZN(N40302));
    NANDX1 U27431 (.A1(n19465), .A2(N2718), .ZN(N40303));
    NOR2X1 U27432 (.A1(N11595), .A2(n25776), .ZN(n40304));
    INVX1 U27433 (.I(N1096), .ZN(n40305));
    INVX1 U27434 (.I(N118), .ZN(N40306));
    NANDX1 U27435 (.A1(n23737), .A2(n14586), .ZN(N40307));
    NANDX1 U27436 (.A1(n13292), .A2(N4324), .ZN(N40308));
    NANDX1 U27437 (.A1(N1681), .A2(n22649), .ZN(N40309));
    NANDX1 U27438 (.A1(N12187), .A2(N9799), .ZN(n40310));
    NANDX1 U27439 (.A1(N8614), .A2(n14240), .ZN(N40311));
    NOR2X1 U27440 (.A1(n25413), .A2(n23904), .ZN(n40312));
    NANDX1 U27441 (.A1(n20891), .A2(N4654), .ZN(N40313));
    NOR2X1 U27442 (.A1(N10218), .A2(n26069), .ZN(N40314));
    NOR2X1 U27443 (.A1(n21812), .A2(N10269), .ZN(N40315));
    NOR2X1 U27444 (.A1(N11469), .A2(n27327), .ZN(N40316));
    NANDX1 U27445 (.A1(n18767), .A2(N9487), .ZN(n40317));
    INVX1 U27446 (.I(n21993), .ZN(N40318));
    INVX1 U27447 (.I(n17128), .ZN(N40319));
    INVX1 U27448 (.I(n13019), .ZN(N40320));
    INVX1 U27449 (.I(n17583), .ZN(N40321));
    NOR2X1 U27450 (.A1(N7998), .A2(n13357), .ZN(N40322));
    INVX1 U27451 (.I(N10798), .ZN(n40323));
    NOR2X1 U27452 (.A1(n17654), .A2(N4565), .ZN(N40324));
    NANDX1 U27453 (.A1(N8408), .A2(n27916), .ZN(N40325));
    INVX1 U27454 (.I(N7186), .ZN(N40326));
    NOR2X1 U27455 (.A1(N4248), .A2(n28998), .ZN(n40327));
    NOR2X1 U27456 (.A1(n13788), .A2(n29027), .ZN(n40328));
    NOR2X1 U27457 (.A1(n23446), .A2(n17656), .ZN(N40329));
    INVX1 U27458 (.I(N6113), .ZN(N40330));
    INVX1 U27459 (.I(N10552), .ZN(N40331));
    NANDX1 U27460 (.A1(n21702), .A2(n23570), .ZN(N40332));
    NOR2X1 U27461 (.A1(N9147), .A2(N7198), .ZN(N40333));
    NOR2X1 U27462 (.A1(N11065), .A2(n29577), .ZN(N40334));
    NOR2X1 U27463 (.A1(n22588), .A2(n17093), .ZN(N40335));
    NANDX1 U27464 (.A1(n21502), .A2(n14061), .ZN(N40336));
    INVX1 U27465 (.I(n26831), .ZN(n40337));
    INVX1 U27466 (.I(n27925), .ZN(N40338));
    NOR2X1 U27467 (.A1(n27366), .A2(n20464), .ZN(N40339));
    NANDX1 U27468 (.A1(n26255), .A2(n28889), .ZN(n40340));
    INVX1 U27469 (.I(n13773), .ZN(N40341));
    INVX1 U27470 (.I(N9970), .ZN(N40342));
    NANDX1 U27471 (.A1(n15776), .A2(N10331), .ZN(n40343));
    NANDX1 U27472 (.A1(N9209), .A2(N8892), .ZN(N40344));
    NANDX1 U27473 (.A1(n16406), .A2(N4010), .ZN(N40345));
    INVX1 U27474 (.I(n15845), .ZN(N40346));
    NANDX1 U27475 (.A1(n23329), .A2(n21499), .ZN(N40347));
    INVX1 U27476 (.I(n14693), .ZN(N40348));
    INVX1 U27477 (.I(N1606), .ZN(N40349));
    NANDX1 U27478 (.A1(N3790), .A2(n29531), .ZN(N40350));
    INVX1 U27479 (.I(n19716), .ZN(N40351));
    INVX1 U27480 (.I(n30134), .ZN(N40352));
    NOR2X1 U27481 (.A1(N7169), .A2(N3854), .ZN(N40353));
    INVX1 U27482 (.I(N12393), .ZN(N40354));
    NANDX1 U27483 (.A1(n30011), .A2(n28169), .ZN(N40355));
    INVX1 U27484 (.I(N3282), .ZN(n40356));
    INVX1 U27485 (.I(N10166), .ZN(N40357));
    NANDX1 U27486 (.A1(N12206), .A2(N2737), .ZN(N40358));
    NOR2X1 U27487 (.A1(n16612), .A2(N1223), .ZN(n40359));
    INVX1 U27488 (.I(n26671), .ZN(N40360));
    NOR2X1 U27489 (.A1(N1584), .A2(N9214), .ZN(N40361));
    INVX1 U27490 (.I(N1531), .ZN(N40362));
    NOR2X1 U27491 (.A1(n25706), .A2(N9678), .ZN(N40363));
    INVX1 U27492 (.I(N3986), .ZN(N40364));
    INVX1 U27493 (.I(N6976), .ZN(N40365));
    NOR2X1 U27494 (.A1(N2088), .A2(n25142), .ZN(n40366));
    NOR2X1 U27495 (.A1(N4471), .A2(n13576), .ZN(N40367));
    NOR2X1 U27496 (.A1(N5746), .A2(n16857), .ZN(n40368));
    INVX1 U27497 (.I(n15911), .ZN(N40369));
    NANDX1 U27498 (.A1(N6706), .A2(n18647), .ZN(N40370));
    INVX1 U27499 (.I(N11878), .ZN(N40371));
    NANDX1 U27500 (.A1(N9104), .A2(N8411), .ZN(N40372));
    NANDX1 U27501 (.A1(N10688), .A2(n17624), .ZN(N40373));
    NANDX1 U27502 (.A1(N779), .A2(n19188), .ZN(n40374));
    INVX1 U27503 (.I(N10456), .ZN(N40375));
    INVX1 U27504 (.I(N10169), .ZN(N40376));
    NOR2X1 U27505 (.A1(N5867), .A2(n28582), .ZN(N40377));
    INVX1 U27506 (.I(n19569), .ZN(n40378));
    INVX1 U27507 (.I(N3810), .ZN(N40379));
    INVX1 U27508 (.I(n27950), .ZN(n40380));
    NOR2X1 U27509 (.A1(N8424), .A2(n22450), .ZN(N40381));
    NANDX1 U27510 (.A1(N6800), .A2(n17716), .ZN(N40382));
    NANDX1 U27511 (.A1(n29013), .A2(n18154), .ZN(n40383));
    NOR2X1 U27512 (.A1(n26677), .A2(n26564), .ZN(N40384));
    INVX1 U27513 (.I(n25925), .ZN(N40385));
    INVX1 U27514 (.I(N5882), .ZN(N40386));
    NOR2X1 U27515 (.A1(N10360), .A2(N12065), .ZN(n40387));
    INVX1 U27516 (.I(N9251), .ZN(n40388));
    INVX1 U27517 (.I(n22971), .ZN(N40389));
    NANDX1 U27518 (.A1(N9239), .A2(n22310), .ZN(N40390));
    NOR2X1 U27519 (.A1(N8352), .A2(n26119), .ZN(n40391));
    INVX1 U27520 (.I(n24863), .ZN(N40392));
    INVX1 U27521 (.I(n23236), .ZN(N40393));
    INVX1 U27522 (.I(N8122), .ZN(N40394));
    INVX1 U27523 (.I(n23451), .ZN(n40395));
    NOR2X1 U27524 (.A1(n17472), .A2(N11467), .ZN(N40396));
    NOR2X1 U27525 (.A1(n14011), .A2(n26591), .ZN(N40397));
    NOR2X1 U27526 (.A1(N9799), .A2(n17762), .ZN(N40398));
    NOR2X1 U27527 (.A1(n25063), .A2(n28121), .ZN(N40399));
    NOR2X1 U27528 (.A1(n20645), .A2(n25932), .ZN(N40400));
    NOR2X1 U27529 (.A1(n13479), .A2(n29609), .ZN(n40401));
    NOR2X1 U27530 (.A1(n24349), .A2(n22717), .ZN(n40402));
    NOR2X1 U27531 (.A1(n20330), .A2(n26090), .ZN(n40403));
    NOR2X1 U27532 (.A1(N2987), .A2(n19189), .ZN(N40404));
    INVX1 U27533 (.I(n29806), .ZN(N40405));
    INVX1 U27534 (.I(n25754), .ZN(N40406));
    INVX1 U27535 (.I(n25119), .ZN(n40407));
    NANDX1 U27536 (.A1(N4889), .A2(N8992), .ZN(N40408));
    NOR2X1 U27537 (.A1(n24857), .A2(n18790), .ZN(N40409));
    NANDX1 U27538 (.A1(n20569), .A2(n13715), .ZN(N40410));
    NOR2X1 U27539 (.A1(N5467), .A2(n22921), .ZN(n40411));
    INVX1 U27540 (.I(N12599), .ZN(N40412));
    INVX1 U27541 (.I(n21806), .ZN(N40413));
    NOR2X1 U27542 (.A1(n19171), .A2(N2947), .ZN(n40414));
    NANDX1 U27543 (.A1(n28061), .A2(n29036), .ZN(N40415));
    NOR2X1 U27544 (.A1(N910), .A2(n18087), .ZN(N40416));
    INVX1 U27545 (.I(N578), .ZN(N40417));
    NOR2X1 U27546 (.A1(n25301), .A2(n18162), .ZN(N40418));
    NOR2X1 U27547 (.A1(n20944), .A2(N11612), .ZN(n40419));
    NOR2X1 U27548 (.A1(n13041), .A2(N6331), .ZN(N40420));
    NOR2X1 U27549 (.A1(n22899), .A2(n15460), .ZN(N40421));
    NANDX1 U27550 (.A1(n19301), .A2(n20926), .ZN(N40422));
    NANDX1 U27551 (.A1(N11498), .A2(n22085), .ZN(N40423));
    NOR2X1 U27552 (.A1(N3167), .A2(N9477), .ZN(N40424));
    NOR2X1 U27553 (.A1(n24811), .A2(n28850), .ZN(N40425));
    NANDX1 U27554 (.A1(n23709), .A2(n26093), .ZN(n40426));
    NANDX1 U27555 (.A1(N220), .A2(n25639), .ZN(N40427));
    INVX1 U27556 (.I(n25953), .ZN(N40428));
    INVX1 U27557 (.I(n25182), .ZN(n40429));
    NANDX1 U27558 (.A1(N170), .A2(N6656), .ZN(n40430));
    NANDX1 U27559 (.A1(n13210), .A2(n12986), .ZN(n40431));
    INVX1 U27560 (.I(n24669), .ZN(n40432));
    NANDX1 U27561 (.A1(N5156), .A2(n13832), .ZN(N40433));
    NOR2X1 U27562 (.A1(n14393), .A2(n13891), .ZN(N40434));
    NANDX1 U27563 (.A1(N7013), .A2(N5618), .ZN(N40435));
    NOR2X1 U27564 (.A1(n18803), .A2(N291), .ZN(N40436));
    NOR2X1 U27565 (.A1(n28516), .A2(N12560), .ZN(N40437));
    NANDX1 U27566 (.A1(n16260), .A2(N12779), .ZN(N40438));
    NOR2X1 U27567 (.A1(N4582), .A2(n27293), .ZN(N40439));
    NOR2X1 U27568 (.A1(n29763), .A2(n20945), .ZN(n40440));
    NOR2X1 U27569 (.A1(N6281), .A2(N2727), .ZN(N40441));
    NOR2X1 U27570 (.A1(N7827), .A2(N10126), .ZN(n40442));
    NOR2X1 U27571 (.A1(n13393), .A2(N3843), .ZN(N40443));
    NANDX1 U27572 (.A1(n21186), .A2(N6796), .ZN(N40444));
    INVX1 U27573 (.I(N9488), .ZN(N40445));
    NOR2X1 U27574 (.A1(N4241), .A2(N7267), .ZN(N40446));
    NANDX1 U27575 (.A1(n23229), .A2(n22455), .ZN(N40447));
    INVX1 U27576 (.I(N5651), .ZN(n40448));
    NANDX1 U27577 (.A1(N5673), .A2(N6991), .ZN(n40449));
    INVX1 U27578 (.I(n28952), .ZN(N40450));
    INVX1 U27579 (.I(n14675), .ZN(n40451));
    INVX1 U27580 (.I(n25090), .ZN(N40452));
    NANDX1 U27581 (.A1(n23418), .A2(n27816), .ZN(n40453));
    INVX1 U27582 (.I(n19805), .ZN(N40454));
    INVX1 U27583 (.I(N8261), .ZN(N40455));
    NOR2X1 U27584 (.A1(n18905), .A2(n23131), .ZN(N40456));
    INVX1 U27585 (.I(n25701), .ZN(N40457));
    INVX1 U27586 (.I(N10855), .ZN(N40458));
    NOR2X1 U27587 (.A1(N3116), .A2(N6682), .ZN(N40459));
    INVX1 U27588 (.I(n14905), .ZN(n40460));
    INVX1 U27589 (.I(n19956), .ZN(N40461));
    INVX1 U27590 (.I(N2461), .ZN(N40462));
    NOR2X1 U27591 (.A1(n27545), .A2(N1128), .ZN(n40463));
    NOR2X1 U27592 (.A1(n20251), .A2(n15802), .ZN(N40464));
    NANDX1 U27593 (.A1(n15203), .A2(N5077), .ZN(N40465));
    NOR2X1 U27594 (.A1(N1442), .A2(N12299), .ZN(N40466));
    NOR2X1 U27595 (.A1(n16505), .A2(N9120), .ZN(N40467));
    NOR2X1 U27596 (.A1(N5272), .A2(N2113), .ZN(N40468));
    NOR2X1 U27597 (.A1(N835), .A2(N988), .ZN(N40469));
    INVX1 U27598 (.I(N10206), .ZN(N40470));
    INVX1 U27599 (.I(N12174), .ZN(n40471));
    NANDX1 U27600 (.A1(N7568), .A2(N11173), .ZN(N40472));
    NOR2X1 U27601 (.A1(n28122), .A2(N2194), .ZN(n40473));
    NANDX1 U27602 (.A1(n14091), .A2(N3321), .ZN(N40474));
    NOR2X1 U27603 (.A1(N4204), .A2(n19123), .ZN(n40475));
    INVX1 U27604 (.I(n19407), .ZN(n40476));
    INVX1 U27605 (.I(n28170), .ZN(N40477));
    NOR2X1 U27606 (.A1(n25058), .A2(n18381), .ZN(N40478));
    NANDX1 U27607 (.A1(n22738), .A2(N11652), .ZN(N40479));
    NOR2X1 U27608 (.A1(n24850), .A2(N6289), .ZN(n40480));
    NOR2X1 U27609 (.A1(n14398), .A2(N11781), .ZN(N40481));
    INVX1 U27610 (.I(N7061), .ZN(n40482));
    NANDX1 U27611 (.A1(N11260), .A2(n14628), .ZN(N40483));
    INVX1 U27612 (.I(N250), .ZN(N40484));
    INVX1 U27613 (.I(n25882), .ZN(n40485));
    NANDX1 U27614 (.A1(n15264), .A2(n17763), .ZN(N40486));
    INVX1 U27615 (.I(n19467), .ZN(n40487));
    NANDX1 U27616 (.A1(n24361), .A2(n27434), .ZN(N40488));
    NOR2X1 U27617 (.A1(n22393), .A2(N6706), .ZN(N40489));
    NANDX1 U27618 (.A1(n29335), .A2(N2481), .ZN(N40490));
    NANDX1 U27619 (.A1(N10849), .A2(n22226), .ZN(N40491));
    INVX1 U27620 (.I(n17137), .ZN(N40492));
    INVX1 U27621 (.I(N11959), .ZN(N40493));
    NOR2X1 U27622 (.A1(n24756), .A2(N7580), .ZN(N40494));
    NANDX1 U27623 (.A1(n24576), .A2(n22208), .ZN(N40495));
    NOR2X1 U27624 (.A1(n24825), .A2(n23381), .ZN(n40496));
    NANDX1 U27625 (.A1(n28254), .A2(N8507), .ZN(N40497));
    INVX1 U27626 (.I(n17729), .ZN(N40498));
    NANDX1 U27627 (.A1(N9481), .A2(N11952), .ZN(N40499));
    NOR2X1 U27628 (.A1(n17549), .A2(n22906), .ZN(N40500));
    NANDX1 U27629 (.A1(n27797), .A2(n22103), .ZN(n40501));
    NOR2X1 U27630 (.A1(N508), .A2(n21512), .ZN(N40502));
    INVX1 U27631 (.I(n28205), .ZN(n40503));
    NOR2X1 U27632 (.A1(n27773), .A2(n28724), .ZN(n40504));
    NOR2X1 U27633 (.A1(N10952), .A2(N6167), .ZN(N40505));
    NANDX1 U27634 (.A1(N5390), .A2(n28374), .ZN(N40506));
    NANDX1 U27635 (.A1(n18775), .A2(N10178), .ZN(N40507));
    NOR2X1 U27636 (.A1(n16892), .A2(n18684), .ZN(n40508));
    INVX1 U27637 (.I(n23181), .ZN(N40509));
    NANDX1 U27638 (.A1(n20616), .A2(n23694), .ZN(N40510));
    INVX1 U27639 (.I(n26725), .ZN(N40511));
    NANDX1 U27640 (.A1(n28006), .A2(n24384), .ZN(n40512));
    NANDX1 U27641 (.A1(N9446), .A2(n24891), .ZN(N40513));
    NANDX1 U27642 (.A1(n13111), .A2(N11520), .ZN(N40514));
    NANDX1 U27643 (.A1(n29444), .A2(N10106), .ZN(n40515));
    NOR2X1 U27644 (.A1(n28956), .A2(n16272), .ZN(N40516));
    NANDX1 U27645 (.A1(N4208), .A2(N3069), .ZN(N40517));
    NOR2X1 U27646 (.A1(N11543), .A2(n13246), .ZN(N40518));
    INVX1 U27647 (.I(n28434), .ZN(n40519));
    INVX1 U27648 (.I(N160), .ZN(n40520));
    NOR2X1 U27649 (.A1(n14131), .A2(n20775), .ZN(n40521));
    NOR2X1 U27650 (.A1(N2903), .A2(n17363), .ZN(N40522));
    NANDX1 U27651 (.A1(n19470), .A2(N170), .ZN(N40523));
    INVX1 U27652 (.I(n28915), .ZN(n40524));
    NOR2X1 U27653 (.A1(N1224), .A2(N11888), .ZN(N40525));
    NOR2X1 U27654 (.A1(n16793), .A2(n29892), .ZN(N40526));
    NOR2X1 U27655 (.A1(N5336), .A2(n28710), .ZN(N40527));
    INVX1 U27656 (.I(n19724), .ZN(N40528));
    NOR2X1 U27657 (.A1(N1571), .A2(N11786), .ZN(n40529));
    INVX1 U27658 (.I(n14817), .ZN(N40530));
    NOR2X1 U27659 (.A1(n19878), .A2(n23867), .ZN(N40531));
    INVX1 U27660 (.I(n18477), .ZN(n40532));
    NOR2X1 U27661 (.A1(N10306), .A2(N10632), .ZN(N40533));
    NANDX1 U27662 (.A1(n16229), .A2(N7809), .ZN(n40534));
    NOR2X1 U27663 (.A1(n16399), .A2(N1973), .ZN(N40535));
    INVX1 U27664 (.I(n30020), .ZN(n40536));
    NANDX1 U27665 (.A1(N6579), .A2(n25023), .ZN(N40537));
    NOR2X1 U27666 (.A1(N6333), .A2(n30131), .ZN(n40538));
    NANDX1 U27667 (.A1(n23603), .A2(n28633), .ZN(n40539));
    INVX1 U27668 (.I(N3504), .ZN(n40540));
    NANDX1 U27669 (.A1(N3817), .A2(N6386), .ZN(n40541));
    INVX1 U27670 (.I(n23326), .ZN(N40542));
    NANDX1 U27671 (.A1(n27310), .A2(N12857), .ZN(n40543));
    NOR2X1 U27672 (.A1(n23731), .A2(n23162), .ZN(N40544));
    NOR2X1 U27673 (.A1(N11615), .A2(N9254), .ZN(N40545));
    NANDX1 U27674 (.A1(n18968), .A2(n14213), .ZN(N40546));
    NANDX1 U27675 (.A1(n25098), .A2(n14095), .ZN(N40547));
    NOR2X1 U27676 (.A1(N1539), .A2(n27678), .ZN(n40548));
    INVX1 U27677 (.I(n26569), .ZN(N40549));
    INVX1 U27678 (.I(N3446), .ZN(N40550));
    NANDX1 U27679 (.A1(n14728), .A2(n14175), .ZN(N40551));
    NANDX1 U27680 (.A1(n14794), .A2(N6552), .ZN(N40552));
    NOR2X1 U27681 (.A1(n18237), .A2(n29877), .ZN(N40553));
    NANDX1 U27682 (.A1(N3970), .A2(N12596), .ZN(N40554));
    INVX1 U27683 (.I(n16261), .ZN(n40555));
    NANDX1 U27684 (.A1(N4507), .A2(n27875), .ZN(n40556));
    INVX1 U27685 (.I(n14669), .ZN(N40557));
    NANDX1 U27686 (.A1(n17647), .A2(n15365), .ZN(N40558));
    NANDX1 U27687 (.A1(n20302), .A2(N7816), .ZN(n40559));
    NANDX1 U27688 (.A1(n17842), .A2(N8816), .ZN(N40560));
    NOR2X1 U27689 (.A1(N3936), .A2(N822), .ZN(N40561));
    INVX1 U27690 (.I(n18663), .ZN(N40562));
    NOR2X1 U27691 (.A1(n26145), .A2(n22017), .ZN(N40563));
    INVX1 U27692 (.I(N3052), .ZN(N40564));
    NOR2X1 U27693 (.A1(N9848), .A2(n13480), .ZN(N40565));
    NOR2X1 U27694 (.A1(N11005), .A2(n15631), .ZN(N40566));
    NOR2X1 U27695 (.A1(N5186), .A2(n20137), .ZN(N40567));
    INVX1 U27696 (.I(N8620), .ZN(N40568));
    NOR2X1 U27697 (.A1(n21910), .A2(n14827), .ZN(n40569));
    NANDX1 U27698 (.A1(N10697), .A2(n23689), .ZN(n40570));
    NOR2X1 U27699 (.A1(N1021), .A2(N11393), .ZN(N40571));
    NOR2X1 U27700 (.A1(n25173), .A2(N3889), .ZN(n40572));
    INVX1 U27701 (.I(N9083), .ZN(N40573));
    NANDX1 U27702 (.A1(n18164), .A2(n23789), .ZN(N40574));
    INVX1 U27703 (.I(n28272), .ZN(N40575));
    NANDX1 U27704 (.A1(N1669), .A2(n26680), .ZN(n40576));
    NOR2X1 U27705 (.A1(n23013), .A2(N7547), .ZN(N40577));
    INVX1 U27706 (.I(N343), .ZN(N40578));
    INVX1 U27707 (.I(n23071), .ZN(N40579));
    INVX1 U27708 (.I(N9912), .ZN(n40580));
    INVX1 U27709 (.I(n16019), .ZN(n40581));
    NOR2X1 U27710 (.A1(n24893), .A2(n26715), .ZN(n40582));
    NOR2X1 U27711 (.A1(N11164), .A2(n16296), .ZN(N40583));
    NANDX1 U27712 (.A1(n13510), .A2(N11331), .ZN(n40584));
    NOR2X1 U27713 (.A1(n16678), .A2(n20414), .ZN(N40585));
    NANDX1 U27714 (.A1(n23402), .A2(N2626), .ZN(n40586));
    NANDX1 U27715 (.A1(n21536), .A2(n18026), .ZN(N40587));
    NOR2X1 U27716 (.A1(N6639), .A2(n16768), .ZN(n40588));
    NOR2X1 U27717 (.A1(N2747), .A2(n19701), .ZN(N40589));
    INVX1 U27718 (.I(n15478), .ZN(N40590));
    INVX1 U27719 (.I(N2350), .ZN(N40591));
    INVX1 U27720 (.I(n28933), .ZN(N40592));
    NANDX1 U27721 (.A1(n15810), .A2(n23688), .ZN(n40593));
    NOR2X1 U27722 (.A1(n22660), .A2(N4715), .ZN(N40594));
    NOR2X1 U27723 (.A1(n18023), .A2(N6785), .ZN(N40595));
    INVX1 U27724 (.I(n17275), .ZN(N40596));
    INVX1 U27725 (.I(n28667), .ZN(n40597));
    INVX1 U27726 (.I(n16726), .ZN(N40598));
    INVX1 U27727 (.I(n29556), .ZN(N40599));
    NANDX1 U27728 (.A1(n19180), .A2(N3003), .ZN(n40600));
    INVX1 U27729 (.I(n24508), .ZN(N40601));
    INVX1 U27730 (.I(n24768), .ZN(N40602));
    NANDX1 U27731 (.A1(N3524), .A2(N10108), .ZN(n40603));
    NANDX1 U27732 (.A1(n24571), .A2(N12619), .ZN(N40604));
    NANDX1 U27733 (.A1(N1363), .A2(n28429), .ZN(N40605));
    NANDX1 U27734 (.A1(N4868), .A2(N9512), .ZN(n40606));
    NANDX1 U27735 (.A1(N1791), .A2(n27534), .ZN(N40607));
    INVX1 U27736 (.I(n21484), .ZN(N40608));
    INVX1 U27737 (.I(N996), .ZN(n40609));
    NANDX1 U27738 (.A1(N734), .A2(N6283), .ZN(N40610));
    INVX1 U27739 (.I(N152), .ZN(n40611));
    INVX1 U27740 (.I(n28908), .ZN(N40612));
    NANDX1 U27741 (.A1(n24988), .A2(n23279), .ZN(N40613));
    NANDX1 U27742 (.A1(n19618), .A2(n25911), .ZN(N40614));
    INVX1 U27743 (.I(n18287), .ZN(N40615));
    NOR2X1 U27744 (.A1(n26530), .A2(n19466), .ZN(N40616));
    INVX1 U27745 (.I(n27892), .ZN(N40617));
    INVX1 U27746 (.I(N2575), .ZN(N40618));
    NOR2X1 U27747 (.A1(n15829), .A2(N3461), .ZN(N40619));
    NOR2X1 U27748 (.A1(N1787), .A2(n29830), .ZN(N40620));
    INVX1 U27749 (.I(N5019), .ZN(N40621));
    INVX1 U27750 (.I(n23031), .ZN(n40622));
    INVX1 U27751 (.I(n25669), .ZN(n40623));
    INVX1 U27752 (.I(n13163), .ZN(n40624));
    INVX1 U27753 (.I(n20090), .ZN(n40625));
    NANDX1 U27754 (.A1(N12047), .A2(N1792), .ZN(N40626));
    NOR2X1 U27755 (.A1(n20225), .A2(n16263), .ZN(N40627));
    INVX1 U27756 (.I(n27072), .ZN(n40628));
    INVX1 U27757 (.I(n20363), .ZN(n40629));
    NOR2X1 U27758 (.A1(N10825), .A2(n18118), .ZN(N40630));
    INVX1 U27759 (.I(N1960), .ZN(N40631));
    INVX1 U27760 (.I(N8410), .ZN(N40632));
    NOR2X1 U27761 (.A1(n20972), .A2(n28894), .ZN(N40633));
    NANDX1 U27762 (.A1(n23990), .A2(N3775), .ZN(N40634));
    NANDX1 U27763 (.A1(N5444), .A2(n16785), .ZN(n40635));
    INVX1 U27764 (.I(n26763), .ZN(N40636));
    NANDX1 U27765 (.A1(n25787), .A2(N5276), .ZN(N40637));
    NOR2X1 U27766 (.A1(n26394), .A2(N7068), .ZN(n40638));
    NOR2X1 U27767 (.A1(N5042), .A2(N11891), .ZN(n40639));
    NOR2X1 U27768 (.A1(N1977), .A2(N9055), .ZN(N40640));
    INVX1 U27769 (.I(N6938), .ZN(n40641));
    NOR2X1 U27770 (.A1(N5996), .A2(n18216), .ZN(N40642));
    INVX1 U27771 (.I(n22555), .ZN(n40643));
    INVX1 U27772 (.I(N4381), .ZN(n40644));
    INVX1 U27773 (.I(n13942), .ZN(N40645));
    NOR2X1 U27774 (.A1(n25939), .A2(N6277), .ZN(n40646));
    INVX1 U27775 (.I(N1245), .ZN(N40647));
    NOR2X1 U27776 (.A1(N8266), .A2(n16568), .ZN(N40648));
    NANDX1 U27777 (.A1(n22613), .A2(n21844), .ZN(N40649));
    NOR2X1 U27778 (.A1(N7430), .A2(n28911), .ZN(N40650));
    NANDX1 U27779 (.A1(N12471), .A2(N10664), .ZN(n40651));
    NOR2X1 U27780 (.A1(N3008), .A2(N8280), .ZN(n40652));
    NOR2X1 U27781 (.A1(n28643), .A2(n16720), .ZN(n40653));
    INVX1 U27782 (.I(n16722), .ZN(N40654));
    NANDX1 U27783 (.A1(N11140), .A2(N1770), .ZN(N40655));
    NOR2X1 U27784 (.A1(n13089), .A2(n15712), .ZN(n40656));
    NOR2X1 U27785 (.A1(n27589), .A2(n21988), .ZN(N40657));
    NOR2X1 U27786 (.A1(n28833), .A2(n14912), .ZN(N40658));
    NOR2X1 U27787 (.A1(N3825), .A2(n14905), .ZN(N40659));
    NANDX1 U27788 (.A1(n25668), .A2(N8145), .ZN(n40660));
    NANDX1 U27789 (.A1(n13002), .A2(N5204), .ZN(N40661));
    NOR2X1 U27790 (.A1(N12226), .A2(n30053), .ZN(N40662));
    NOR2X1 U27791 (.A1(n20505), .A2(N12643), .ZN(n40663));
    NANDX1 U27792 (.A1(n25785), .A2(N1228), .ZN(N40664));
    NANDX1 U27793 (.A1(N11328), .A2(N928), .ZN(N40665));
    NOR2X1 U27794 (.A1(N1251), .A2(N2578), .ZN(n40666));
    NOR2X1 U27795 (.A1(n19365), .A2(N29), .ZN(n40667));
    NANDX1 U27796 (.A1(N7016), .A2(n17422), .ZN(N40668));
    NOR2X1 U27797 (.A1(N2933), .A2(n21246), .ZN(n40669));
    NOR2X1 U27798 (.A1(N10022), .A2(n16776), .ZN(N40670));
    NOR2X1 U27799 (.A1(n13102), .A2(n29777), .ZN(N40671));
    NANDX1 U27800 (.A1(n28652), .A2(N11866), .ZN(n40672));
    INVX1 U27801 (.I(N5633), .ZN(N40673));
    NANDX1 U27802 (.A1(n22944), .A2(n22696), .ZN(n40674));
    INVX1 U27803 (.I(N12732), .ZN(N40675));
    NOR2X1 U27804 (.A1(n16467), .A2(n13660), .ZN(N40676));
    INVX1 U27805 (.I(n17717), .ZN(N40677));
    NANDX1 U27806 (.A1(n18570), .A2(n25642), .ZN(N40678));
    NOR2X1 U27807 (.A1(N8670), .A2(N2520), .ZN(n40679));
    INVX1 U27808 (.I(n13682), .ZN(N40680));
    NOR2X1 U27809 (.A1(N1917), .A2(n22158), .ZN(N40681));
    NANDX1 U27810 (.A1(N7253), .A2(N8642), .ZN(N40682));
    NANDX1 U27811 (.A1(n25591), .A2(n19027), .ZN(N40683));
    INVX1 U27812 (.I(n26017), .ZN(N40684));
    INVX1 U27813 (.I(N9843), .ZN(N40685));
    INVX1 U27814 (.I(n22133), .ZN(N40686));
    NANDX1 U27815 (.A1(N10510), .A2(N4728), .ZN(N40687));
    NANDX1 U27816 (.A1(n26976), .A2(N6948), .ZN(N40688));
    NOR2X1 U27817 (.A1(N3116), .A2(N11745), .ZN(n40689));
    NOR2X1 U27818 (.A1(n28757), .A2(N5131), .ZN(n40690));
    NANDX1 U27819 (.A1(n19838), .A2(n15938), .ZN(N40691));
    NOR2X1 U27820 (.A1(n13850), .A2(N6415), .ZN(n40692));
    NOR2X1 U27821 (.A1(N6445), .A2(n13668), .ZN(N40693));
    NANDX1 U27822 (.A1(N702), .A2(n27819), .ZN(N40694));
    NOR2X1 U27823 (.A1(N4912), .A2(n23698), .ZN(N40695));
    INVX1 U27824 (.I(N3316), .ZN(N40696));
    NANDX1 U27825 (.A1(N5165), .A2(n12976), .ZN(N40697));
    INVX1 U27826 (.I(N9892), .ZN(N40698));
    INVX1 U27827 (.I(n24977), .ZN(N40699));
    NANDX1 U27828 (.A1(n17969), .A2(n16654), .ZN(N40700));
    NANDX1 U27829 (.A1(n16968), .A2(N3834), .ZN(N40701));
    INVX1 U27830 (.I(n24636), .ZN(N40702));
    NANDX1 U27831 (.A1(n15333), .A2(N4410), .ZN(n40703));
    NANDX1 U27832 (.A1(n21748), .A2(N6341), .ZN(n40704));
    INVX1 U27833 (.I(n23976), .ZN(n40705));
    INVX1 U27834 (.I(N3091), .ZN(n40706));
    INVX1 U27835 (.I(N755), .ZN(n40707));
    NANDX1 U27836 (.A1(N3778), .A2(n25362), .ZN(N40708));
    NANDX1 U27837 (.A1(N2708), .A2(N389), .ZN(N40709));
    NOR2X1 U27838 (.A1(N709), .A2(n28978), .ZN(N40710));
    NANDX1 U27839 (.A1(n14247), .A2(n22938), .ZN(N40711));
    NANDX1 U27840 (.A1(n19461), .A2(n28642), .ZN(N40712));
    NANDX1 U27841 (.A1(n23294), .A2(n28037), .ZN(N40713));
    INVX1 U27842 (.I(N5389), .ZN(N40714));
    NOR2X1 U27843 (.A1(N8341), .A2(N1333), .ZN(N40715));
    NANDX1 U27844 (.A1(N3242), .A2(n22419), .ZN(N40716));
    NANDX1 U27845 (.A1(n27413), .A2(n25509), .ZN(n40717));
    NANDX1 U27846 (.A1(n16728), .A2(N10633), .ZN(n40718));
    NANDX1 U27847 (.A1(N514), .A2(n29208), .ZN(N40719));
    NANDX1 U27848 (.A1(n19600), .A2(n19183), .ZN(N40720));
    INVX1 U27849 (.I(N7002), .ZN(N40721));
    INVX1 U27850 (.I(n26157), .ZN(N40722));
    NANDX1 U27851 (.A1(N9025), .A2(n15480), .ZN(N40723));
    INVX1 U27852 (.I(n18458), .ZN(N40724));
    INVX1 U27853 (.I(n14904), .ZN(n40725));
    INVX1 U27854 (.I(n21283), .ZN(n40726));
    NANDX1 U27855 (.A1(N593), .A2(n22615), .ZN(n40727));
    NOR2X1 U27856 (.A1(n22532), .A2(n14897), .ZN(N40728));
    INVX1 U27857 (.I(N8369), .ZN(N40729));
    INVX1 U27858 (.I(n24936), .ZN(n40730));
    INVX1 U27859 (.I(N9461), .ZN(N40731));
    INVX1 U27860 (.I(n14170), .ZN(N40732));
    INVX1 U27861 (.I(n18675), .ZN(N40733));
    NANDX1 U27862 (.A1(n16275), .A2(N448), .ZN(n40734));
    INVX1 U27863 (.I(N9955), .ZN(N40735));
    NOR2X1 U27864 (.A1(n29133), .A2(n18979), .ZN(N40736));
    INVX1 U27865 (.I(n16000), .ZN(n40737));
    NOR2X1 U27866 (.A1(n16401), .A2(n19465), .ZN(N40738));
    NOR2X1 U27867 (.A1(n26245), .A2(n24722), .ZN(N40739));
    INVX1 U27868 (.I(n18722), .ZN(N40740));
    NANDX1 U27869 (.A1(n29933), .A2(n22179), .ZN(n40741));
    NOR2X1 U27870 (.A1(N8164), .A2(n21008), .ZN(N40742));
    INVX1 U27871 (.I(n21820), .ZN(n40743));
    NANDX1 U27872 (.A1(n18814), .A2(n24551), .ZN(N40744));
    NANDX1 U27873 (.A1(n26049), .A2(n28183), .ZN(n40745));
    NANDX1 U27874 (.A1(n15057), .A2(n27377), .ZN(N40746));
    NANDX1 U27875 (.A1(N84), .A2(n14933), .ZN(N40747));
    INVX1 U27876 (.I(n19288), .ZN(N40748));
    NOR2X1 U27877 (.A1(N4171), .A2(n24250), .ZN(N40749));
    NOR2X1 U27878 (.A1(N10980), .A2(n20357), .ZN(N40750));
    INVX1 U27879 (.I(n18380), .ZN(n40751));
    NANDX1 U27880 (.A1(n15348), .A2(N6736), .ZN(n40752));
    NANDX1 U27881 (.A1(n24632), .A2(N3460), .ZN(n40753));
    NOR2X1 U27882 (.A1(n28714), .A2(n13841), .ZN(n40754));
    NANDX1 U27883 (.A1(N5951), .A2(N8254), .ZN(n40755));
    NANDX1 U27884 (.A1(N1863), .A2(N6299), .ZN(N40756));
    NOR2X1 U27885 (.A1(n16919), .A2(n22236), .ZN(N40757));
    NOR2X1 U27886 (.A1(N5564), .A2(N7031), .ZN(N40758));
    INVX1 U27887 (.I(n24851), .ZN(n40759));
    NOR2X1 U27888 (.A1(N11276), .A2(n18963), .ZN(N40760));
    NANDX1 U27889 (.A1(n22255), .A2(n27880), .ZN(N40761));
    NOR2X1 U27890 (.A1(n29195), .A2(n25382), .ZN(N40762));
    NANDX1 U27891 (.A1(n24492), .A2(N3486), .ZN(N40763));
    NANDX1 U27892 (.A1(n27951), .A2(N2597), .ZN(n40764));
    NOR2X1 U27893 (.A1(N11654), .A2(n27995), .ZN(n40765));
    NOR2X1 U27894 (.A1(N8468), .A2(N9240), .ZN(N40766));
    NOR2X1 U27895 (.A1(N3327), .A2(N2), .ZN(N40767));
    INVX1 U27896 (.I(n25562), .ZN(N40768));
    INVX1 U27897 (.I(N8826), .ZN(N40769));
    NOR2X1 U27898 (.A1(n28777), .A2(N3540), .ZN(N40770));
    NANDX1 U27899 (.A1(N9915), .A2(N11063), .ZN(N40771));
    INVX1 U27900 (.I(N2032), .ZN(N40772));
    NOR2X1 U27901 (.A1(N11559), .A2(n19788), .ZN(N40773));
    NOR2X1 U27902 (.A1(n19898), .A2(n14142), .ZN(n40774));
    INVX1 U27903 (.I(N4034), .ZN(N40775));
    NANDX1 U27904 (.A1(n17390), .A2(n24141), .ZN(N40776));
    NOR2X1 U27905 (.A1(n15247), .A2(n20062), .ZN(n40777));
    INVX1 U27906 (.I(n24487), .ZN(N40778));
    INVX1 U27907 (.I(N12525), .ZN(N40779));
    INVX1 U27908 (.I(N9669), .ZN(N40780));
    NOR2X1 U27909 (.A1(n23282), .A2(n18494), .ZN(n40781));
    NOR2X1 U27910 (.A1(n21921), .A2(N10594), .ZN(n40782));
    NOR2X1 U27911 (.A1(N1699), .A2(N10218), .ZN(n40783));
    NOR2X1 U27912 (.A1(n22428), .A2(n19023), .ZN(n40784));
    INVX1 U27913 (.I(N12078), .ZN(n40785));
    INVX1 U27914 (.I(n20770), .ZN(N40786));
    NOR2X1 U27915 (.A1(n26426), .A2(n24803), .ZN(N40787));
    NANDX1 U27916 (.A1(N2239), .A2(N7368), .ZN(N40788));
    INVX1 U27917 (.I(n17485), .ZN(N40789));
    NANDX1 U27918 (.A1(n25223), .A2(N395), .ZN(N40790));
    INVX1 U27919 (.I(N7610), .ZN(N40791));
    NANDX1 U27920 (.A1(n13366), .A2(n15559), .ZN(n40792));
    NOR2X1 U27921 (.A1(n20420), .A2(n21782), .ZN(N40793));
    INVX1 U27922 (.I(N877), .ZN(N40794));
    NANDX1 U27923 (.A1(N7328), .A2(N11094), .ZN(N40795));
    NANDX1 U27924 (.A1(n29755), .A2(n18677), .ZN(n40796));
    NANDX1 U27925 (.A1(N257), .A2(n18870), .ZN(N40797));
    NANDX1 U27926 (.A1(n15036), .A2(N3719), .ZN(N40798));
    NOR2X1 U27927 (.A1(N194), .A2(n24655), .ZN(n40799));
    NOR2X1 U27928 (.A1(n16219), .A2(N563), .ZN(n40800));
    NANDX1 U27929 (.A1(N11305), .A2(N958), .ZN(N40801));
    NOR2X1 U27930 (.A1(n18914), .A2(N2961), .ZN(n40802));
    NANDX1 U27931 (.A1(n23033), .A2(n28246), .ZN(n40803));
    NOR2X1 U27932 (.A1(n14678), .A2(n15177), .ZN(N40804));
    INVX1 U27933 (.I(N7207), .ZN(N40805));
    NOR2X1 U27934 (.A1(n29382), .A2(N490), .ZN(n40806));
    INVX1 U27935 (.I(N6482), .ZN(n40807));
    NANDX1 U27936 (.A1(N10938), .A2(n13912), .ZN(n40808));
    NOR2X1 U27937 (.A1(n25974), .A2(N6191), .ZN(N40809));
    NOR2X1 U27938 (.A1(n26167), .A2(N708), .ZN(N40810));
    NOR2X1 U27939 (.A1(N810), .A2(N1271), .ZN(N40811));
    NANDX1 U27940 (.A1(N12114), .A2(n20926), .ZN(n40812));
    INVX1 U27941 (.I(N890), .ZN(N40813));
    NOR2X1 U27942 (.A1(n15364), .A2(N12484), .ZN(n40814));
    NANDX1 U27943 (.A1(N2640), .A2(n27161), .ZN(n40815));
    NANDX1 U27944 (.A1(n20928), .A2(n22928), .ZN(N40816));
    NANDX1 U27945 (.A1(N8734), .A2(n23417), .ZN(n40817));
    NOR2X1 U27946 (.A1(n15215), .A2(n18061), .ZN(n40818));
    INVX1 U27947 (.I(n17688), .ZN(n40819));
    INVX1 U27948 (.I(N1235), .ZN(n40820));
    INVX1 U27949 (.I(N12468), .ZN(n40821));
    NOR2X1 U27950 (.A1(n13147), .A2(n14265), .ZN(N40822));
    NOR2X1 U27951 (.A1(N2978), .A2(n26129), .ZN(N40823));
    INVX1 U27952 (.I(N12464), .ZN(n40824));
    INVX1 U27953 (.I(N6896), .ZN(n40825));
    NOR2X1 U27954 (.A1(n18287), .A2(n19379), .ZN(N40826));
    NANDX1 U27955 (.A1(n20926), .A2(N4963), .ZN(N40827));
    INVX1 U27956 (.I(N11717), .ZN(N40828));
    NOR2X1 U27957 (.A1(N3399), .A2(n20450), .ZN(N40829));
    INVX1 U27958 (.I(N9299), .ZN(N40830));
    INVX1 U27959 (.I(n27791), .ZN(N40831));
    NANDX1 U27960 (.A1(N336), .A2(n13843), .ZN(N40832));
    INVX1 U27961 (.I(N12775), .ZN(N40833));
    INVX1 U27962 (.I(N9016), .ZN(N40834));
    NOR2X1 U27963 (.A1(n29135), .A2(n14348), .ZN(n40835));
    NOR2X1 U27964 (.A1(n13688), .A2(N1656), .ZN(N40836));
    NOR2X1 U27965 (.A1(n28050), .A2(n27249), .ZN(N40837));
    NANDX1 U27966 (.A1(n16199), .A2(N5052), .ZN(N40838));
    INVX1 U27967 (.I(N6988), .ZN(N40839));
    INVX1 U27968 (.I(n26762), .ZN(N40840));
    NANDX1 U27969 (.A1(n26465), .A2(N23), .ZN(N40841));
    INVX1 U27970 (.I(N6059), .ZN(n40842));
    NOR2X1 U27971 (.A1(N10362), .A2(N3712), .ZN(N40843));
    NANDX1 U27972 (.A1(N10698), .A2(N6115), .ZN(N40844));
    NOR2X1 U27973 (.A1(n23472), .A2(n20986), .ZN(N40845));
    NOR2X1 U27974 (.A1(N7816), .A2(N8544), .ZN(N40846));
    NOR2X1 U27975 (.A1(n13835), .A2(n22231), .ZN(n40847));
    INVX1 U27976 (.I(n13619), .ZN(n40848));
    NOR2X1 U27977 (.A1(n23580), .A2(n26873), .ZN(N40849));
    NOR2X1 U27978 (.A1(n28631), .A2(n15318), .ZN(N40850));
    NOR2X1 U27979 (.A1(N8507), .A2(N11942), .ZN(n40851));
    INVX1 U27980 (.I(n23533), .ZN(N40852));
    NOR2X1 U27981 (.A1(N2413), .A2(n29591), .ZN(n40853));
    NOR2X1 U27982 (.A1(N1335), .A2(n21863), .ZN(N40854));
    INVX1 U27983 (.I(N593), .ZN(N40855));
    NANDX1 U27984 (.A1(N12434), .A2(n24064), .ZN(N40856));
    INVX1 U27985 (.I(N4201), .ZN(N40857));
    NOR2X1 U27986 (.A1(n23189), .A2(N10316), .ZN(N40858));
    INVX1 U27987 (.I(N3844), .ZN(N40859));
    NOR2X1 U27988 (.A1(n17755), .A2(N12547), .ZN(N40860));
    NOR2X1 U27989 (.A1(N3052), .A2(n14571), .ZN(N40861));
    NOR2X1 U27990 (.A1(n18369), .A2(n23582), .ZN(N40862));
    NANDX1 U27991 (.A1(n18871), .A2(n28418), .ZN(N40863));
    INVX1 U27992 (.I(N7956), .ZN(n40864));
    NOR2X1 U27993 (.A1(N7195), .A2(n25059), .ZN(N40865));
    NANDX1 U27994 (.A1(n17618), .A2(N1724), .ZN(N40866));
    INVX1 U27995 (.I(N4019), .ZN(n40867));
    NANDX1 U27996 (.A1(N3806), .A2(n30103), .ZN(N40868));
    NOR2X1 U27997 (.A1(n24245), .A2(n23155), .ZN(N40869));
    INVX1 U27998 (.I(n16943), .ZN(N40870));
    INVX1 U27999 (.I(N12440), .ZN(N40871));
    NANDX1 U28000 (.A1(n28105), .A2(N12528), .ZN(N40872));
    NOR2X1 U28001 (.A1(N12539), .A2(n29806), .ZN(n40873));
    NANDX1 U28002 (.A1(n24681), .A2(n25454), .ZN(n40874));
    NANDX1 U28003 (.A1(n22962), .A2(N3058), .ZN(N40875));
    NANDX1 U28004 (.A1(N776), .A2(n28950), .ZN(N40876));
    NANDX1 U28005 (.A1(n21501), .A2(n16431), .ZN(n40877));
    NOR2X1 U28006 (.A1(N1243), .A2(n20449), .ZN(N40878));
    INVX1 U28007 (.I(N5048), .ZN(N40879));
    NANDX1 U28008 (.A1(n13328), .A2(n17853), .ZN(N40880));
    INVX1 U28009 (.I(N424), .ZN(n40881));
    NOR2X1 U28010 (.A1(n17551), .A2(N1425), .ZN(n40882));
    NOR2X1 U28011 (.A1(N4079), .A2(n13952), .ZN(n40883));
    NANDX1 U28012 (.A1(n16617), .A2(N2181), .ZN(n40884));
    INVX1 U28013 (.I(n29859), .ZN(n40885));
    INVX1 U28014 (.I(n26280), .ZN(N40886));
    NANDX1 U28015 (.A1(N7814), .A2(n26069), .ZN(n40887));
    NOR2X1 U28016 (.A1(N6627), .A2(n28037), .ZN(N40888));
    INVX1 U28017 (.I(N11618), .ZN(n40889));
    NOR2X1 U28018 (.A1(n23323), .A2(n20627), .ZN(n40890));
    NANDX1 U28019 (.A1(n16931), .A2(n29602), .ZN(n40891));
    NANDX1 U28020 (.A1(N4646), .A2(n20155), .ZN(N40892));
    INVX1 U28021 (.I(n28002), .ZN(N40893));
    NOR2X1 U28022 (.A1(n23177), .A2(n14341), .ZN(n40894));
    INVX1 U28023 (.I(n25689), .ZN(n40895));
    INVX1 U28024 (.I(N5385), .ZN(N40896));
    NOR2X1 U28025 (.A1(n19858), .A2(n23804), .ZN(n40897));
    INVX1 U28026 (.I(n16001), .ZN(n40898));
    INVX1 U28027 (.I(N10302), .ZN(N40899));
    INVX1 U28028 (.I(n16929), .ZN(n40900));
    NOR2X1 U28029 (.A1(n28529), .A2(N8872), .ZN(n40901));
    NOR2X1 U28030 (.A1(n30121), .A2(N2057), .ZN(N40902));
    NOR2X1 U28031 (.A1(n19424), .A2(N7548), .ZN(N40903));
    NOR2X1 U28032 (.A1(n22054), .A2(N12193), .ZN(N40904));
    INVX1 U28033 (.I(n13669), .ZN(N40905));
    NOR2X1 U28034 (.A1(N465), .A2(N6708), .ZN(N40906));
    NANDX1 U28035 (.A1(n19370), .A2(N2259), .ZN(N40907));
    NOR2X1 U28036 (.A1(n24754), .A2(n18689), .ZN(N40908));
    INVX1 U28037 (.I(n18421), .ZN(N40909));
    NOR2X1 U28038 (.A1(n22788), .A2(N11891), .ZN(N40910));
    NANDX1 U28039 (.A1(N11841), .A2(n28819), .ZN(N40911));
    INVX1 U28040 (.I(N10233), .ZN(n40912));
    INVX1 U28041 (.I(N12494), .ZN(N40913));
    NANDX1 U28042 (.A1(n16868), .A2(N8650), .ZN(n40914));
    INVX1 U28043 (.I(n24415), .ZN(N40915));
    NOR2X1 U28044 (.A1(N10116), .A2(n25169), .ZN(n40916));
    NOR2X1 U28045 (.A1(n23785), .A2(n23786), .ZN(N40917));
    NANDX1 U28046 (.A1(n19053), .A2(n25305), .ZN(n40918));
    INVX1 U28047 (.I(n21312), .ZN(N40919));
    NOR2X1 U28048 (.A1(N11616), .A2(n28561), .ZN(N40920));
    NOR2X1 U28049 (.A1(n18597), .A2(N8160), .ZN(n40921));
    NOR2X1 U28050 (.A1(N350), .A2(n28198), .ZN(N40922));
    NANDX1 U28051 (.A1(n17730), .A2(n23586), .ZN(N40923));
    NOR2X1 U28052 (.A1(n13843), .A2(n24641), .ZN(N40924));
    NANDX1 U28053 (.A1(N574), .A2(N3153), .ZN(n40925));
    NANDX1 U28054 (.A1(n13549), .A2(N7422), .ZN(N40926));
    INVX1 U28055 (.I(N8580), .ZN(n40927));
    INVX1 U28056 (.I(n20166), .ZN(n40928));
    NOR2X1 U28057 (.A1(n25095), .A2(N9081), .ZN(N40929));
    NOR2X1 U28058 (.A1(N11956), .A2(n18953), .ZN(N40930));
    NANDX1 U28059 (.A1(n23571), .A2(n17376), .ZN(N40931));
    NANDX1 U28060 (.A1(N12030), .A2(n14097), .ZN(n40932));
    NANDX1 U28061 (.A1(N941), .A2(N12157), .ZN(N40933));
    NANDX1 U28062 (.A1(n18670), .A2(n24303), .ZN(N40934));
    INVX1 U28063 (.I(N2375), .ZN(N40935));
    NANDX1 U28064 (.A1(N7351), .A2(n21646), .ZN(N40936));
    NOR2X1 U28065 (.A1(n23753), .A2(N5058), .ZN(N40937));
    INVX1 U28066 (.I(n20134), .ZN(n40938));
    NOR2X1 U28067 (.A1(n22527), .A2(N10162), .ZN(N40939));
    NANDX1 U28068 (.A1(n17484), .A2(n19243), .ZN(N40940));
    NANDX1 U28069 (.A1(n18000), .A2(n26756), .ZN(n40941));
    NOR2X1 U28070 (.A1(N11434), .A2(n13995), .ZN(N40942));
    NOR2X1 U28071 (.A1(N12024), .A2(n16652), .ZN(n40943));
    INVX1 U28072 (.I(n12964), .ZN(N40944));
    INVX1 U28073 (.I(N8968), .ZN(N40945));
    INVX1 U28074 (.I(n22973), .ZN(N40946));
    INVX1 U28075 (.I(n22569), .ZN(N40947));
    INVX1 U28076 (.I(N2587), .ZN(n40948));
    NOR2X1 U28077 (.A1(N10721), .A2(n14900), .ZN(N40949));
    INVX1 U28078 (.I(n17222), .ZN(N40950));
    NOR2X1 U28079 (.A1(N2634), .A2(N9611), .ZN(n40951));
    NOR2X1 U28080 (.A1(N7059), .A2(n15655), .ZN(n40952));
    NOR2X1 U28081 (.A1(n27578), .A2(N3517), .ZN(n40953));
    NANDX1 U28082 (.A1(n23408), .A2(N3511), .ZN(N40954));
    INVX1 U28083 (.I(N2133), .ZN(N40955));
    NANDX1 U28084 (.A1(n27247), .A2(n20080), .ZN(N40956));
    NANDX1 U28085 (.A1(n25917), .A2(n17608), .ZN(N40957));
    NOR2X1 U28086 (.A1(N7313), .A2(N12844), .ZN(n40958));
    NANDX1 U28087 (.A1(n26213), .A2(n15430), .ZN(N40959));
    NANDX1 U28088 (.A1(N6797), .A2(n18891), .ZN(N40960));
    NOR2X1 U28089 (.A1(n24018), .A2(n23787), .ZN(N40961));
    INVX1 U28090 (.I(N3491), .ZN(N40962));
    NOR2X1 U28091 (.A1(N872), .A2(n19145), .ZN(N40963));
    NOR2X1 U28092 (.A1(n17010), .A2(N11222), .ZN(n40964));
    INVX1 U28093 (.I(n28979), .ZN(N40965));
    NOR2X1 U28094 (.A1(n15886), .A2(n19672), .ZN(n40966));
    NANDX1 U28095 (.A1(N1556), .A2(n28312), .ZN(n40967));
    NOR2X1 U28096 (.A1(n27472), .A2(n15783), .ZN(n40968));
    NOR2X1 U28097 (.A1(n23345), .A2(n17187), .ZN(N40969));
    NANDX1 U28098 (.A1(n19421), .A2(n21178), .ZN(n40970));
    INVX1 U28099 (.I(n14778), .ZN(N40971));
    NOR2X1 U28100 (.A1(n17213), .A2(N8658), .ZN(n40972));
    NOR2X1 U28101 (.A1(N11026), .A2(N709), .ZN(N40973));
    NANDX1 U28102 (.A1(N458), .A2(N8414), .ZN(N40974));
    INVX1 U28103 (.I(N6029), .ZN(n40975));
    NOR2X1 U28104 (.A1(n29344), .A2(N4870), .ZN(n40976));
    NOR2X1 U28105 (.A1(N3653), .A2(n13102), .ZN(n40977));
    INVX1 U28106 (.I(N5208), .ZN(N40978));
    NANDX1 U28107 (.A1(N5928), .A2(N2542), .ZN(N40979));
    NOR2X1 U28108 (.A1(n18791), .A2(n14448), .ZN(n40980));
    NANDX1 U28109 (.A1(n19762), .A2(N3731), .ZN(N40981));
    INVX1 U28110 (.I(n15657), .ZN(n40982));
    NOR2X1 U28111 (.A1(N3639), .A2(N2732), .ZN(N40983));
    NOR2X1 U28112 (.A1(n25916), .A2(N2318), .ZN(N40984));
    NOR2X1 U28113 (.A1(n22583), .A2(N2775), .ZN(n40985));
    INVX1 U28114 (.I(n27938), .ZN(N40986));
    NOR2X1 U28115 (.A1(n21603), .A2(n27145), .ZN(N40987));
    INVX1 U28116 (.I(n14394), .ZN(n40988));
    NOR2X1 U28117 (.A1(n15335), .A2(n14572), .ZN(N40989));
    NANDX1 U28118 (.A1(n15172), .A2(n20499), .ZN(N40990));
    INVX1 U28119 (.I(N12093), .ZN(N40991));
    NANDX1 U28120 (.A1(n30115), .A2(N3322), .ZN(n40992));
    NANDX1 U28121 (.A1(n22406), .A2(n27168), .ZN(N40993));
    NANDX1 U28122 (.A1(n29474), .A2(n19367), .ZN(N40994));
    NOR2X1 U28123 (.A1(N3623), .A2(n15146), .ZN(N40995));
    NANDX1 U28124 (.A1(N8617), .A2(N7591), .ZN(n40996));
    INVX1 U28125 (.I(N10585), .ZN(N40997));
    NOR2X1 U28126 (.A1(N4000), .A2(n20749), .ZN(N40998));
    INVX1 U28127 (.I(n24930), .ZN(N40999));
    NOR2X1 U28128 (.A1(n29015), .A2(n28825), .ZN(N41000));
    INVX1 U28129 (.I(n23443), .ZN(n41001));
    NOR2X1 U28130 (.A1(n28636), .A2(n20412), .ZN(n41002));
    INVX1 U28131 (.I(n14910), .ZN(N41003));
    INVX1 U28132 (.I(n17834), .ZN(n41004));
    INVX1 U28133 (.I(N1219), .ZN(n41005));
    INVX1 U28134 (.I(n23938), .ZN(N41006));
    INVX1 U28135 (.I(N4093), .ZN(n41007));
    NOR2X1 U28136 (.A1(N4178), .A2(N7799), .ZN(N41008));
    INVX1 U28137 (.I(N1356), .ZN(n41009));
    NANDX1 U28138 (.A1(n28719), .A2(N11940), .ZN(N41010));
    NOR2X1 U28139 (.A1(n21279), .A2(n21249), .ZN(n41011));
    NOR2X1 U28140 (.A1(n16072), .A2(n14814), .ZN(N41012));
    INVX1 U28141 (.I(n14759), .ZN(N41013));
    INVX1 U28142 (.I(n18438), .ZN(n41014));
    NOR2X1 U28143 (.A1(N10010), .A2(n27411), .ZN(n41015));
    NOR2X1 U28144 (.A1(n24919), .A2(N6224), .ZN(n41016));
    NOR2X1 U28145 (.A1(n27165), .A2(N7442), .ZN(N41017));
    INVX1 U28146 (.I(N9526), .ZN(N41018));
    INVX1 U28147 (.I(n15464), .ZN(n41019));
    NOR2X1 U28148 (.A1(N736), .A2(N11823), .ZN(N41020));
    NOR2X1 U28149 (.A1(n20789), .A2(N4334), .ZN(N41021));
    INVX1 U28150 (.I(N2591), .ZN(N41022));
    NOR2X1 U28151 (.A1(N5237), .A2(n23840), .ZN(N41023));
    NANDX1 U28152 (.A1(n21308), .A2(N8516), .ZN(N41024));
    INVX1 U28153 (.I(n24627), .ZN(n41025));
    NOR2X1 U28154 (.A1(N7606), .A2(N11668), .ZN(N41026));
    NANDX1 U28155 (.A1(n23577), .A2(N1782), .ZN(N41027));
    NANDX1 U28156 (.A1(n29800), .A2(N9728), .ZN(N41028));
    NOR2X1 U28157 (.A1(n25803), .A2(N2401), .ZN(N41029));
    NOR2X1 U28158 (.A1(N10921), .A2(N6425), .ZN(n41030));
    NOR2X1 U28159 (.A1(N11656), .A2(n18247), .ZN(N41031));
    NANDX1 U28160 (.A1(N2307), .A2(n22580), .ZN(N41032));
    INVX1 U28161 (.I(n23596), .ZN(N41033));
    NOR2X1 U28162 (.A1(N10808), .A2(N5859), .ZN(N41034));
    NOR2X1 U28163 (.A1(n20676), .A2(N2935), .ZN(N41035));
    INVX1 U28164 (.I(n15165), .ZN(N41036));
    NANDX1 U28165 (.A1(n15760), .A2(n15394), .ZN(N41037));
    INVX1 U28166 (.I(n27898), .ZN(N41038));
    INVX1 U28167 (.I(N1921), .ZN(N41039));
    NANDX1 U28168 (.A1(n15463), .A2(N886), .ZN(n41040));
    INVX1 U28169 (.I(n17863), .ZN(N41041));
    INVX1 U28170 (.I(n22707), .ZN(n41042));
    INVX1 U28171 (.I(N11297), .ZN(N41043));
    INVX1 U28172 (.I(N958), .ZN(n41044));
    NOR2X1 U28173 (.A1(n13791), .A2(N12098), .ZN(N41045));
    INVX1 U28174 (.I(n25947), .ZN(N41046));
    INVX1 U28175 (.I(n26411), .ZN(N41047));
    INVX1 U28176 (.I(N2883), .ZN(N41048));
    NANDX1 U28177 (.A1(N4602), .A2(n29735), .ZN(N41049));
    NOR2X1 U28178 (.A1(n16124), .A2(N3918), .ZN(N41050));
    INVX1 U28179 (.I(n16106), .ZN(n41051));
    INVX1 U28180 (.I(N226), .ZN(N41052));
    NOR2X1 U28181 (.A1(n17799), .A2(n15689), .ZN(N41053));
    NOR2X1 U28182 (.A1(n18145), .A2(n22112), .ZN(N41054));
    NOR2X1 U28183 (.A1(N10714), .A2(N4823), .ZN(N41055));
    INVX1 U28184 (.I(n22198), .ZN(n41056));
    INVX1 U28185 (.I(N3860), .ZN(N41057));
    NANDX1 U28186 (.A1(N6438), .A2(n19463), .ZN(n41058));
    NOR2X1 U28187 (.A1(n20471), .A2(n15736), .ZN(N41059));
    NOR2X1 U28188 (.A1(N11914), .A2(n21245), .ZN(N41060));
    NANDX1 U28189 (.A1(N72), .A2(N342), .ZN(n41061));
    INVX1 U28190 (.I(N3990), .ZN(N41062));
    INVX1 U28191 (.I(N5840), .ZN(N41063));
    NANDX1 U28192 (.A1(n25195), .A2(N12426), .ZN(N41064));
    NANDX1 U28193 (.A1(n29444), .A2(N8458), .ZN(N41065));
    INVX1 U28194 (.I(N9980), .ZN(N41066));
    NANDX1 U28195 (.A1(n29445), .A2(N3363), .ZN(N41067));
    NOR2X1 U28196 (.A1(n21505), .A2(n16401), .ZN(N41068));
    NOR2X1 U28197 (.A1(n27355), .A2(n22838), .ZN(N41069));
    INVX1 U28198 (.I(n17575), .ZN(N41070));
    INVX1 U28199 (.I(n19692), .ZN(N41071));
    INVX1 U28200 (.I(N2207), .ZN(N41072));
    INVX1 U28201 (.I(n24649), .ZN(N41073));
    NOR2X1 U28202 (.A1(N11140), .A2(n25822), .ZN(N41074));
    NOR2X1 U28203 (.A1(n24670), .A2(n20222), .ZN(N41075));
    NANDX1 U28204 (.A1(N8289), .A2(N2510), .ZN(N41076));
    INVX1 U28205 (.I(n26293), .ZN(n41077));
    NOR2X1 U28206 (.A1(N8374), .A2(N6135), .ZN(N41078));
    NANDX1 U28207 (.A1(n26379), .A2(n28195), .ZN(N41079));
    INVX1 U28208 (.I(n17747), .ZN(N41080));
    NANDX1 U28209 (.A1(N8660), .A2(N3525), .ZN(N41081));
    NOR2X1 U28210 (.A1(n24055), .A2(n21100), .ZN(n41082));
    INVX1 U28211 (.I(N2170), .ZN(N41083));
    NANDX1 U28212 (.A1(N6917), .A2(n12968), .ZN(N41084));
    NANDX1 U28213 (.A1(n27893), .A2(N12669), .ZN(N41085));
    NANDX1 U28214 (.A1(N11282), .A2(n25899), .ZN(n41086));
    NOR2X1 U28215 (.A1(n19036), .A2(N4050), .ZN(n41087));
    INVX1 U28216 (.I(n27376), .ZN(N41088));
    NOR2X1 U28217 (.A1(N8697), .A2(n24310), .ZN(n41089));
    NANDX1 U28218 (.A1(n17910), .A2(n20551), .ZN(n41090));
    INVX1 U28219 (.I(N500), .ZN(n41091));
    NANDX1 U28220 (.A1(n26114), .A2(n27857), .ZN(n41092));
    NOR2X1 U28221 (.A1(N10394), .A2(n21775), .ZN(N41093));
    INVX1 U28222 (.I(n26543), .ZN(N41094));
    NANDX1 U28223 (.A1(n29027), .A2(N3323), .ZN(N41095));
    NOR2X1 U28224 (.A1(N12523), .A2(n19776), .ZN(N41096));
    INVX1 U28225 (.I(N10400), .ZN(N41097));
    INVX1 U28226 (.I(n22463), .ZN(N41098));
    NOR2X1 U28227 (.A1(N8517), .A2(n15074), .ZN(n41099));
    INVX1 U28228 (.I(N5755), .ZN(N41100));
    INVX1 U28229 (.I(n16226), .ZN(N41101));
    NOR2X1 U28230 (.A1(n28877), .A2(n22697), .ZN(n41102));
    INVX1 U28231 (.I(N10396), .ZN(N41103));
    NOR2X1 U28232 (.A1(N5759), .A2(n25071), .ZN(N41104));
    INVX1 U28233 (.I(N6004), .ZN(N41105));
    NOR2X1 U28234 (.A1(N1113), .A2(n15909), .ZN(N41106));
    INVX1 U28235 (.I(n13618), .ZN(N41107));
    INVX1 U28236 (.I(N12314), .ZN(N41108));
    INVX1 U28237 (.I(n15881), .ZN(n41109));
    NANDX1 U28238 (.A1(N12776), .A2(n26281), .ZN(N41110));
    NANDX1 U28239 (.A1(n23799), .A2(n13203), .ZN(N41111));
    NOR2X1 U28240 (.A1(N8735), .A2(n20732), .ZN(n41112));
    NOR2X1 U28241 (.A1(N1135), .A2(n25519), .ZN(n41113));
    NOR2X1 U28242 (.A1(n18573), .A2(n18078), .ZN(N41114));
    INVX1 U28243 (.I(n28968), .ZN(N41115));
    INVX1 U28244 (.I(N8986), .ZN(n41116));
    NANDX1 U28245 (.A1(N9172), .A2(N3550), .ZN(N41117));
    NOR2X1 U28246 (.A1(N10285), .A2(n19458), .ZN(n41118));
    NOR2X1 U28247 (.A1(N12463), .A2(n22816), .ZN(N41119));
    NANDX1 U28248 (.A1(n28674), .A2(N8560), .ZN(N41120));
    NOR2X1 U28249 (.A1(N11312), .A2(n23401), .ZN(N41121));
    NOR2X1 U28250 (.A1(N4973), .A2(N6466), .ZN(N41122));
    NANDX1 U28251 (.A1(N2269), .A2(n27197), .ZN(N41123));
    NOR2X1 U28252 (.A1(N3403), .A2(N11139), .ZN(N41124));
    NOR2X1 U28253 (.A1(n21975), .A2(n29216), .ZN(n41125));
    INVX1 U28254 (.I(N9367), .ZN(n41126));
    NOR2X1 U28255 (.A1(n28910), .A2(n21828), .ZN(N41127));
    NANDX1 U28256 (.A1(N2322), .A2(n28177), .ZN(N41128));
    NANDX1 U28257 (.A1(N10340), .A2(n13380), .ZN(N41129));
    NANDX1 U28258 (.A1(N3019), .A2(n22335), .ZN(N41130));
    NOR2X1 U28259 (.A1(N139), .A2(n21803), .ZN(N41131));
    NANDX1 U28260 (.A1(n23539), .A2(N12703), .ZN(N41132));
    NANDX1 U28261 (.A1(n30004), .A2(N3551), .ZN(n41133));
    NOR2X1 U28262 (.A1(n15624), .A2(n18800), .ZN(N41134));
    INVX1 U28263 (.I(n26763), .ZN(N41135));
    INVX1 U28264 (.I(N8703), .ZN(N41136));
    INVX1 U28265 (.I(n18026), .ZN(n41137));
    NOR2X1 U28266 (.A1(n13177), .A2(n16799), .ZN(N41138));
    NANDX1 U28267 (.A1(n21123), .A2(N7681), .ZN(N41139));
    NANDX1 U28268 (.A1(n16475), .A2(n18021), .ZN(n41140));
    NANDX1 U28269 (.A1(N5591), .A2(n21039), .ZN(n41141));
    NOR2X1 U28270 (.A1(N11941), .A2(N9738), .ZN(n41142));
    NANDX1 U28271 (.A1(n29602), .A2(N3139), .ZN(n41143));
    NOR2X1 U28272 (.A1(n22098), .A2(n21703), .ZN(N41144));
    NANDX1 U28273 (.A1(N5424), .A2(n25887), .ZN(N41145));
    NANDX1 U28274 (.A1(n22289), .A2(N11073), .ZN(N41146));
    NOR2X1 U28275 (.A1(n19552), .A2(n25475), .ZN(N41147));
    NANDX1 U28276 (.A1(n26182), .A2(N8514), .ZN(N41148));
    NANDX1 U28277 (.A1(n24502), .A2(n18197), .ZN(N41149));
    NANDX1 U28278 (.A1(N9422), .A2(N4534), .ZN(N41150));
    NOR2X1 U28279 (.A1(n26420), .A2(n28822), .ZN(N41151));
    INVX1 U28280 (.I(N5479), .ZN(N41152));
    NOR2X1 U28281 (.A1(N7844), .A2(n25037), .ZN(N41153));
    INVX1 U28282 (.I(n29680), .ZN(N41154));
    NANDX1 U28283 (.A1(N9308), .A2(n21245), .ZN(n41155));
    NOR2X1 U28284 (.A1(n14731), .A2(n16995), .ZN(n41156));
    NANDX1 U28285 (.A1(n25580), .A2(n16628), .ZN(n41157));
    NANDX1 U28286 (.A1(n14995), .A2(N11965), .ZN(n41158));
    INVX1 U28287 (.I(N11039), .ZN(N41159));
    NANDX1 U28288 (.A1(N10476), .A2(n24101), .ZN(N41160));
    NANDX1 U28289 (.A1(N11100), .A2(n22083), .ZN(N41161));
    INVX1 U28290 (.I(n29745), .ZN(N41162));
    NANDX1 U28291 (.A1(N7574), .A2(n27851), .ZN(n41163));
    NANDX1 U28292 (.A1(n18198), .A2(n24256), .ZN(n41164));
    NOR2X1 U28293 (.A1(N5408), .A2(n23798), .ZN(N41165));
    INVX1 U28294 (.I(n14716), .ZN(N41166));
    INVX1 U28295 (.I(N10103), .ZN(N41167));
    INVX1 U28296 (.I(N9022), .ZN(N41168));
    NOR2X1 U28297 (.A1(n13450), .A2(n25649), .ZN(n41169));
    NANDX1 U28298 (.A1(n28444), .A2(N7477), .ZN(N41170));
    NANDX1 U28299 (.A1(n28043), .A2(n16515), .ZN(N41171));
    INVX1 U28300 (.I(n22006), .ZN(N41172));
    NOR2X1 U28301 (.A1(N295), .A2(n13951), .ZN(N41173));
    INVX1 U28302 (.I(n18600), .ZN(N41174));
    INVX1 U28303 (.I(n18637), .ZN(n41175));
    NOR2X1 U28304 (.A1(N3144), .A2(n25395), .ZN(N41176));
    NOR2X1 U28305 (.A1(n29146), .A2(n19364), .ZN(n41177));
    NOR2X1 U28306 (.A1(n29292), .A2(N3942), .ZN(N41178));
    INVX1 U28307 (.I(n27956), .ZN(N41179));
    INVX1 U28308 (.I(n23838), .ZN(n41180));
    INVX1 U28309 (.I(N5260), .ZN(N41181));
    INVX1 U28310 (.I(N10799), .ZN(N41182));
    INVX1 U28311 (.I(n26826), .ZN(N41183));
    INVX1 U28312 (.I(n20169), .ZN(N41184));
    INVX1 U28313 (.I(n27549), .ZN(N41185));
    NANDX1 U28314 (.A1(n22635), .A2(n16404), .ZN(N41186));
    INVX1 U28315 (.I(n22259), .ZN(N41187));
    INVX1 U28316 (.I(n23986), .ZN(n41188));
    INVX1 U28317 (.I(N9741), .ZN(N41189));
    INVX1 U28318 (.I(n13274), .ZN(N41190));
    NOR2X1 U28319 (.A1(n14699), .A2(N2500), .ZN(n41191));
    NOR2X1 U28320 (.A1(N2414), .A2(N6441), .ZN(n41192));
    INVX1 U28321 (.I(N232), .ZN(N41193));
    INVX1 U28322 (.I(n28600), .ZN(N41194));
    NANDX1 U28323 (.A1(n22209), .A2(n17812), .ZN(N41195));
    NOR2X1 U28324 (.A1(n14336), .A2(N3061), .ZN(N41196));
    INVX1 U28325 (.I(n23065), .ZN(n41197));
    INVX1 U28326 (.I(n13251), .ZN(n41198));
    INVX1 U28327 (.I(N4581), .ZN(N41199));
    NOR2X1 U28328 (.A1(n26772), .A2(n26839), .ZN(N41200));
    NOR2X1 U28329 (.A1(N9181), .A2(n14718), .ZN(N41201));
    NOR2X1 U28330 (.A1(N6173), .A2(n27992), .ZN(N41202));
    NOR2X1 U28331 (.A1(N9432), .A2(N354), .ZN(n41203));
    NANDX1 U28332 (.A1(N11846), .A2(n25493), .ZN(N41204));
    NANDX1 U28333 (.A1(N638), .A2(n23744), .ZN(n41205));
    NANDX1 U28334 (.A1(N8903), .A2(N4376), .ZN(n41206));
    INVX1 U28335 (.I(n16526), .ZN(n41207));
    NOR2X1 U28336 (.A1(n21279), .A2(N2229), .ZN(N41208));
    INVX1 U28337 (.I(n14664), .ZN(N41209));
    INVX1 U28338 (.I(N12423), .ZN(N41210));
    NOR2X1 U28339 (.A1(N3557), .A2(n27755), .ZN(N41211));
    NANDX1 U28340 (.A1(n26638), .A2(N6798), .ZN(N41212));
    NOR2X1 U28341 (.A1(N10624), .A2(N1532), .ZN(N41213));
    NANDX1 U28342 (.A1(N10601), .A2(n29661), .ZN(N41214));
    NOR2X1 U28343 (.A1(N11963), .A2(n30067), .ZN(N41215));
    NOR2X1 U28344 (.A1(N6647), .A2(N568), .ZN(N41216));
    INVX1 U28345 (.I(n18492), .ZN(n41217));
    NOR2X1 U28346 (.A1(N6588), .A2(n18012), .ZN(n41218));
    NANDX1 U28347 (.A1(n13860), .A2(N9153), .ZN(N41219));
    NANDX1 U28348 (.A1(N2620), .A2(n23816), .ZN(N41220));
    INVX1 U28349 (.I(n15042), .ZN(n41221));
    INVX1 U28350 (.I(n12941), .ZN(n41222));
    NOR2X1 U28351 (.A1(n13248), .A2(N9442), .ZN(N41223));
    INVX1 U28352 (.I(n21033), .ZN(N41224));
    NOR2X1 U28353 (.A1(n28246), .A2(n15232), .ZN(N41225));
    NOR2X1 U28354 (.A1(n16331), .A2(N9785), .ZN(N41226));
    INVX1 U28355 (.I(n16260), .ZN(N41227));
    NANDX1 U28356 (.A1(n26396), .A2(N5388), .ZN(N41228));
    NANDX1 U28357 (.A1(n14751), .A2(N3418), .ZN(N41229));
    NOR2X1 U28358 (.A1(N2625), .A2(n17974), .ZN(n41230));
    NANDX1 U28359 (.A1(N338), .A2(n23318), .ZN(n41231));
    NANDX1 U28360 (.A1(N12714), .A2(N2565), .ZN(N41232));
    NOR2X1 U28361 (.A1(N2757), .A2(n15506), .ZN(n41233));
    NOR2X1 U28362 (.A1(n16005), .A2(n13508), .ZN(N41234));
    NOR2X1 U28363 (.A1(N6900), .A2(n22133), .ZN(N41235));
    NOR2X1 U28364 (.A1(n22131), .A2(N11222), .ZN(N41236));
    INVX1 U28365 (.I(n20477), .ZN(N41237));
    NANDX1 U28366 (.A1(N11311), .A2(n20169), .ZN(n41238));
    INVX1 U28367 (.I(n16699), .ZN(N41239));
    NOR2X1 U28368 (.A1(N404), .A2(n20116), .ZN(N41240));
    NANDX1 U28369 (.A1(n21726), .A2(n26650), .ZN(n41241));
    INVX1 U28370 (.I(n22063), .ZN(N41242));
    INVX1 U28371 (.I(N9253), .ZN(n41243));
    INVX1 U28372 (.I(N10956), .ZN(N41244));
    NOR2X1 U28373 (.A1(N7395), .A2(n15022), .ZN(n41245));
    NANDX1 U28374 (.A1(n23399), .A2(n17090), .ZN(N41246));
    NANDX1 U28375 (.A1(n18859), .A2(N9086), .ZN(N41247));
    INVX1 U28376 (.I(n29551), .ZN(N41248));
    INVX1 U28377 (.I(n29259), .ZN(N41249));
    INVX1 U28378 (.I(N9702), .ZN(N41250));
    NOR2X1 U28379 (.A1(n28619), .A2(n25492), .ZN(n41251));
    INVX1 U28380 (.I(n27814), .ZN(N41252));
    INVX1 U28381 (.I(N5670), .ZN(N41253));
    NOR2X1 U28382 (.A1(N6044), .A2(n20881), .ZN(n41254));
    NOR2X1 U28383 (.A1(n28106), .A2(n29272), .ZN(N41255));
    NOR2X1 U28384 (.A1(n21305), .A2(n28788), .ZN(N41256));
    NANDX1 U28385 (.A1(n28699), .A2(N2234), .ZN(N41257));
    NOR2X1 U28386 (.A1(N10522), .A2(n19323), .ZN(n41258));
    NANDX1 U28387 (.A1(n17941), .A2(n16969), .ZN(N41259));
    NOR2X1 U28388 (.A1(N5915), .A2(n25837), .ZN(N41260));
    NOR2X1 U28389 (.A1(n25804), .A2(n24099), .ZN(n41261));
    NANDX1 U28390 (.A1(N12847), .A2(N8014), .ZN(N41262));
    NOR2X1 U28391 (.A1(N10523), .A2(n22469), .ZN(N41263));
    NANDX1 U28392 (.A1(n23146), .A2(n17073), .ZN(n41264));
    INVX1 U28393 (.I(N12791), .ZN(N41265));
    NOR2X1 U28394 (.A1(n28719), .A2(N11689), .ZN(N41266));
    NANDX1 U28395 (.A1(n15931), .A2(n25532), .ZN(N41267));
    NANDX1 U28396 (.A1(n18164), .A2(n19659), .ZN(n41268));
    NOR2X1 U28397 (.A1(n26047), .A2(n27696), .ZN(n41269));
    NANDX1 U28398 (.A1(n12879), .A2(N9666), .ZN(n41270));
    INVX1 U28399 (.I(N8578), .ZN(N41271));
    INVX1 U28400 (.I(N7754), .ZN(n41272));
    NANDX1 U28401 (.A1(N8239), .A2(n20600), .ZN(N41273));
    INVX1 U28402 (.I(N11274), .ZN(n41274));
    NANDX1 U28403 (.A1(N10142), .A2(n19979), .ZN(n41275));
    NOR2X1 U28404 (.A1(n15775), .A2(n19426), .ZN(N41276));
    NANDX1 U28405 (.A1(n19376), .A2(N6569), .ZN(n41277));
    INVX1 U28406 (.I(n14144), .ZN(N41278));
    INVX1 U28407 (.I(n21125), .ZN(N41279));
    INVX1 U28408 (.I(n29223), .ZN(N41280));
    INVX1 U28409 (.I(n25842), .ZN(n41281));
    NANDX1 U28410 (.A1(n26902), .A2(n13316), .ZN(N41282));
    NANDX1 U28411 (.A1(n25129), .A2(N6704), .ZN(N41283));
    NOR2X1 U28412 (.A1(n23145), .A2(n14457), .ZN(N41284));
    NANDX1 U28413 (.A1(n19945), .A2(N4919), .ZN(N41285));
    NANDX1 U28414 (.A1(N1081), .A2(n13163), .ZN(N41286));
    INVX1 U28415 (.I(n21059), .ZN(N41287));
    NOR2X1 U28416 (.A1(n16957), .A2(n29046), .ZN(n41288));
    NANDX1 U28417 (.A1(N6195), .A2(n24175), .ZN(N41289));
    NANDX1 U28418 (.A1(N8899), .A2(N5097), .ZN(N41290));
    NOR2X1 U28419 (.A1(n23631), .A2(N4182), .ZN(n41291));
    NOR2X1 U28420 (.A1(n19335), .A2(n17874), .ZN(n41292));
    INVX1 U28421 (.I(N2513), .ZN(N41293));
    NOR2X1 U28422 (.A1(n24697), .A2(N9216), .ZN(N41294));
    NANDX1 U28423 (.A1(n17704), .A2(n23673), .ZN(N41295));
    INVX1 U28424 (.I(N7511), .ZN(N41296));
    NOR2X1 U28425 (.A1(n25167), .A2(n27290), .ZN(N41297));
    NOR2X1 U28426 (.A1(n26350), .A2(n18211), .ZN(n41298));
    INVX1 U28427 (.I(n13169), .ZN(N41299));
    NOR2X1 U28428 (.A1(n12909), .A2(n19364), .ZN(N41300));
    INVX1 U28429 (.I(N6821), .ZN(n41301));
    INVX1 U28430 (.I(N4813), .ZN(N41302));
    NANDX1 U28431 (.A1(n21755), .A2(n27692), .ZN(N41303));
    NANDX1 U28432 (.A1(n29650), .A2(n15429), .ZN(N41304));
    NANDX1 U28433 (.A1(N2025), .A2(n29736), .ZN(N41305));
    INVX1 U28434 (.I(n29939), .ZN(N41306));
    NANDX1 U28435 (.A1(n25052), .A2(n23474), .ZN(n41307));
    NOR2X1 U28436 (.A1(n21123), .A2(n29186), .ZN(n41308));
    NOR2X1 U28437 (.A1(n18275), .A2(n17924), .ZN(N41309));
    NOR2X1 U28438 (.A1(n25047), .A2(n21075), .ZN(N41310));
    NANDX1 U28439 (.A1(N589), .A2(N3846), .ZN(N41311));
    NOR2X1 U28440 (.A1(n19004), .A2(N10666), .ZN(N41312));
    NANDX1 U28441 (.A1(n23816), .A2(n21083), .ZN(N41313));
    NANDX1 U28442 (.A1(N9932), .A2(n15606), .ZN(n41314));
    NOR2X1 U28443 (.A1(n25360), .A2(N9696), .ZN(N41315));
    INVX1 U28444 (.I(n13519), .ZN(N41316));
    INVX1 U28445 (.I(n29397), .ZN(n41317));
    INVX1 U28446 (.I(N11958), .ZN(N41318));
    NOR2X1 U28447 (.A1(N9582), .A2(N2943), .ZN(N41319));
    NANDX1 U28448 (.A1(N4637), .A2(n21218), .ZN(n41320));
    NOR2X1 U28449 (.A1(n14602), .A2(N4688), .ZN(N41321));
    NANDX1 U28450 (.A1(n19037), .A2(n23974), .ZN(N41322));
    INVX1 U28451 (.I(n19958), .ZN(N41323));
    NOR2X1 U28452 (.A1(n22275), .A2(n19003), .ZN(N41324));
    NANDX1 U28453 (.A1(N1781), .A2(n28363), .ZN(N41325));
    INVX1 U28454 (.I(n17386), .ZN(n41326));
    NANDX1 U28455 (.A1(n18931), .A2(n27082), .ZN(n41327));
    NOR2X1 U28456 (.A1(N2312), .A2(n13988), .ZN(n41328));
    NANDX1 U28457 (.A1(N11867), .A2(n14506), .ZN(N41329));
    NOR2X1 U28458 (.A1(n21448), .A2(n17448), .ZN(N41330));
    INVX1 U28459 (.I(n14645), .ZN(N41331));
    NOR2X1 U28460 (.A1(N2703), .A2(n29246), .ZN(n41332));
    INVX1 U28461 (.I(n21905), .ZN(N41333));
    NOR2X1 U28462 (.A1(n25750), .A2(n22074), .ZN(N41334));
    NANDX1 U28463 (.A1(N8452), .A2(n14211), .ZN(n41335));
    NANDX1 U28464 (.A1(n22229), .A2(N4553), .ZN(N41336));
    INVX1 U28465 (.I(n27239), .ZN(N41337));
    NOR2X1 U28466 (.A1(n28112), .A2(N4593), .ZN(n41338));
    NOR2X1 U28467 (.A1(N11791), .A2(n25602), .ZN(N41339));
    INVX1 U28468 (.I(N6168), .ZN(n41340));
    NOR2X1 U28469 (.A1(n24496), .A2(N11839), .ZN(N41341));
    NANDX1 U28470 (.A1(N11807), .A2(n16413), .ZN(N41342));
    NOR2X1 U28471 (.A1(N8895), .A2(n19115), .ZN(N41343));
    NANDX1 U28472 (.A1(N10671), .A2(n29580), .ZN(N41344));
    INVX1 U28473 (.I(n24981), .ZN(n41345));
    NOR2X1 U28474 (.A1(N11447), .A2(N3295), .ZN(n41346));
    INVX1 U28475 (.I(n15536), .ZN(n41347));
    NANDX1 U28476 (.A1(n28840), .A2(n17851), .ZN(N41348));
    NOR2X1 U28477 (.A1(N9202), .A2(N4386), .ZN(N41349));
    NANDX1 U28478 (.A1(n16644), .A2(N4737), .ZN(N41350));
    INVX1 U28479 (.I(n26635), .ZN(n41351));
    NOR2X1 U28480 (.A1(N7135), .A2(n20993), .ZN(N41352));
    INVX1 U28481 (.I(n13036), .ZN(N41353));
    INVX1 U28482 (.I(n16277), .ZN(N41354));
    NANDX1 U28483 (.A1(N118), .A2(n23953), .ZN(N41355));
    INVX1 U28484 (.I(n29486), .ZN(N41356));
    NOR2X1 U28485 (.A1(n26579), .A2(n24329), .ZN(N41357));
    NOR2X1 U28486 (.A1(N7888), .A2(n16184), .ZN(n41358));
    NANDX1 U28487 (.A1(n23424), .A2(N131), .ZN(N41359));
    NANDX1 U28488 (.A1(n29835), .A2(N11317), .ZN(N41360));
    NOR2X1 U28489 (.A1(n22781), .A2(n15656), .ZN(n41361));
    NANDX1 U28490 (.A1(n27517), .A2(n15459), .ZN(N41362));
    NOR2X1 U28491 (.A1(n26981), .A2(N11155), .ZN(N41363));
    NANDX1 U28492 (.A1(N8147), .A2(N12751), .ZN(N41364));
    INVX1 U28493 (.I(n24424), .ZN(n41365));
    NANDX1 U28494 (.A1(n26682), .A2(n18239), .ZN(n41366));
    NANDX1 U28495 (.A1(n26030), .A2(N57), .ZN(N41367));
    INVX1 U28496 (.I(n20221), .ZN(N41368));
    NOR2X1 U28497 (.A1(N9302), .A2(n24965), .ZN(N41369));
    INVX1 U28498 (.I(N2588), .ZN(n41370));
    INVX1 U28499 (.I(n23021), .ZN(N41371));
    NANDX1 U28500 (.A1(N6275), .A2(N5532), .ZN(N41372));
    NANDX1 U28501 (.A1(N10491), .A2(n23384), .ZN(N41373));
    INVX1 U28502 (.I(n14510), .ZN(N41374));
    INVX1 U28503 (.I(N7848), .ZN(N41375));
    NOR2X1 U28504 (.A1(n24239), .A2(N4556), .ZN(N41376));
    NOR2X1 U28505 (.A1(n20666), .A2(n17540), .ZN(N41377));
    INVX1 U28506 (.I(N5771), .ZN(N41378));
    NANDX1 U28507 (.A1(n18004), .A2(N1663), .ZN(N41379));
    NOR2X1 U28508 (.A1(n19417), .A2(N10444), .ZN(N41380));
    NANDX1 U28509 (.A1(n28718), .A2(N5272), .ZN(N41381));
    NANDX1 U28510 (.A1(n19866), .A2(N230), .ZN(N41382));
    NANDX1 U28511 (.A1(N10711), .A2(n25202), .ZN(n41383));
    NANDX1 U28512 (.A1(n24336), .A2(n24253), .ZN(N41384));
    NOR2X1 U28513 (.A1(N5203), .A2(N8625), .ZN(n41385));
    INVX1 U28514 (.I(N1612), .ZN(N41386));
    INVX1 U28515 (.I(n13659), .ZN(N41387));
    NANDX1 U28516 (.A1(n19687), .A2(n22886), .ZN(N41388));
    INVX1 U28517 (.I(n21279), .ZN(N41389));
    NANDX1 U28518 (.A1(n17907), .A2(N9145), .ZN(N41390));
    NOR2X1 U28519 (.A1(N725), .A2(n17122), .ZN(N41391));
    NOR2X1 U28520 (.A1(N5633), .A2(n15703), .ZN(N41392));
    NOR2X1 U28521 (.A1(n18675), .A2(N5431), .ZN(N41393));
    INVX1 U28522 (.I(n13162), .ZN(N41394));
    NOR2X1 U28523 (.A1(n25707), .A2(N1741), .ZN(N41395));
    NOR2X1 U28524 (.A1(N8383), .A2(n13703), .ZN(n41396));
    NANDX1 U28525 (.A1(n17008), .A2(n14562), .ZN(N41397));
    INVX1 U28526 (.I(n28418), .ZN(n41398));
    NOR2X1 U28527 (.A1(n19140), .A2(n17967), .ZN(N41399));
    NANDX1 U28528 (.A1(N1269), .A2(n27806), .ZN(N41400));
    INVX1 U28529 (.I(N7736), .ZN(N41401));
    NOR2X1 U28530 (.A1(n15488), .A2(N8460), .ZN(n41402));
    INVX1 U28531 (.I(N3235), .ZN(N41403));
    NOR2X1 U28532 (.A1(n28198), .A2(n14950), .ZN(N41404));
    INVX1 U28533 (.I(n22189), .ZN(N41405));
    NANDX1 U28534 (.A1(n23050), .A2(N8193), .ZN(N41406));
    INVX1 U28535 (.I(n24791), .ZN(N41407));
    NANDX1 U28536 (.A1(N7969), .A2(N8356), .ZN(n41408));
    INVX1 U28537 (.I(n24976), .ZN(N41409));
    INVX1 U28538 (.I(N12731), .ZN(N41410));
    INVX1 U28539 (.I(n28260), .ZN(n41411));
    INVX1 U28540 (.I(n29783), .ZN(N41412));
    INVX1 U28541 (.I(N3001), .ZN(n41413));
    NOR2X1 U28542 (.A1(n22958), .A2(n29434), .ZN(N41414));
    NANDX1 U28543 (.A1(N8309), .A2(N7756), .ZN(N41415));
    NANDX1 U28544 (.A1(N104), .A2(n29107), .ZN(n41416));
    INVX1 U28545 (.I(N3614), .ZN(N41417));
    NOR2X1 U28546 (.A1(N2554), .A2(n19069), .ZN(N41418));
    NOR2X1 U28547 (.A1(n29444), .A2(n18655), .ZN(N41419));
    NANDX1 U28548 (.A1(n25098), .A2(n15184), .ZN(n41420));
    NOR2X1 U28549 (.A1(n13416), .A2(n28720), .ZN(N41421));
    INVX1 U28550 (.I(n14707), .ZN(n41422));
    NANDX1 U28551 (.A1(N2940), .A2(n16439), .ZN(n41423));
    INVX1 U28552 (.I(n29289), .ZN(N41424));
    INVX1 U28553 (.I(n14617), .ZN(N41425));
    NANDX1 U28554 (.A1(N7296), .A2(n26003), .ZN(N41426));
    INVX1 U28555 (.I(N3613), .ZN(n41427));
    INVX1 U28556 (.I(n19081), .ZN(N41428));
    NANDX1 U28557 (.A1(n18809), .A2(n22695), .ZN(n41429));
    INVX1 U28558 (.I(N9923), .ZN(N41430));
    INVX1 U28559 (.I(N1769), .ZN(N41431));
    NOR2X1 U28560 (.A1(n18841), .A2(n28329), .ZN(N41432));
    INVX1 U28561 (.I(N3887), .ZN(N41433));
    NANDX1 U28562 (.A1(n13425), .A2(N2469), .ZN(N41434));
    NANDX1 U28563 (.A1(n28132), .A2(N1428), .ZN(N41435));
    NANDX1 U28564 (.A1(N2994), .A2(N33), .ZN(n41436));
    NANDX1 U28565 (.A1(N10994), .A2(n14649), .ZN(N41437));
    INVX1 U28566 (.I(N6850), .ZN(N41438));
    NANDX1 U28567 (.A1(n16646), .A2(n29160), .ZN(N41439));
    INVX1 U28568 (.I(n24287), .ZN(N41440));
    NANDX1 U28569 (.A1(n26190), .A2(n16844), .ZN(N41441));
    NANDX1 U28570 (.A1(n24673), .A2(n17031), .ZN(n41442));
    NOR2X1 U28571 (.A1(N11023), .A2(n24432), .ZN(N41443));
    NANDX1 U28572 (.A1(n22471), .A2(n16880), .ZN(n41444));
    NOR2X1 U28573 (.A1(N5759), .A2(N7909), .ZN(N41445));
    NANDX1 U28574 (.A1(n22451), .A2(N9337), .ZN(N41446));
    INVX1 U28575 (.I(n25444), .ZN(n41447));
    NOR2X1 U28576 (.A1(n16199), .A2(n24998), .ZN(n41448));
    NOR2X1 U28577 (.A1(n13866), .A2(N1711), .ZN(n41449));
    NOR2X1 U28578 (.A1(N374), .A2(n19431), .ZN(N41450));
    NOR2X1 U28579 (.A1(n24661), .A2(n28294), .ZN(n41451));
    NANDX1 U28580 (.A1(n30065), .A2(N7018), .ZN(N41452));
    NOR2X1 U28581 (.A1(N5519), .A2(n17648), .ZN(N41453));
    NOR2X1 U28582 (.A1(n29951), .A2(n15030), .ZN(n41454));
    INVX1 U28583 (.I(n16693), .ZN(n41455));
    INVX1 U28584 (.I(n25994), .ZN(N41456));
    NOR2X1 U28585 (.A1(n26597), .A2(n18307), .ZN(N41457));
    INVX1 U28586 (.I(n25660), .ZN(N41458));
    INVX1 U28587 (.I(N1729), .ZN(N41459));
    NANDX1 U28588 (.A1(N8474), .A2(n14307), .ZN(N41460));
    NANDX1 U28589 (.A1(n28882), .A2(N7261), .ZN(N41461));
    NOR2X1 U28590 (.A1(N6736), .A2(n26294), .ZN(N41462));
    NANDX1 U28591 (.A1(N4892), .A2(n29940), .ZN(n41463));
    NANDX1 U28592 (.A1(N11910), .A2(n28121), .ZN(N41464));
    NOR2X1 U28593 (.A1(n29557), .A2(N7187), .ZN(n41465));
    NANDX1 U28594 (.A1(N3011), .A2(n27422), .ZN(N41466));
    NANDX1 U28595 (.A1(n25650), .A2(n23278), .ZN(N41467));
    NANDX1 U28596 (.A1(N10671), .A2(N8), .ZN(n41468));
    NOR2X1 U28597 (.A1(N6193), .A2(n13621), .ZN(n41469));
    NANDX1 U28598 (.A1(n17914), .A2(N10655), .ZN(N41470));
    NOR2X1 U28599 (.A1(N1924), .A2(n28097), .ZN(N41471));
    INVX1 U28600 (.I(n16444), .ZN(n41472));
    NOR2X1 U28601 (.A1(N10212), .A2(N2610), .ZN(N41473));
    NANDX1 U28602 (.A1(n28712), .A2(N142), .ZN(N41474));
    NANDX1 U28603 (.A1(n26695), .A2(n21890), .ZN(n41475));
    INVX1 U28604 (.I(n22442), .ZN(N41476));
    INVX1 U28605 (.I(n19745), .ZN(n41477));
    NANDX1 U28606 (.A1(n28690), .A2(N3819), .ZN(n41478));
    INVX1 U28607 (.I(N8392), .ZN(N41479));
    NOR2X1 U28608 (.A1(N1436), .A2(N10592), .ZN(n41480));
    NOR2X1 U28609 (.A1(N3617), .A2(n14520), .ZN(N41481));
    INVX1 U28610 (.I(N2832), .ZN(n41482));
    NANDX1 U28611 (.A1(n29078), .A2(n19489), .ZN(N41483));
    NANDX1 U28612 (.A1(N3946), .A2(N12744), .ZN(N41484));
    NOR2X1 U28613 (.A1(N6555), .A2(n29589), .ZN(n41485));
    NOR2X1 U28614 (.A1(n25394), .A2(n16767), .ZN(N41486));
    NANDX1 U28615 (.A1(N5707), .A2(N3365), .ZN(n41487));
    INVX1 U28616 (.I(N7582), .ZN(n41488));
    NANDX1 U28617 (.A1(n29864), .A2(n24833), .ZN(N41489));
    INVX1 U28618 (.I(N1155), .ZN(N41490));
    NOR2X1 U28619 (.A1(n18537), .A2(n21288), .ZN(N41491));
    INVX1 U28620 (.I(n27779), .ZN(n41492));
    NOR2X1 U28621 (.A1(n28197), .A2(n13357), .ZN(N41493));
    INVX1 U28622 (.I(n19374), .ZN(N41494));
    INVX1 U28623 (.I(N5647), .ZN(N41495));
    NOR2X1 U28624 (.A1(N4804), .A2(N6951), .ZN(N41496));
    NOR2X1 U28625 (.A1(n30056), .A2(N6403), .ZN(N41497));
    NANDX1 U28626 (.A1(n25312), .A2(N11730), .ZN(n41498));
    INVX1 U28627 (.I(n19579), .ZN(N41499));
    INVX1 U28628 (.I(N3065), .ZN(N41500));
    INVX1 U28629 (.I(n15325), .ZN(n41501));
    NANDX1 U28630 (.A1(N10417), .A2(n19373), .ZN(n41502));
    NANDX1 U28631 (.A1(n13503), .A2(n26471), .ZN(n41503));
    NANDX1 U28632 (.A1(n15742), .A2(N12673), .ZN(N41504));
    INVX1 U28633 (.I(n13801), .ZN(N41505));
    NANDX1 U28634 (.A1(N1976), .A2(N3038), .ZN(N41506));
    NANDX1 U28635 (.A1(N7622), .A2(n27643), .ZN(n41507));
    INVX1 U28636 (.I(n14573), .ZN(n41508));
    NOR2X1 U28637 (.A1(n20169), .A2(N9536), .ZN(n41509));
    NANDX1 U28638 (.A1(n15343), .A2(N9826), .ZN(n41510));
    INVX1 U28639 (.I(n23483), .ZN(N41511));
    INVX1 U28640 (.I(N11718), .ZN(N41512));
    NOR2X1 U28641 (.A1(n17366), .A2(N3069), .ZN(N41513));
    NOR2X1 U28642 (.A1(n25299), .A2(n14273), .ZN(N41514));
    NANDX1 U28643 (.A1(n21632), .A2(n16626), .ZN(N41515));
    NOR2X1 U28644 (.A1(n22865), .A2(N2307), .ZN(n41516));
    NANDX1 U28645 (.A1(n18757), .A2(N4282), .ZN(n41517));
    NANDX1 U28646 (.A1(n15506), .A2(N11904), .ZN(N41518));
    NANDX1 U28647 (.A1(N5620), .A2(n15037), .ZN(N41519));
    NANDX1 U28648 (.A1(n14349), .A2(n13133), .ZN(N41520));
    NANDX1 U28649 (.A1(n18253), .A2(N11519), .ZN(N41521));
    NANDX1 U28650 (.A1(N11598), .A2(n24999), .ZN(N41522));
    INVX1 U28651 (.I(n20664), .ZN(n41523));
    INVX1 U28652 (.I(N7801), .ZN(n41524));
    NOR2X1 U28653 (.A1(n26087), .A2(N10634), .ZN(N41525));
    NANDX1 U28654 (.A1(N6142), .A2(n27260), .ZN(N41526));
    NOR2X1 U28655 (.A1(n29007), .A2(n18127), .ZN(N41527));
    NANDX1 U28656 (.A1(N6187), .A2(n22408), .ZN(N41528));
    NOR2X1 U28657 (.A1(N10253), .A2(n22872), .ZN(N41529));
    NANDX1 U28658 (.A1(N4433), .A2(n26469), .ZN(N41530));
    INVX1 U28659 (.I(n18782), .ZN(N41531));
    NOR2X1 U28660 (.A1(n15454), .A2(N6897), .ZN(N41532));
    NOR2X1 U28661 (.A1(n27167), .A2(n18494), .ZN(n41533));
    NOR2X1 U28662 (.A1(N1762), .A2(n27718), .ZN(n41534));
    INVX1 U28663 (.I(n28260), .ZN(n41535));
    INVX1 U28664 (.I(N8401), .ZN(N41536));
    INVX1 U28665 (.I(n27703), .ZN(N41537));
    INVX1 U28666 (.I(n24577), .ZN(n41538));
    NANDX1 U28667 (.A1(N1972), .A2(N12566), .ZN(n41539));
    NOR2X1 U28668 (.A1(N8158), .A2(n23534), .ZN(N41540));
    NOR2X1 U28669 (.A1(n18411), .A2(n16269), .ZN(N41541));
    NANDX1 U28670 (.A1(n22843), .A2(N12600), .ZN(N41542));
    NOR2X1 U28671 (.A1(N11487), .A2(N10625), .ZN(N41543));
    NANDX1 U28672 (.A1(N6944), .A2(N8729), .ZN(N41544));
    NANDX1 U28673 (.A1(n13998), .A2(N1694), .ZN(N41545));
    NANDX1 U28674 (.A1(N11578), .A2(n25584), .ZN(n41546));
    INVX1 U28675 (.I(n19166), .ZN(N41547));
    INVX1 U28676 (.I(n18817), .ZN(n41548));
    INVX1 U28677 (.I(N6950), .ZN(N41549));
    NOR2X1 U28678 (.A1(N11424), .A2(N8921), .ZN(N41550));
    NOR2X1 U28679 (.A1(N5496), .A2(N5640), .ZN(N41551));
    NOR2X1 U28680 (.A1(N7314), .A2(n24050), .ZN(N41552));
    NOR2X1 U28681 (.A1(n26933), .A2(N5316), .ZN(N41553));
    INVX1 U28682 (.I(n28808), .ZN(N41554));
    NANDX1 U28683 (.A1(n24392), .A2(N4560), .ZN(N41555));
    NOR2X1 U28684 (.A1(N2983), .A2(n26176), .ZN(N41556));
    INVX1 U28685 (.I(n23375), .ZN(n41557));
    NOR2X1 U28686 (.A1(n26443), .A2(n18821), .ZN(N41558));
    INVX1 U28687 (.I(n15472), .ZN(N41559));
    NANDX1 U28688 (.A1(n29595), .A2(n20764), .ZN(N41560));
    INVX1 U28689 (.I(N1275), .ZN(N41561));
    NANDX1 U28690 (.A1(n15659), .A2(N4217), .ZN(N41562));
    NANDX1 U28691 (.A1(n21298), .A2(N11995), .ZN(n41563));
    NANDX1 U28692 (.A1(N3771), .A2(n24602), .ZN(N41564));
    INVX1 U28693 (.I(n27785), .ZN(N41565));
    NOR2X1 U28694 (.A1(N6145), .A2(N3011), .ZN(N41566));
    NOR2X1 U28695 (.A1(n29402), .A2(N3878), .ZN(N41567));
    INVX1 U28696 (.I(n25441), .ZN(N41568));
    NANDX1 U28697 (.A1(n17405), .A2(n14719), .ZN(N41569));
    NOR2X1 U28698 (.A1(n24786), .A2(n25497), .ZN(N41570));
    NANDX1 U28699 (.A1(n24575), .A2(n13516), .ZN(N41571));
    NANDX1 U28700 (.A1(N12615), .A2(n14790), .ZN(N41572));
    INVX1 U28701 (.I(n16835), .ZN(N41573));
    NOR2X1 U28702 (.A1(n15121), .A2(N7995), .ZN(N41574));
    NOR2X1 U28703 (.A1(N7101), .A2(N327), .ZN(N41575));
    INVX1 U28704 (.I(n26013), .ZN(N41576));
    INVX1 U28705 (.I(N10819), .ZN(N41577));
    NANDX1 U28706 (.A1(n19682), .A2(N1867), .ZN(N41578));
    INVX1 U28707 (.I(N12120), .ZN(N41579));
    INVX1 U28708 (.I(n15286), .ZN(N41580));
    INVX1 U28709 (.I(n20560), .ZN(n41581));
    INVX1 U28710 (.I(N4335), .ZN(N41582));
    INVX1 U28711 (.I(n13925), .ZN(N41583));
    NOR2X1 U28712 (.A1(n28344), .A2(n27440), .ZN(N41584));
    INVX1 U28713 (.I(n29519), .ZN(n41585));
    NOR2X1 U28714 (.A1(n29257), .A2(n16216), .ZN(N41586));
    NANDX1 U28715 (.A1(N2801), .A2(N12772), .ZN(N41587));
    NANDX1 U28716 (.A1(N9901), .A2(n13098), .ZN(N41588));
    NOR2X1 U28717 (.A1(n24475), .A2(n29769), .ZN(N41589));
    NANDX1 U28718 (.A1(n15055), .A2(n19313), .ZN(N41590));
    NANDX1 U28719 (.A1(N4900), .A2(N1295), .ZN(N41591));
    NANDX1 U28720 (.A1(N8746), .A2(n20718), .ZN(n41592));
    NOR2X1 U28721 (.A1(N8613), .A2(n13613), .ZN(N41593));
    INVX1 U28722 (.I(N11098), .ZN(n41594));
    INVX1 U28723 (.I(n27164), .ZN(N41595));
    NOR2X1 U28724 (.A1(n24391), .A2(n26545), .ZN(N41596));
    NANDX1 U28725 (.A1(n23511), .A2(N12624), .ZN(N41597));
    INVX1 U28726 (.I(n26311), .ZN(N41598));
    INVX1 U28727 (.I(n14913), .ZN(n41599));
    NOR2X1 U28728 (.A1(n27053), .A2(n15142), .ZN(N41600));
    NANDX1 U28729 (.A1(n15245), .A2(n14750), .ZN(N41601));
    NANDX1 U28730 (.A1(n23118), .A2(N4786), .ZN(n41602));
    NANDX1 U28731 (.A1(n24412), .A2(n20854), .ZN(N41603));
    NANDX1 U28732 (.A1(N3554), .A2(n15906), .ZN(N41604));
    NANDX1 U28733 (.A1(n17166), .A2(n14726), .ZN(n41605));
    INVX1 U28734 (.I(N1178), .ZN(N41606));
    NANDX1 U28735 (.A1(N24), .A2(n25568), .ZN(N41607));
    NANDX1 U28736 (.A1(n27773), .A2(n18941), .ZN(N41608));
    INVX1 U28737 (.I(N3467), .ZN(N41609));
    INVX1 U28738 (.I(n23298), .ZN(n41610));
    NOR2X1 U28739 (.A1(n17009), .A2(N8774), .ZN(n41611));
    NANDX1 U28740 (.A1(n13240), .A2(n24018), .ZN(N41612));
    NOR2X1 U28741 (.A1(n24525), .A2(n16998), .ZN(N41613));
    NOR2X1 U28742 (.A1(n29271), .A2(n29971), .ZN(n41614));
    NOR2X1 U28743 (.A1(N12626), .A2(N3387), .ZN(n41615));
    INVX1 U28744 (.I(n23290), .ZN(N41616));
    INVX1 U28745 (.I(n28645), .ZN(n41617));
    NANDX1 U28746 (.A1(N10290), .A2(n28957), .ZN(n41618));
    NANDX1 U28747 (.A1(n24419), .A2(n25676), .ZN(N41619));
    INVX1 U28748 (.I(N1783), .ZN(n41620));
    INVX1 U28749 (.I(N4601), .ZN(N41621));
    NOR2X1 U28750 (.A1(N5301), .A2(N11540), .ZN(N41622));
    NOR2X1 U28751 (.A1(n14075), .A2(n22181), .ZN(N41623));
    NANDX1 U28752 (.A1(n26653), .A2(n17434), .ZN(n41624));
    INVX1 U28753 (.I(N2075), .ZN(n41625));
    NOR2X1 U28754 (.A1(N6348), .A2(N1908), .ZN(n41626));
    NANDX1 U28755 (.A1(n18973), .A2(n23992), .ZN(n41627));
    NOR2X1 U28756 (.A1(N687), .A2(n21665), .ZN(N41628));
    NANDX1 U28757 (.A1(n15601), .A2(n20516), .ZN(n41629));
    NOR2X1 U28758 (.A1(n19099), .A2(n14797), .ZN(n41630));
    NANDX1 U28759 (.A1(N8794), .A2(n16579), .ZN(n41631));
    NOR2X1 U28760 (.A1(N1955), .A2(N10598), .ZN(N41632));
    NOR2X1 U28761 (.A1(n13494), .A2(N10185), .ZN(N41633));
    NANDX1 U28762 (.A1(n24235), .A2(n23012), .ZN(n41634));
    NANDX1 U28763 (.A1(N11532), .A2(N89), .ZN(n41635));
    INVX1 U28764 (.I(n17565), .ZN(N41636));
    NOR2X1 U28765 (.A1(N8525), .A2(n21612), .ZN(n41637));
    NANDX1 U28766 (.A1(n21077), .A2(n20880), .ZN(N41638));
    INVX1 U28767 (.I(N12605), .ZN(N41639));
    INVX1 U28768 (.I(n18817), .ZN(N41640));
    NANDX1 U28769 (.A1(n22508), .A2(N7778), .ZN(n41641));
    NANDX1 U28770 (.A1(n21899), .A2(N5133), .ZN(N41642));
    NANDX1 U28771 (.A1(n21992), .A2(N7087), .ZN(N41643));
    NOR2X1 U28772 (.A1(N8687), .A2(N9142), .ZN(n41644));
    INVX1 U28773 (.I(n16715), .ZN(N41645));
    NOR2X1 U28774 (.A1(n13696), .A2(N9819), .ZN(N41646));
    NOR2X1 U28775 (.A1(n13784), .A2(n16437), .ZN(n41647));
    NANDX1 U28776 (.A1(N8780), .A2(n13522), .ZN(n41648));
    NANDX1 U28777 (.A1(N11310), .A2(N4462), .ZN(N41649));
    INVX1 U28778 (.I(n25965), .ZN(N41650));
    NANDX1 U28779 (.A1(n29024), .A2(n14644), .ZN(N41651));
    INVX1 U28780 (.I(n21394), .ZN(N41652));
    NOR2X1 U28781 (.A1(N3509), .A2(N1717), .ZN(n41653));
    INVX1 U28782 (.I(n14987), .ZN(N41654));
    INVX1 U28783 (.I(N11762), .ZN(N41655));
    INVX1 U28784 (.I(n20955), .ZN(n41656));
    INVX1 U28785 (.I(n27747), .ZN(N41657));
    INVX1 U28786 (.I(N12703), .ZN(N41658));
    NOR2X1 U28787 (.A1(N5911), .A2(N4594), .ZN(N41659));
    INVX1 U28788 (.I(n22347), .ZN(N41660));
    NOR2X1 U28789 (.A1(n22428), .A2(n24430), .ZN(N41661));
    NANDX1 U28790 (.A1(N3601), .A2(n28891), .ZN(N41662));
    NOR2X1 U28791 (.A1(n29565), .A2(n23078), .ZN(n41663));
    NANDX1 U28792 (.A1(N2633), .A2(n20247), .ZN(N41664));
    INVX1 U28793 (.I(N2176), .ZN(N41665));
    NOR2X1 U28794 (.A1(n24467), .A2(N6851), .ZN(N41666));
    NOR2X1 U28795 (.A1(n18037), .A2(n18612), .ZN(N41667));
    NOR2X1 U28796 (.A1(N8854), .A2(n16637), .ZN(N41668));
    INVX1 U28797 (.I(N4946), .ZN(N41669));
    INVX1 U28798 (.I(n13003), .ZN(N41670));
    NANDX1 U28799 (.A1(n22493), .A2(n26651), .ZN(N41671));
    NANDX1 U28800 (.A1(n25103), .A2(n18942), .ZN(n41672));
    NOR2X1 U28801 (.A1(n28643), .A2(n22542), .ZN(N41673));
    NANDX1 U28802 (.A1(n23854), .A2(N10530), .ZN(N41674));
    NANDX1 U28803 (.A1(N6512), .A2(n13162), .ZN(N41675));
    NOR2X1 U28804 (.A1(n29262), .A2(n15337), .ZN(n41676));
    NANDX1 U28805 (.A1(n23591), .A2(N10748), .ZN(n41677));
    INVX1 U28806 (.I(N51), .ZN(n41678));
    NANDX1 U28807 (.A1(N7247), .A2(n27602), .ZN(N41679));
    INVX1 U28808 (.I(N8945), .ZN(N41680));
    NOR2X1 U28809 (.A1(n22319), .A2(N10509), .ZN(N41681));
    NANDX1 U28810 (.A1(n14674), .A2(N7022), .ZN(n41682));
    INVX1 U28811 (.I(N9640), .ZN(n41683));
    NOR2X1 U28812 (.A1(n16767), .A2(n26843), .ZN(n41684));
    NOR2X1 U28813 (.A1(n20136), .A2(N9120), .ZN(N41685));
    NANDX1 U28814 (.A1(N5006), .A2(N4192), .ZN(n41686));
    INVX1 U28815 (.I(n28820), .ZN(N41687));
    NANDX1 U28816 (.A1(N4380), .A2(n16114), .ZN(n41688));
    NANDX1 U28817 (.A1(n15127), .A2(n19270), .ZN(n41689));
    NANDX1 U28818 (.A1(N2910), .A2(n26516), .ZN(n41690));
    NOR2X1 U28819 (.A1(N7329), .A2(n24022), .ZN(n41691));
    INVX1 U28820 (.I(n18208), .ZN(N41692));
    NOR2X1 U28821 (.A1(n24478), .A2(n21443), .ZN(n41693));
    NANDX1 U28822 (.A1(n25189), .A2(n19643), .ZN(n41694));
    NANDX1 U28823 (.A1(N11818), .A2(n16348), .ZN(N41695));
    NANDX1 U28824 (.A1(n20514), .A2(n25467), .ZN(n41696));
    INVX1 U28825 (.I(n25519), .ZN(N41697));
    INVX1 U28826 (.I(N1969), .ZN(N41698));
    INVX1 U28827 (.I(n21535), .ZN(N41699));
    NOR2X1 U28828 (.A1(n17436), .A2(N6866), .ZN(N41700));
    NANDX1 U28829 (.A1(N6568), .A2(N10945), .ZN(N41701));
    NOR2X1 U28830 (.A1(n21645), .A2(n23927), .ZN(n41702));
    INVX1 U28831 (.I(N4090), .ZN(n41703));
    INVX1 U28832 (.I(n15603), .ZN(n41704));
    INVX1 U28833 (.I(n29479), .ZN(n41705));
    INVX1 U28834 (.I(n19895), .ZN(n41706));
    INVX1 U28835 (.I(n26550), .ZN(N41707));
    INVX1 U28836 (.I(N6210), .ZN(N41708));
    NOR2X1 U28837 (.A1(n18423), .A2(n26723), .ZN(N41709));
    INVX1 U28838 (.I(N8470), .ZN(N41710));
    NOR2X1 U28839 (.A1(n26307), .A2(N10438), .ZN(n41711));
    NOR2X1 U28840 (.A1(n17705), .A2(N5346), .ZN(N41712));
    NOR2X1 U28841 (.A1(n13131), .A2(N3942), .ZN(n41713));
    NANDX1 U28842 (.A1(n24075), .A2(N5447), .ZN(N41714));
    NOR2X1 U28843 (.A1(N6425), .A2(N2841), .ZN(N41715));
    INVX1 U28844 (.I(N11427), .ZN(N41716));
    NOR2X1 U28845 (.A1(n17189), .A2(N10768), .ZN(N41717));
    NOR2X1 U28846 (.A1(n25644), .A2(N5161), .ZN(n41718));
    NANDX1 U28847 (.A1(N11202), .A2(n30068), .ZN(n41719));
    NANDX1 U28848 (.A1(n18185), .A2(n26654), .ZN(N41720));
    NANDX1 U28849 (.A1(n26654), .A2(n25879), .ZN(n41721));
    INVX1 U28850 (.I(n25653), .ZN(n41722));
    NANDX1 U28851 (.A1(N10727), .A2(n19559), .ZN(n41723));
    INVX1 U28852 (.I(n23857), .ZN(N41724));
    NANDX1 U28853 (.A1(N1426), .A2(N6355), .ZN(N41725));
    INVX1 U28854 (.I(N6044), .ZN(N41726));
    INVX1 U28855 (.I(n20348), .ZN(N41727));
    NOR2X1 U28856 (.A1(N1327), .A2(N8653), .ZN(N41728));
    NANDX1 U28857 (.A1(N12095), .A2(n22564), .ZN(n41729));
    NOR2X1 U28858 (.A1(N5816), .A2(N2749), .ZN(n41730));
    NANDX1 U28859 (.A1(N5746), .A2(n25831), .ZN(N41731));
    INVX1 U28860 (.I(n20960), .ZN(N41732));
    INVX1 U28861 (.I(N332), .ZN(N41733));
    NANDX1 U28862 (.A1(N8446), .A2(n25984), .ZN(n41734));
    NOR2X1 U28863 (.A1(n19172), .A2(N3967), .ZN(n41735));
    INVX1 U28864 (.I(N1452), .ZN(N41736));
    NOR2X1 U28865 (.A1(N9990), .A2(n26504), .ZN(N41737));
    NANDX1 U28866 (.A1(n16033), .A2(n16405), .ZN(n41738));
    NANDX1 U28867 (.A1(N647), .A2(n17731), .ZN(n41739));
    NANDX1 U28868 (.A1(N2448), .A2(n18386), .ZN(n41740));
    NANDX1 U28869 (.A1(n29893), .A2(n24201), .ZN(N41741));
    NANDX1 U28870 (.A1(n26963), .A2(n18508), .ZN(n41742));
    INVX1 U28871 (.I(N641), .ZN(N41743));
    INVX1 U28872 (.I(N4370), .ZN(n41744));
    NANDX1 U28873 (.A1(n14592), .A2(N1377), .ZN(N41745));
    NANDX1 U28874 (.A1(n16143), .A2(N9109), .ZN(n41746));
    NOR2X1 U28875 (.A1(n24707), .A2(N10561), .ZN(n41747));
    INVX1 U28876 (.I(n23257), .ZN(n41748));
    NOR2X1 U28877 (.A1(N8769), .A2(N9152), .ZN(N41749));
    NANDX1 U28878 (.A1(N2375), .A2(n28496), .ZN(N41750));
    INVX1 U28879 (.I(N11892), .ZN(N41751));
    INVX1 U28880 (.I(N6432), .ZN(N41752));
    INVX1 U28881 (.I(n19260), .ZN(N41753));
    INVX1 U28882 (.I(n29967), .ZN(N41754));
    INVX1 U28883 (.I(n19003), .ZN(n41755));
    NOR2X1 U28884 (.A1(n23985), .A2(n16893), .ZN(n41756));
    INVX1 U28885 (.I(n24957), .ZN(n41757));
    NOR2X1 U28886 (.A1(n24658), .A2(n29035), .ZN(N41758));
    INVX1 U28887 (.I(n22328), .ZN(N41759));
    INVX1 U28888 (.I(n19318), .ZN(N41760));
    INVX1 U28889 (.I(n23752), .ZN(N41761));
    INVX1 U28890 (.I(n16936), .ZN(n41762));
    NOR2X1 U28891 (.A1(N10150), .A2(n28828), .ZN(N41763));
    NOR2X1 U28892 (.A1(N8508), .A2(n16874), .ZN(N41764));
    NANDX1 U28893 (.A1(n16573), .A2(n23305), .ZN(N41765));
    NOR2X1 U28894 (.A1(N5696), .A2(N12361), .ZN(N41766));
    NANDX1 U28895 (.A1(n29040), .A2(N1226), .ZN(N41767));
    NANDX1 U28896 (.A1(n22887), .A2(N6680), .ZN(N41768));
    NOR2X1 U28897 (.A1(N6268), .A2(n26725), .ZN(N41769));
    INVX1 U28898 (.I(N5165), .ZN(N41770));
    NANDX1 U28899 (.A1(n13461), .A2(N12105), .ZN(n41771));
    INVX1 U28900 (.I(N4772), .ZN(n41772));
    NOR2X1 U28901 (.A1(N11514), .A2(n21707), .ZN(n41773));
    NANDX1 U28902 (.A1(N10224), .A2(N8958), .ZN(n41774));
    NANDX1 U28903 (.A1(N7293), .A2(n14392), .ZN(N41775));
    INVX1 U28904 (.I(n23865), .ZN(N41776));
    NANDX1 U28905 (.A1(n17313), .A2(n18121), .ZN(N41777));
    INVX1 U28906 (.I(n13308), .ZN(N41778));
    INVX1 U28907 (.I(n28405), .ZN(n41779));
    INVX1 U28908 (.I(n28471), .ZN(n41780));
    INVX1 U28909 (.I(N6129), .ZN(N41781));
    NANDX1 U28910 (.A1(n20232), .A2(n15960), .ZN(n41782));
    NANDX1 U28911 (.A1(N11430), .A2(n29420), .ZN(N41783));
    NANDX1 U28912 (.A1(N10507), .A2(n22752), .ZN(n41784));
    INVX1 U28913 (.I(N10582), .ZN(n41785));
    NOR2X1 U28914 (.A1(N8632), .A2(n20805), .ZN(N41786));
    NOR2X1 U28915 (.A1(N5871), .A2(n16658), .ZN(N41787));
    NANDX1 U28916 (.A1(N4139), .A2(N10386), .ZN(N41788));
    INVX1 U28917 (.I(n21451), .ZN(n41789));
    NANDX1 U28918 (.A1(n19393), .A2(n23319), .ZN(n41790));
    INVX1 U28919 (.I(N6221), .ZN(n41791));
    INVX1 U28920 (.I(N2286), .ZN(N41792));
    INVX1 U28921 (.I(n16085), .ZN(N41793));
    NANDX1 U28922 (.A1(n19959), .A2(N1908), .ZN(n41794));
    INVX1 U28923 (.I(N1252), .ZN(N41795));
    NANDX1 U28924 (.A1(N4201), .A2(N319), .ZN(N41796));
    INVX1 U28925 (.I(n27609), .ZN(N41797));
    NANDX1 U28926 (.A1(N3946), .A2(N6103), .ZN(N41798));
    NOR2X1 U28927 (.A1(n15785), .A2(N534), .ZN(n41799));
    INVX1 U28928 (.I(N440), .ZN(N41800));
    NANDX1 U28929 (.A1(N5732), .A2(N11352), .ZN(n41801));
    INVX1 U28930 (.I(N4101), .ZN(N41802));
    NOR2X1 U28931 (.A1(N7864), .A2(n26751), .ZN(N41803));
    NOR2X1 U28932 (.A1(n29259), .A2(n29036), .ZN(N41804));
    NANDX1 U28933 (.A1(N3767), .A2(n24482), .ZN(N41805));
    INVX1 U28934 (.I(N5674), .ZN(N41806));
    NANDX1 U28935 (.A1(N4887), .A2(n14123), .ZN(N41807));
    INVX1 U28936 (.I(N5206), .ZN(n41808));
    NOR2X1 U28937 (.A1(N8485), .A2(n23364), .ZN(n41809));
    NANDX1 U28938 (.A1(n14587), .A2(N2053), .ZN(N41810));
    INVX1 U28939 (.I(n15120), .ZN(N41811));
    INVX1 U28940 (.I(n23916), .ZN(N41812));
    INVX1 U28941 (.I(N3131), .ZN(N41813));
    NOR2X1 U28942 (.A1(N4336), .A2(n25929), .ZN(N41814));
    NANDX1 U28943 (.A1(N760), .A2(n22542), .ZN(N41815));
    NOR2X1 U28944 (.A1(n30018), .A2(N10001), .ZN(n41816));
    INVX1 U28945 (.I(n22346), .ZN(n41817));
    NANDX1 U28946 (.A1(N7136), .A2(n16580), .ZN(N41818));
    NOR2X1 U28947 (.A1(N584), .A2(N565), .ZN(n41819));
    INVX1 U28948 (.I(n24487), .ZN(N41820));
    INVX1 U28949 (.I(N519), .ZN(n41821));
    NOR2X1 U28950 (.A1(N12002), .A2(n15106), .ZN(N41822));
    NOR2X1 U28951 (.A1(N5341), .A2(n18786), .ZN(N41823));
    NOR2X1 U28952 (.A1(n17817), .A2(n27138), .ZN(n41824));
    NOR2X1 U28953 (.A1(N11507), .A2(n20034), .ZN(n41825));
    NANDX1 U28954 (.A1(n13064), .A2(n20794), .ZN(n41826));
    NOR2X1 U28955 (.A1(N10009), .A2(N9235), .ZN(N41827));
    INVX1 U28956 (.I(n20768), .ZN(n41828));
    NANDX1 U28957 (.A1(n18656), .A2(n16464), .ZN(N41829));
    INVX1 U28958 (.I(n29814), .ZN(N41830));
    NANDX1 U28959 (.A1(N7148), .A2(N3150), .ZN(N41831));
    NANDX1 U28960 (.A1(N11459), .A2(n22366), .ZN(N41832));
    NANDX1 U28961 (.A1(n23460), .A2(N7334), .ZN(N41833));
    INVX1 U28962 (.I(n17361), .ZN(n41834));
    NOR2X1 U28963 (.A1(n24462), .A2(N5040), .ZN(N41835));
    INVX1 U28964 (.I(N3180), .ZN(N41836));
    NANDX1 U28965 (.A1(n20275), .A2(n26525), .ZN(N41837));
    INVX1 U28966 (.I(N10931), .ZN(N41838));
    NOR2X1 U28967 (.A1(n16740), .A2(n20166), .ZN(N41839));
    INVX1 U28968 (.I(n26068), .ZN(N41840));
    NANDX1 U28969 (.A1(N3528), .A2(N12394), .ZN(n41841));
    NANDX1 U28970 (.A1(N3204), .A2(n29441), .ZN(N41842));
    NANDX1 U28971 (.A1(n25051), .A2(N10699), .ZN(N41843));
    INVX1 U28972 (.I(n17280), .ZN(N41844));
    NOR2X1 U28973 (.A1(n17241), .A2(n13174), .ZN(N41845));
    INVX1 U28974 (.I(N4465), .ZN(N41846));
    NANDX1 U28975 (.A1(N11291), .A2(N9504), .ZN(n41847));
    NOR2X1 U28976 (.A1(N3032), .A2(N3172), .ZN(N41848));
    INVX1 U28977 (.I(n18117), .ZN(N41849));
    NOR2X1 U28978 (.A1(n17724), .A2(n18815), .ZN(n41850));
    NOR2X1 U28979 (.A1(n26450), .A2(N3687), .ZN(N41851));
    NOR2X1 U28980 (.A1(N6482), .A2(N7215), .ZN(n41852));
    NANDX1 U28981 (.A1(n23233), .A2(n29116), .ZN(n41853));
    NANDX1 U28982 (.A1(n16995), .A2(n24030), .ZN(n41854));
    NOR2X1 U28983 (.A1(N10776), .A2(N11172), .ZN(n41855));
    INVX1 U28984 (.I(n28017), .ZN(N41856));
    INVX1 U28985 (.I(n18588), .ZN(n41857));
    NANDX1 U28986 (.A1(n29321), .A2(n18440), .ZN(n41858));
    NOR2X1 U28987 (.A1(n15839), .A2(N10032), .ZN(N41859));
    NOR2X1 U28988 (.A1(n22632), .A2(n28148), .ZN(N41860));
    NANDX1 U28989 (.A1(N10219), .A2(n16826), .ZN(N41861));
    NOR2X1 U28990 (.A1(N6531), .A2(n20512), .ZN(N41862));
    NANDX1 U28991 (.A1(N1573), .A2(n16287), .ZN(n41863));
    NOR2X1 U28992 (.A1(n13367), .A2(n15266), .ZN(n41864));
    INVX1 U28993 (.I(n18922), .ZN(N41865));
    NANDX1 U28994 (.A1(n17850), .A2(n29698), .ZN(N41866));
    NOR2X1 U28995 (.A1(N8032), .A2(n27577), .ZN(N41867));
    NOR2X1 U28996 (.A1(n15180), .A2(n18481), .ZN(n41868));
    NOR2X1 U28997 (.A1(N3482), .A2(n18888), .ZN(N41869));
    NANDX1 U28998 (.A1(n13513), .A2(N11028), .ZN(n41870));
    NOR2X1 U28999 (.A1(N85), .A2(n24510), .ZN(N41871));
    INVX1 U29000 (.I(n16910), .ZN(n41872));
    NANDX1 U29001 (.A1(N11743), .A2(n25982), .ZN(N41873));
    INVX1 U29002 (.I(N1876), .ZN(N41874));
    NANDX1 U29003 (.A1(n24366), .A2(n15242), .ZN(N41875));
    NOR2X1 U29004 (.A1(N8687), .A2(N4027), .ZN(N41876));
    INVX1 U29005 (.I(n15097), .ZN(N41877));
    NOR2X1 U29006 (.A1(n29824), .A2(n23128), .ZN(N41878));
    NANDX1 U29007 (.A1(N10042), .A2(N8171), .ZN(n41879));
    INVX1 U29008 (.I(N8142), .ZN(N41880));
    INVX1 U29009 (.I(n15515), .ZN(N41881));
    INVX1 U29010 (.I(N2287), .ZN(N41882));
    NANDX1 U29011 (.A1(n17073), .A2(N2371), .ZN(N41883));
    NANDX1 U29012 (.A1(N3587), .A2(N7841), .ZN(n41884));
    INVX1 U29013 (.I(N3890), .ZN(N41885));
    NANDX1 U29014 (.A1(N12252), .A2(n24463), .ZN(n41886));
    NOR2X1 U29015 (.A1(n25178), .A2(N9568), .ZN(N41887));
    NANDX1 U29016 (.A1(n22426), .A2(N2155), .ZN(N41888));
    NANDX1 U29017 (.A1(n26083), .A2(n24439), .ZN(N41889));
    INVX1 U29018 (.I(N7635), .ZN(N41890));
    NOR2X1 U29019 (.A1(n28118), .A2(N4366), .ZN(N41891));
    NOR2X1 U29020 (.A1(N6122), .A2(N4578), .ZN(N41892));
    INVX1 U29021 (.I(n16762), .ZN(N41893));
    NANDX1 U29022 (.A1(n18391), .A2(N3697), .ZN(N41894));
    NANDX1 U29023 (.A1(n16427), .A2(n25981), .ZN(N41895));
    NOR2X1 U29024 (.A1(N7382), .A2(n18431), .ZN(N41896));
    NOR2X1 U29025 (.A1(N8195), .A2(N12757), .ZN(N41897));
    NANDX1 U29026 (.A1(n21933), .A2(N10885), .ZN(N41898));
    INVX1 U29027 (.I(n14221), .ZN(N41899));
    NOR2X1 U29028 (.A1(n13922), .A2(n28865), .ZN(N41900));
    NOR2X1 U29029 (.A1(N1861), .A2(N6362), .ZN(N41901));
    NOR2X1 U29030 (.A1(n29978), .A2(N10727), .ZN(N41902));
    NOR2X1 U29031 (.A1(n24660), .A2(N3865), .ZN(N41903));
    NOR2X1 U29032 (.A1(n29982), .A2(n17988), .ZN(N41904));
    INVX1 U29033 (.I(n22239), .ZN(n41905));
    NOR2X1 U29034 (.A1(N1485), .A2(n18083), .ZN(N41906));
    INVX1 U29035 (.I(n27565), .ZN(N41907));
    NOR2X1 U29036 (.A1(n22376), .A2(N5622), .ZN(N41908));
    NOR2X1 U29037 (.A1(n20452), .A2(n27554), .ZN(n41909));
    NOR2X1 U29038 (.A1(N4545), .A2(N199), .ZN(N41910));
    NANDX1 U29039 (.A1(N7028), .A2(n29063), .ZN(N41911));
    NANDX1 U29040 (.A1(N8888), .A2(n23985), .ZN(N41912));
    NANDX1 U29041 (.A1(n27426), .A2(N4574), .ZN(n41913));
    INVX1 U29042 (.I(N10509), .ZN(n41914));
    INVX1 U29043 (.I(N12142), .ZN(N41915));
    INVX1 U29044 (.I(n14986), .ZN(N41916));
    NOR2X1 U29045 (.A1(N2454), .A2(N7890), .ZN(N41917));
    INVX1 U29046 (.I(N9097), .ZN(N41918));
    NOR2X1 U29047 (.A1(n14809), .A2(N4034), .ZN(N41919));
    NANDX1 U29048 (.A1(n20430), .A2(N11726), .ZN(N41920));
    NOR2X1 U29049 (.A1(N6408), .A2(n18864), .ZN(N41921));
    NOR2X1 U29050 (.A1(N6606), .A2(n27600), .ZN(n41922));
    NOR2X1 U29051 (.A1(n24229), .A2(n20798), .ZN(N41923));
    NOR2X1 U29052 (.A1(n18076), .A2(n19739), .ZN(N41924));
    NOR2X1 U29053 (.A1(N11210), .A2(N4939), .ZN(n41925));
    INVX1 U29054 (.I(N8208), .ZN(n41926));
    NOR2X1 U29055 (.A1(n19227), .A2(N11755), .ZN(N41927));
    NANDX1 U29056 (.A1(n21680), .A2(n19644), .ZN(n41928));
    NOR2X1 U29057 (.A1(N640), .A2(n14632), .ZN(N41929));
    NOR2X1 U29058 (.A1(n23371), .A2(n20556), .ZN(n41930));
    NOR2X1 U29059 (.A1(n23657), .A2(N5355), .ZN(N41931));
    INVX1 U29060 (.I(N12383), .ZN(N41932));
    NANDX1 U29061 (.A1(N11276), .A2(n28544), .ZN(N41933));
    INVX1 U29062 (.I(N5367), .ZN(n41934));
    NANDX1 U29063 (.A1(n22285), .A2(n23442), .ZN(N41935));
    INVX1 U29064 (.I(n20651), .ZN(N41936));
    NANDX1 U29065 (.A1(N2304), .A2(N10827), .ZN(N41937));
    NOR2X1 U29066 (.A1(n26642), .A2(n18614), .ZN(N41938));
    NANDX1 U29067 (.A1(N6603), .A2(N10157), .ZN(n41939));
    NOR2X1 U29068 (.A1(N3946), .A2(n29494), .ZN(n41940));
    INVX1 U29069 (.I(N4658), .ZN(N41941));
    NANDX1 U29070 (.A1(n26290), .A2(n14360), .ZN(N41942));
    NOR2X1 U29071 (.A1(N1507), .A2(N333), .ZN(N41943));
    NANDX1 U29072 (.A1(n14904), .A2(N169), .ZN(N41944));
    NOR2X1 U29073 (.A1(n13232), .A2(N5536), .ZN(N41945));
    INVX1 U29074 (.I(n24078), .ZN(n41946));
    NOR2X1 U29075 (.A1(N9286), .A2(n14591), .ZN(N41947));
    NOR2X1 U29076 (.A1(N151), .A2(n13979), .ZN(N41948));
    NOR2X1 U29077 (.A1(n26792), .A2(N2455), .ZN(n41949));
    INVX1 U29078 (.I(N3258), .ZN(N41950));
    NANDX1 U29079 (.A1(n16034), .A2(n25901), .ZN(N41951));
    INVX1 U29080 (.I(n21768), .ZN(N41952));
    INVX1 U29081 (.I(N11815), .ZN(N41953));
    INVX1 U29082 (.I(N3341), .ZN(n41954));
    NOR2X1 U29083 (.A1(n26685), .A2(n22371), .ZN(n41955));
    NANDX1 U29084 (.A1(N11451), .A2(n22540), .ZN(N41956));
    INVX1 U29085 (.I(n24683), .ZN(N41957));
    NANDX1 U29086 (.A1(N8311), .A2(N7184), .ZN(N41958));
    NANDX1 U29087 (.A1(N6157), .A2(n21774), .ZN(N41959));
    NANDX1 U29088 (.A1(N6307), .A2(N5615), .ZN(N41960));
    INVX1 U29089 (.I(n21660), .ZN(n41961));
    NANDX1 U29090 (.A1(n21335), .A2(n13478), .ZN(N41962));
    NOR2X1 U29091 (.A1(N7231), .A2(N9241), .ZN(n41963));
    NANDX1 U29092 (.A1(n17559), .A2(n28359), .ZN(N41964));
    INVX1 U29093 (.I(n24039), .ZN(N41965));
    NOR2X1 U29094 (.A1(N3887), .A2(n20587), .ZN(N41966));
    NANDX1 U29095 (.A1(n14819), .A2(N1900), .ZN(n41967));
    NOR2X1 U29096 (.A1(N11209), .A2(n15143), .ZN(N41968));
    NANDX1 U29097 (.A1(N8080), .A2(n22326), .ZN(N41969));
    INVX1 U29098 (.I(n14237), .ZN(N41970));
    NANDX1 U29099 (.A1(N10077), .A2(N9104), .ZN(n41971));
    NOR2X1 U29100 (.A1(n17920), .A2(N626), .ZN(N41972));
    INVX1 U29101 (.I(n27816), .ZN(N41973));
    INVX1 U29102 (.I(N9829), .ZN(n41974));
    NANDX1 U29103 (.A1(N11904), .A2(n26856), .ZN(N41975));
    NANDX1 U29104 (.A1(n28823), .A2(n14121), .ZN(n41976));
    NANDX1 U29105 (.A1(n18946), .A2(n18008), .ZN(N41977));
    INVX1 U29106 (.I(N1302), .ZN(n41978));
    INVX1 U29107 (.I(n15977), .ZN(N41979));
    NANDX1 U29108 (.A1(N2459), .A2(n19680), .ZN(N41980));
    INVX1 U29109 (.I(n29236), .ZN(n41981));
    NOR2X1 U29110 (.A1(N277), .A2(N1896), .ZN(N41982));
    NANDX1 U29111 (.A1(n29051), .A2(N11000), .ZN(N41983));
    INVX1 U29112 (.I(N5395), .ZN(N41984));
    NOR2X1 U29113 (.A1(N11678), .A2(N3073), .ZN(N41985));
    INVX1 U29114 (.I(n21506), .ZN(N41986));
    NANDX1 U29115 (.A1(N3314), .A2(n18224), .ZN(n41987));
    INVX1 U29116 (.I(N2000), .ZN(N41988));
    NOR2X1 U29117 (.A1(n23939), .A2(n20945), .ZN(n41989));
    NANDX1 U29118 (.A1(N7878), .A2(n22246), .ZN(N41990));
    INVX1 U29119 (.I(N12415), .ZN(N41991));
    NANDX1 U29120 (.A1(N2483), .A2(N1958), .ZN(N41992));
    NANDX1 U29121 (.A1(N1581), .A2(N2387), .ZN(N41993));
    NOR2X1 U29122 (.A1(N3477), .A2(N5339), .ZN(N41994));
    NANDX1 U29123 (.A1(N3037), .A2(n23687), .ZN(N41995));
    NANDX1 U29124 (.A1(N3222), .A2(N5227), .ZN(N41996));
    NANDX1 U29125 (.A1(n24769), .A2(n26732), .ZN(n41997));
    INVX1 U29126 (.I(n28083), .ZN(N41998));
    INVX1 U29127 (.I(N10740), .ZN(n41999));
    NANDX1 U29128 (.A1(n24284), .A2(n23239), .ZN(N42000));
    NOR2X1 U29129 (.A1(N2921), .A2(N979), .ZN(N42001));
    NOR2X1 U29130 (.A1(N2945), .A2(n13394), .ZN(N42002));
    INVX1 U29131 (.I(n24125), .ZN(N42003));
    NOR2X1 U29132 (.A1(n17532), .A2(n14267), .ZN(N42004));
    NANDX1 U29133 (.A1(n16780), .A2(n17743), .ZN(N42005));
    NOR2X1 U29134 (.A1(N3503), .A2(N9340), .ZN(N42006));
    INVX1 U29135 (.I(N7059), .ZN(n42007));
    NOR2X1 U29136 (.A1(n29110), .A2(N2248), .ZN(N42008));
    NOR2X1 U29137 (.A1(n14265), .A2(N5418), .ZN(n42009));
    NOR2X1 U29138 (.A1(n17644), .A2(N4718), .ZN(n42010));
    INVX1 U29139 (.I(N11790), .ZN(N42011));
    NOR2X1 U29140 (.A1(n14531), .A2(N3271), .ZN(N42012));
    NOR2X1 U29141 (.A1(n16088), .A2(n24914), .ZN(N42013));
    NOR2X1 U29142 (.A1(n23208), .A2(N7462), .ZN(N42014));
    NANDX1 U29143 (.A1(n29300), .A2(n21728), .ZN(N42015));
    NOR2X1 U29144 (.A1(N4503), .A2(n28031), .ZN(N42016));
    NANDX1 U29145 (.A1(N8006), .A2(N7233), .ZN(n42017));
    INVX1 U29146 (.I(n15064), .ZN(N42018));
    NOR2X1 U29147 (.A1(N11132), .A2(N5873), .ZN(N42019));
    NANDX1 U29148 (.A1(n13957), .A2(N11290), .ZN(N42020));
    INVX1 U29149 (.I(N1463), .ZN(n42021));
    NOR2X1 U29150 (.A1(N10146), .A2(N1813), .ZN(N42022));
    NOR2X1 U29151 (.A1(n24676), .A2(n23782), .ZN(n42023));
    NANDX1 U29152 (.A1(n29324), .A2(N7119), .ZN(N42024));
    NANDX1 U29153 (.A1(N10955), .A2(n14580), .ZN(N42025));
    NOR2X1 U29154 (.A1(n28815), .A2(N6171), .ZN(N42026));
    INVX1 U29155 (.I(N3180), .ZN(n42027));
    INVX1 U29156 (.I(N8908), .ZN(N42028));
    NANDX1 U29157 (.A1(n29995), .A2(n21067), .ZN(N42029));
    NANDX1 U29158 (.A1(n26910), .A2(N2061), .ZN(N42030));
    INVX1 U29159 (.I(n19578), .ZN(N42031));
    INVX1 U29160 (.I(n20532), .ZN(n42032));
    NANDX1 U29161 (.A1(N6041), .A2(n25099), .ZN(N42033));
    NOR2X1 U29162 (.A1(n26552), .A2(n27484), .ZN(n42034));
    INVX1 U29163 (.I(N8757), .ZN(N42035));
    NANDX1 U29164 (.A1(n28511), .A2(n15875), .ZN(n42036));
    NOR2X1 U29165 (.A1(N9328), .A2(n19015), .ZN(n42037));
    INVX1 U29166 (.I(N8005), .ZN(n42038));
    NANDX1 U29167 (.A1(n26584), .A2(n29882), .ZN(N42039));
    NOR2X1 U29168 (.A1(N5354), .A2(N10930), .ZN(N42040));
    NOR2X1 U29169 (.A1(n14982), .A2(n14300), .ZN(N42041));
    NANDX1 U29170 (.A1(n17042), .A2(n23542), .ZN(n42042));
    INVX1 U29171 (.I(n21620), .ZN(n42043));
    NANDX1 U29172 (.A1(n17081), .A2(n16222), .ZN(n42044));
    NANDX1 U29173 (.A1(N3032), .A2(N1197), .ZN(N42045));
    NANDX1 U29174 (.A1(N2219), .A2(n28651), .ZN(n42046));
    NOR2X1 U29175 (.A1(N592), .A2(N2949), .ZN(N42047));
    INVX1 U29176 (.I(n28617), .ZN(n42048));
    NOR2X1 U29177 (.A1(n28779), .A2(n25182), .ZN(n42049));
    NANDX1 U29178 (.A1(n13786), .A2(n24926), .ZN(n42050));
    NANDX1 U29179 (.A1(N7700), .A2(n24416), .ZN(N42051));
    INVX1 U29180 (.I(n22681), .ZN(n42052));
    INVX1 U29181 (.I(N5549), .ZN(n42053));
    INVX1 U29182 (.I(N1982), .ZN(N42054));
    NOR2X1 U29183 (.A1(N8327), .A2(N4478), .ZN(N42055));
    NANDX1 U29184 (.A1(n13109), .A2(n20633), .ZN(N42056));
    INVX1 U29185 (.I(N2866), .ZN(n42057));
    NOR2X1 U29186 (.A1(n23396), .A2(N1379), .ZN(n42058));
    INVX1 U29187 (.I(n23987), .ZN(N42059));
    INVX1 U29188 (.I(n23233), .ZN(n42060));
    NANDX1 U29189 (.A1(n14851), .A2(N10435), .ZN(N42061));
    INVX1 U29190 (.I(N8983), .ZN(N42062));
    NOR2X1 U29191 (.A1(N859), .A2(N9485), .ZN(n42063));
    NANDX1 U29192 (.A1(n25275), .A2(n23473), .ZN(N42064));
    INVX1 U29193 (.I(n22413), .ZN(n42065));
    NANDX1 U29194 (.A1(N11170), .A2(n24395), .ZN(N42066));
    NANDX1 U29195 (.A1(n19496), .A2(n17433), .ZN(n42067));
    INVX1 U29196 (.I(N2468), .ZN(N42068));
    NOR2X1 U29197 (.A1(n13316), .A2(N5333), .ZN(N42069));
    NANDX1 U29198 (.A1(N6574), .A2(n25410), .ZN(N42070));
    NANDX1 U29199 (.A1(N423), .A2(n29736), .ZN(N42071));
    NOR2X1 U29200 (.A1(N11449), .A2(N3010), .ZN(N42072));
    NANDX1 U29201 (.A1(N6080), .A2(N11992), .ZN(n42073));
    INVX1 U29202 (.I(n25636), .ZN(N42074));
    INVX1 U29203 (.I(n14803), .ZN(n42075));
    NOR2X1 U29204 (.A1(N3372), .A2(n16387), .ZN(N42076));
    NANDX1 U29205 (.A1(n20953), .A2(n27556), .ZN(n42077));
    INVX1 U29206 (.I(N2204), .ZN(N42078));
    NOR2X1 U29207 (.A1(N1860), .A2(n24479), .ZN(n42079));
    INVX1 U29208 (.I(n17047), .ZN(N42080));
    NANDX1 U29209 (.A1(N1836), .A2(n24792), .ZN(n42081));
    INVX1 U29210 (.I(n27245), .ZN(N42082));
    NOR2X1 U29211 (.A1(N3213), .A2(n15404), .ZN(n42083));
    NOR2X1 U29212 (.A1(N3222), .A2(n18414), .ZN(N42084));
    INVX1 U29213 (.I(n27999), .ZN(N42085));
    NANDX1 U29214 (.A1(n17312), .A2(n23498), .ZN(N42086));
    NOR2X1 U29215 (.A1(n20675), .A2(N2694), .ZN(N42087));
    NANDX1 U29216 (.A1(N6924), .A2(N4303), .ZN(N42088));
    INVX1 U29217 (.I(n23040), .ZN(N42089));
    NANDX1 U29218 (.A1(n25393), .A2(n28514), .ZN(n42090));
    INVX1 U29219 (.I(N8296), .ZN(N42091));
    INVX1 U29220 (.I(n26334), .ZN(N42092));
    NANDX1 U29221 (.A1(n26852), .A2(n20988), .ZN(n42093));
    NOR2X1 U29222 (.A1(n23959), .A2(n23793), .ZN(N42094));
    INVX1 U29223 (.I(N9225), .ZN(N42095));
    INVX1 U29224 (.I(n20997), .ZN(N42096));
    NOR2X1 U29225 (.A1(n20694), .A2(n18858), .ZN(N42097));
    NANDX1 U29226 (.A1(n26566), .A2(N12218), .ZN(n42098));
    INVX1 U29227 (.I(n17103), .ZN(n42099));
    NANDX1 U29228 (.A1(n24827), .A2(N12587), .ZN(N42100));
    NOR2X1 U29229 (.A1(n17879), .A2(N5489), .ZN(N42101));
    NOR2X1 U29230 (.A1(N1696), .A2(N3866), .ZN(n42102));
    NOR2X1 U29231 (.A1(n28689), .A2(n28882), .ZN(N42103));
    NOR2X1 U29232 (.A1(N3064), .A2(n14157), .ZN(N42104));
    NANDX1 U29233 (.A1(N10367), .A2(N7978), .ZN(N42105));
    NANDX1 U29234 (.A1(N9444), .A2(N5763), .ZN(N42106));
    NANDX1 U29235 (.A1(n19001), .A2(N10523), .ZN(N42107));
    NOR2X1 U29236 (.A1(N7721), .A2(N4111), .ZN(N42108));
    NANDX1 U29237 (.A1(N8500), .A2(N8003), .ZN(N42109));
    INVX1 U29238 (.I(n23411), .ZN(N42110));
    NOR2X1 U29239 (.A1(N3952), .A2(N1048), .ZN(n42111));
    INVX1 U29240 (.I(n28138), .ZN(n42112));
    INVX1 U29241 (.I(n29525), .ZN(N42113));
    INVX1 U29242 (.I(n22041), .ZN(N42114));
    NOR2X1 U29243 (.A1(n19308), .A2(n24029), .ZN(N42115));
    NOR2X1 U29244 (.A1(N3327), .A2(N5428), .ZN(N42116));
    NANDX1 U29245 (.A1(n30002), .A2(n29317), .ZN(n42117));
    NANDX1 U29246 (.A1(n24326), .A2(N9335), .ZN(N42118));
    NOR2X1 U29247 (.A1(N4711), .A2(n28744), .ZN(n42119));
    NANDX1 U29248 (.A1(N8821), .A2(n14445), .ZN(n42120));
    NANDX1 U29249 (.A1(N5384), .A2(N5810), .ZN(n42121));
    INVX1 U29250 (.I(n26773), .ZN(n42122));
    INVX1 U29251 (.I(N4596), .ZN(n42123));
    NANDX1 U29252 (.A1(N7761), .A2(n20845), .ZN(n42124));
    NOR2X1 U29253 (.A1(n28325), .A2(N12749), .ZN(N42125));
    NOR2X1 U29254 (.A1(N6056), .A2(n25338), .ZN(n42126));
    INVX1 U29255 (.I(N9383), .ZN(N42127));
    NANDX1 U29256 (.A1(n25800), .A2(n27945), .ZN(N42128));
    NANDX1 U29257 (.A1(n23733), .A2(n22133), .ZN(N42129));
    NANDX1 U29258 (.A1(n29227), .A2(n15404), .ZN(n42130));
    INVX1 U29259 (.I(N865), .ZN(N42131));
    NANDX1 U29260 (.A1(n29451), .A2(n22579), .ZN(N42132));
    NOR2X1 U29261 (.A1(N5123), .A2(n26126), .ZN(N42133));
    NANDX1 U29262 (.A1(N3444), .A2(n19282), .ZN(n42134));
    NOR2X1 U29263 (.A1(N11204), .A2(n28688), .ZN(n42135));
    INVX1 U29264 (.I(N9391), .ZN(N42136));
    NANDX1 U29265 (.A1(N4836), .A2(n15447), .ZN(n42137));
    NANDX1 U29266 (.A1(N12008), .A2(n13390), .ZN(N42138));
    NOR2X1 U29267 (.A1(N7670), .A2(n29895), .ZN(n42139));
    NANDX1 U29268 (.A1(n19963), .A2(N10452), .ZN(N42140));
    INVX1 U29269 (.I(N7613), .ZN(N42141));
    NOR2X1 U29270 (.A1(N11278), .A2(N8478), .ZN(N42142));
    NANDX1 U29271 (.A1(n29289), .A2(N919), .ZN(n42143));
    NANDX1 U29272 (.A1(n22972), .A2(n15605), .ZN(N42144));
    INVX1 U29273 (.I(n26415), .ZN(N42145));
    INVX1 U29274 (.I(N12107), .ZN(N42146));
    NANDX1 U29275 (.A1(N3300), .A2(n18031), .ZN(n42147));
    NANDX1 U29276 (.A1(N3159), .A2(n22866), .ZN(n42148));
    NANDX1 U29277 (.A1(n16916), .A2(n23435), .ZN(N42149));
    NOR2X1 U29278 (.A1(n19861), .A2(N967), .ZN(N42150));
    INVX1 U29279 (.I(n29871), .ZN(N42151));
    NOR2X1 U29280 (.A1(n21599), .A2(n26143), .ZN(N42152));
    INVX1 U29281 (.I(n17316), .ZN(N42153));
    NANDX1 U29282 (.A1(n14141), .A2(n14379), .ZN(N42154));
    NANDX1 U29283 (.A1(N3620), .A2(n18171), .ZN(n42155));
    NANDX1 U29284 (.A1(n19225), .A2(n13887), .ZN(N42156));
    INVX1 U29285 (.I(N12535), .ZN(n42157));
    INVX1 U29286 (.I(N10287), .ZN(N42158));
    INVX1 U29287 (.I(N2447), .ZN(n42159));
    INVX1 U29288 (.I(N7553), .ZN(N42160));
    INVX1 U29289 (.I(n25159), .ZN(n42161));
    NANDX1 U29290 (.A1(N7171), .A2(N6411), .ZN(N42162));
    NOR2X1 U29291 (.A1(n26835), .A2(n17558), .ZN(n42163));
    NOR2X1 U29292 (.A1(N6188), .A2(N9019), .ZN(N42164));
    INVX1 U29293 (.I(N11852), .ZN(n42165));
    INVX1 U29294 (.I(n13031), .ZN(n42166));
    NANDX1 U29295 (.A1(n17835), .A2(n26724), .ZN(n42167));
    NANDX1 U29296 (.A1(n24566), .A2(N3115), .ZN(N42168));
    INVX1 U29297 (.I(N8316), .ZN(N42169));
    NANDX1 U29298 (.A1(N8355), .A2(n22869), .ZN(N42170));
    INVX1 U29299 (.I(N12749), .ZN(n42171));
    INVX1 U29300 (.I(n20485), .ZN(n42172));
    NOR2X1 U29301 (.A1(N9052), .A2(n15506), .ZN(n42173));
    INVX1 U29302 (.I(n16222), .ZN(N42174));
    NANDX1 U29303 (.A1(n13202), .A2(N1480), .ZN(N42175));
    INVX1 U29304 (.I(N4247), .ZN(N42176));
    NANDX1 U29305 (.A1(n25615), .A2(n21434), .ZN(N42177));
    INVX1 U29306 (.I(n29071), .ZN(N42178));
    NOR2X1 U29307 (.A1(n22632), .A2(N5329), .ZN(n42179));
    NANDX1 U29308 (.A1(n29365), .A2(n18456), .ZN(N42180));
    NANDX1 U29309 (.A1(n25185), .A2(n15332), .ZN(N42181));
    NOR2X1 U29310 (.A1(N3402), .A2(N8063), .ZN(N42182));
    INVX1 U29311 (.I(N4711), .ZN(n42183));
    NANDX1 U29312 (.A1(N12319), .A2(n13572), .ZN(n42184));
    INVX1 U29313 (.I(n16386), .ZN(N42185));
    NOR2X1 U29314 (.A1(n24333), .A2(n26863), .ZN(N42186));
    INVX1 U29315 (.I(n25813), .ZN(N42187));
    NOR2X1 U29316 (.A1(n30030), .A2(n22041), .ZN(N42188));
    NANDX1 U29317 (.A1(N9887), .A2(n30120), .ZN(N42189));
    INVX1 U29318 (.I(N2775), .ZN(n42190));
    NANDX1 U29319 (.A1(n20319), .A2(N10947), .ZN(N42191));
    NOR2X1 U29320 (.A1(N8637), .A2(N10794), .ZN(N42192));
    NOR2X1 U29321 (.A1(N12529), .A2(n27999), .ZN(n42193));
    INVX1 U29322 (.I(N9152), .ZN(N42194));
    NANDX1 U29323 (.A1(N2123), .A2(N954), .ZN(N42195));
    NOR2X1 U29324 (.A1(N4256), .A2(N9065), .ZN(n42196));
    NOR2X1 U29325 (.A1(n28277), .A2(N3261), .ZN(N42197));
    INVX1 U29326 (.I(n23924), .ZN(N42198));
    INVX1 U29327 (.I(N5567), .ZN(N42199));
    INVX1 U29328 (.I(n28235), .ZN(N42200));
    NOR2X1 U29329 (.A1(n22264), .A2(n28217), .ZN(N42201));
    NANDX1 U29330 (.A1(n13599), .A2(n27952), .ZN(n42202));
    NOR2X1 U29331 (.A1(n13106), .A2(n26915), .ZN(N42203));
    INVX1 U29332 (.I(n23899), .ZN(N42204));
    NANDX1 U29333 (.A1(n17821), .A2(N10321), .ZN(n42205));
    NANDX1 U29334 (.A1(n26972), .A2(n18714), .ZN(N42206));
    NANDX1 U29335 (.A1(n16486), .A2(N9288), .ZN(N42207));
    INVX1 U29336 (.I(n14112), .ZN(N42208));
    NANDX1 U29337 (.A1(n22855), .A2(N5933), .ZN(N42209));
    NOR2X1 U29338 (.A1(N5202), .A2(n23566), .ZN(N42210));
    INVX1 U29339 (.I(N6139), .ZN(N42211));
    NANDX1 U29340 (.A1(N5545), .A2(n16963), .ZN(N42212));
    NANDX1 U29341 (.A1(N12020), .A2(N424), .ZN(N42213));
    INVX1 U29342 (.I(N8676), .ZN(N42214));
    NOR2X1 U29343 (.A1(n21593), .A2(n13968), .ZN(n42215));
    NANDX1 U29344 (.A1(n23820), .A2(n20349), .ZN(n42216));
    NOR2X1 U29345 (.A1(N12020), .A2(N5744), .ZN(N42217));
    INVX1 U29346 (.I(N2342), .ZN(N42218));
    INVX1 U29347 (.I(n22733), .ZN(N42219));
    NOR2X1 U29348 (.A1(n24902), .A2(n16102), .ZN(N42220));
    NOR2X1 U29349 (.A1(N697), .A2(n13155), .ZN(N42221));
    NOR2X1 U29350 (.A1(N12823), .A2(N4336), .ZN(N42222));
    NOR2X1 U29351 (.A1(n23046), .A2(n28578), .ZN(n42223));
    INVX1 U29352 (.I(N1211), .ZN(N42224));
    NOR2X1 U29353 (.A1(n14182), .A2(n14586), .ZN(N42225));
    NANDX1 U29354 (.A1(n16272), .A2(N6041), .ZN(n42226));
    NANDX1 U29355 (.A1(N12122), .A2(n18421), .ZN(N42227));
    NANDX1 U29356 (.A1(n18293), .A2(n19001), .ZN(n42228));
    INVX1 U29357 (.I(N1600), .ZN(N42229));
    NANDX1 U29358 (.A1(N5529), .A2(n24332), .ZN(N42230));
    INVX1 U29359 (.I(N293), .ZN(n42231));
    NOR2X1 U29360 (.A1(n22416), .A2(n19687), .ZN(N42232));
    NANDX1 U29361 (.A1(n13073), .A2(N2372), .ZN(N42233));
    INVX1 U29362 (.I(N9868), .ZN(N42234));
    INVX1 U29363 (.I(n14787), .ZN(N42235));
    NANDX1 U29364 (.A1(n15188), .A2(n13807), .ZN(n42236));
    INVX1 U29365 (.I(n18335), .ZN(N42237));
    NOR2X1 U29366 (.A1(N1064), .A2(n24375), .ZN(N42238));
    INVX1 U29367 (.I(n13185), .ZN(n42239));
    NOR2X1 U29368 (.A1(N2022), .A2(N1340), .ZN(N42240));
    NANDX1 U29369 (.A1(n26897), .A2(N2940), .ZN(N42241));
    NOR2X1 U29370 (.A1(N2289), .A2(n15832), .ZN(N42242));
    NOR2X1 U29371 (.A1(n21279), .A2(n14689), .ZN(N42243));
    NANDX1 U29372 (.A1(N10829), .A2(n26700), .ZN(n42244));
    INVX1 U29373 (.I(N1761), .ZN(N42245));
    NANDX1 U29374 (.A1(n29285), .A2(n15739), .ZN(N42246));
    NOR2X1 U29375 (.A1(n30032), .A2(n19487), .ZN(N42247));
    NOR2X1 U29376 (.A1(n26263), .A2(N7684), .ZN(N42248));
    NANDX1 U29377 (.A1(n15887), .A2(N1922), .ZN(N42249));
    NOR2X1 U29378 (.A1(n29072), .A2(n21839), .ZN(N42250));
    NANDX1 U29379 (.A1(n18972), .A2(N11921), .ZN(n42251));
    NANDX1 U29380 (.A1(N10472), .A2(N11907), .ZN(N42252));
    INVX1 U29381 (.I(n14865), .ZN(n42253));
    NOR2X1 U29382 (.A1(N3784), .A2(n29553), .ZN(N42254));
    NOR2X1 U29383 (.A1(N3173), .A2(n26115), .ZN(N42255));
    NOR2X1 U29384 (.A1(N4933), .A2(n16145), .ZN(N42256));
    NANDX1 U29385 (.A1(n20671), .A2(n20961), .ZN(N42257));
    NOR2X1 U29386 (.A1(N10021), .A2(n28144), .ZN(N42258));
    INVX1 U29387 (.I(n17704), .ZN(N42259));
    NOR2X1 U29388 (.A1(N9773), .A2(N8186), .ZN(N42260));
    NANDX1 U29389 (.A1(n27405), .A2(n30024), .ZN(n42261));
    INVX1 U29390 (.I(n16239), .ZN(N42262));
    NOR2X1 U29391 (.A1(N9196), .A2(n15272), .ZN(N42263));
    NANDX1 U29392 (.A1(N10399), .A2(n30136), .ZN(N42264));
    NANDX1 U29393 (.A1(n14182), .A2(n29551), .ZN(N42265));
    INVX1 U29394 (.I(N5915), .ZN(n42266));
    NANDX1 U29395 (.A1(n20448), .A2(N10847), .ZN(N42267));
    NOR2X1 U29396 (.A1(n29752), .A2(n20079), .ZN(n42268));
    INVX1 U29397 (.I(N8814), .ZN(N42269));
    INVX1 U29398 (.I(n26321), .ZN(N42270));
    NANDX1 U29399 (.A1(n24924), .A2(n22874), .ZN(N42271));
    INVX1 U29400 (.I(n21671), .ZN(N42272));
    NOR2X1 U29401 (.A1(N9739), .A2(n21557), .ZN(N42273));
    INVX1 U29402 (.I(n14538), .ZN(n42274));
    NOR2X1 U29403 (.A1(n27598), .A2(n29809), .ZN(n42275));
    NANDX1 U29404 (.A1(N7859), .A2(n18368), .ZN(N42276));
    INVX1 U29405 (.I(N10601), .ZN(n42277));
    NANDX1 U29406 (.A1(N6842), .A2(n16515), .ZN(n42278));
    INVX1 U29407 (.I(n27289), .ZN(N42279));
    NOR2X1 U29408 (.A1(N9086), .A2(n15465), .ZN(N42280));
    NOR2X1 U29409 (.A1(N7263), .A2(n24278), .ZN(N42281));
    INVX1 U29410 (.I(N3446), .ZN(n42282));
    NOR2X1 U29411 (.A1(N7870), .A2(n26319), .ZN(N42283));
    INVX1 U29412 (.I(n29540), .ZN(N42284));
    NOR2X1 U29413 (.A1(n26308), .A2(N9521), .ZN(n42285));
    NOR2X1 U29414 (.A1(n29407), .A2(n20006), .ZN(N42286));
    NOR2X1 U29415 (.A1(n17639), .A2(N1190), .ZN(N42287));
    INVX1 U29416 (.I(N5870), .ZN(N42288));
    NOR2X1 U29417 (.A1(n27186), .A2(N12211), .ZN(n42289));
    INVX1 U29418 (.I(N2124), .ZN(N42290));
    INVX1 U29419 (.I(n20433), .ZN(n42291));
    NANDX1 U29420 (.A1(N150), .A2(N5760), .ZN(N42292));
    NANDX1 U29421 (.A1(N7413), .A2(n18598), .ZN(n42293));
    NANDX1 U29422 (.A1(N10858), .A2(N3999), .ZN(N42294));
    NANDX1 U29423 (.A1(n25738), .A2(n20568), .ZN(N42295));
    NOR2X1 U29424 (.A1(n18601), .A2(N5300), .ZN(N42296));
    INVX1 U29425 (.I(N11169), .ZN(N42297));
    INVX1 U29426 (.I(N9336), .ZN(n42298));
    NOR2X1 U29427 (.A1(N10768), .A2(n29223), .ZN(N42299));
    INVX1 U29428 (.I(N5198), .ZN(N42300));
    NOR2X1 U29429 (.A1(n22088), .A2(N5970), .ZN(N42301));
    NOR2X1 U29430 (.A1(n24212), .A2(n27171), .ZN(N42302));
    NANDX1 U29431 (.A1(N681), .A2(n27320), .ZN(N42303));
    NANDX1 U29432 (.A1(n13151), .A2(n23293), .ZN(N42304));
    NOR2X1 U29433 (.A1(n27264), .A2(n22712), .ZN(N42305));
    NOR2X1 U29434 (.A1(n19110), .A2(N6873), .ZN(N42306));
    INVX1 U29435 (.I(N10359), .ZN(n42307));
    INVX1 U29436 (.I(N11608), .ZN(N42308));
    INVX1 U29437 (.I(n25202), .ZN(n42309));
    INVX1 U29438 (.I(N9023), .ZN(N42310));
    INVX1 U29439 (.I(n15505), .ZN(N42311));
    NANDX1 U29440 (.A1(n28560), .A2(N9263), .ZN(n42312));
    INVX1 U29441 (.I(N9071), .ZN(N42313));
    NOR2X1 U29442 (.A1(n25041), .A2(n21843), .ZN(n42314));
    NANDX1 U29443 (.A1(n16744), .A2(n22524), .ZN(N42315));
    NANDX1 U29444 (.A1(N2768), .A2(n24235), .ZN(n42316));
    NOR2X1 U29445 (.A1(n26087), .A2(n21361), .ZN(N42317));
    NANDX1 U29446 (.A1(n23267), .A2(N10334), .ZN(N42318));
    NOR2X1 U29447 (.A1(N10877), .A2(N9253), .ZN(n42319));
    INVX1 U29448 (.I(n22485), .ZN(N42320));
    NOR2X1 U29449 (.A1(N6967), .A2(n15782), .ZN(n42321));
    INVX1 U29450 (.I(N10487), .ZN(N42322));
    NOR2X1 U29451 (.A1(n14631), .A2(n27607), .ZN(N42323));
    NOR2X1 U29452 (.A1(N8126), .A2(N6540), .ZN(n42324));
    NOR2X1 U29453 (.A1(N3029), .A2(n16944), .ZN(n42325));
    NANDX1 U29454 (.A1(n19772), .A2(N9330), .ZN(N42326));
    NOR2X1 U29455 (.A1(N11100), .A2(n22125), .ZN(N42327));
    NOR2X1 U29456 (.A1(n25747), .A2(N1909), .ZN(N42328));
    NANDX1 U29457 (.A1(n18876), .A2(N12242), .ZN(n42329));
    NANDX1 U29458 (.A1(n18314), .A2(N10055), .ZN(N42330));
    NANDX1 U29459 (.A1(n29359), .A2(n18995), .ZN(N42331));
    NANDX1 U29460 (.A1(n15003), .A2(n25518), .ZN(N42332));
    NANDX1 U29461 (.A1(N4713), .A2(n28709), .ZN(n42333));
    NOR2X1 U29462 (.A1(N3685), .A2(N6697), .ZN(n42334));
    INVX1 U29463 (.I(n25147), .ZN(n42335));
    NANDX1 U29464 (.A1(n23573), .A2(n28737), .ZN(N42336));
    INVX1 U29465 (.I(n21463), .ZN(N42337));
    INVX1 U29466 (.I(n17718), .ZN(n42338));
    NANDX1 U29467 (.A1(n26176), .A2(n13328), .ZN(n42339));
    NANDX1 U29468 (.A1(n24452), .A2(N2066), .ZN(n42340));
    INVX1 U29469 (.I(n20596), .ZN(n42341));
    NANDX1 U29470 (.A1(n14777), .A2(n28643), .ZN(N42342));
    INVX1 U29471 (.I(N3634), .ZN(N42343));
    NOR2X1 U29472 (.A1(n23164), .A2(n17712), .ZN(N42344));
    INVX1 U29473 (.I(n16437), .ZN(N42345));
    NANDX1 U29474 (.A1(n27669), .A2(N8682), .ZN(n42346));
    NOR2X1 U29475 (.A1(n22859), .A2(N3691), .ZN(n42347));
    NANDX1 U29476 (.A1(N4856), .A2(N2291), .ZN(n42348));
    NOR2X1 U29477 (.A1(n26318), .A2(n28445), .ZN(n42349));
    INVX1 U29478 (.I(n28329), .ZN(N42350));
    INVX1 U29479 (.I(N5913), .ZN(N42351));
    NOR2X1 U29480 (.A1(N7358), .A2(n26676), .ZN(N42352));
    NOR2X1 U29481 (.A1(n16515), .A2(N5479), .ZN(N42353));
    NOR2X1 U29482 (.A1(N3581), .A2(n13639), .ZN(N42354));
    NANDX1 U29483 (.A1(N5660), .A2(n25363), .ZN(N42355));
    NOR2X1 U29484 (.A1(n21799), .A2(N223), .ZN(N42356));
    NANDX1 U29485 (.A1(N7891), .A2(N8904), .ZN(N42357));
    NANDX1 U29486 (.A1(N612), .A2(N12595), .ZN(n42358));
    NOR2X1 U29487 (.A1(n24165), .A2(N3446), .ZN(n42359));
    INVX1 U29488 (.I(n20346), .ZN(N42360));
    NOR2X1 U29489 (.A1(n25175), .A2(N7098), .ZN(n42361));
    INVX1 U29490 (.I(N950), .ZN(N42362));
    NANDX1 U29491 (.A1(n29413), .A2(n27625), .ZN(N42363));
    NANDX1 U29492 (.A1(n15790), .A2(n21664), .ZN(N42364));
    NOR2X1 U29493 (.A1(n19370), .A2(N5166), .ZN(N42365));
    NANDX1 U29494 (.A1(n13590), .A2(n19089), .ZN(n42366));
    NANDX1 U29495 (.A1(N5251), .A2(N7873), .ZN(N42367));
    INVX1 U29496 (.I(n13141), .ZN(N42368));
    NOR2X1 U29497 (.A1(n23787), .A2(N2314), .ZN(N42369));
    INVX1 U29498 (.I(n28493), .ZN(N42370));
    NANDX1 U29499 (.A1(N9937), .A2(n19506), .ZN(n42371));
    INVX1 U29500 (.I(N251), .ZN(n42372));
    NOR2X1 U29501 (.A1(N905), .A2(N3608), .ZN(n42373));
    INVX1 U29502 (.I(N10112), .ZN(n42374));
    NANDX1 U29503 (.A1(n20239), .A2(n26151), .ZN(n42375));
    INVX1 U29504 (.I(N11765), .ZN(N42376));
    NOR2X1 U29505 (.A1(n15164), .A2(N5491), .ZN(n42377));
    NANDX1 U29506 (.A1(n28754), .A2(n13141), .ZN(N42378));
    NOR2X1 U29507 (.A1(n22565), .A2(n21013), .ZN(n42379));
    INVX1 U29508 (.I(n24267), .ZN(n42380));
    NANDX1 U29509 (.A1(N5619), .A2(n26580), .ZN(N42381));
    NOR2X1 U29510 (.A1(n22673), .A2(N11481), .ZN(N42382));
    INVX1 U29511 (.I(N602), .ZN(n42383));
    NANDX1 U29512 (.A1(n12890), .A2(n22404), .ZN(N42384));
    NANDX1 U29513 (.A1(N5058), .A2(n15017), .ZN(N42385));
    NANDX1 U29514 (.A1(n26639), .A2(n23816), .ZN(N42386));
    NANDX1 U29515 (.A1(n22433), .A2(n24142), .ZN(n42387));
    NANDX1 U29516 (.A1(n26157), .A2(n18193), .ZN(N42388));
    NOR2X1 U29517 (.A1(n13334), .A2(N1196), .ZN(N42389));
    INVX1 U29518 (.I(N5762), .ZN(N42390));
    NOR2X1 U29519 (.A1(N12828), .A2(n30028), .ZN(n42391));
    NOR2X1 U29520 (.A1(N7008), .A2(n15031), .ZN(N42392));
    NOR2X1 U29521 (.A1(n18241), .A2(n15072), .ZN(N42393));
    NOR2X1 U29522 (.A1(n18842), .A2(N8921), .ZN(n42394));
    INVX1 U29523 (.I(n29806), .ZN(N42395));
    INVX1 U29524 (.I(n17392), .ZN(n42396));
    INVX1 U29525 (.I(n19979), .ZN(N42397));
    INVX1 U29526 (.I(n27062), .ZN(N42398));
    INVX1 U29527 (.I(n13447), .ZN(N42399));
    NOR2X1 U29528 (.A1(n21077), .A2(n28165), .ZN(N42400));
    NOR2X1 U29529 (.A1(n15992), .A2(N11361), .ZN(n42401));
    INVX1 U29530 (.I(n16850), .ZN(n42402));
    NOR2X1 U29531 (.A1(n28345), .A2(n29678), .ZN(n42403));
    NANDX1 U29532 (.A1(n23886), .A2(n25246), .ZN(N42404));
    INVX1 U29533 (.I(n22130), .ZN(n42405));
    INVX1 U29534 (.I(n24236), .ZN(N42406));
    NOR2X1 U29535 (.A1(n20751), .A2(N3019), .ZN(N42407));
    INVX1 U29536 (.I(n20420), .ZN(n42408));
    NOR2X1 U29537 (.A1(n21163), .A2(n23666), .ZN(n42409));
    NANDX1 U29538 (.A1(N12177), .A2(N9151), .ZN(N42410));
    NOR2X1 U29539 (.A1(n25624), .A2(N80), .ZN(N42411));
    NANDX1 U29540 (.A1(n23651), .A2(n27899), .ZN(N42412));
    NANDX1 U29541 (.A1(n23572), .A2(n15337), .ZN(N42413));
    NANDX1 U29542 (.A1(n29255), .A2(N2105), .ZN(N42414));
    NANDX1 U29543 (.A1(N4690), .A2(n14551), .ZN(N42415));
    INVX1 U29544 (.I(n13854), .ZN(n42416));
    NOR2X1 U29545 (.A1(n22108), .A2(N7952), .ZN(N42417));
    NOR2X1 U29546 (.A1(N12722), .A2(N10970), .ZN(N42418));
    NOR2X1 U29547 (.A1(n21702), .A2(n17663), .ZN(n42419));
    INVX1 U29548 (.I(N3791), .ZN(N42420));
    INVX1 U29549 (.I(N12211), .ZN(N42421));
    NANDX1 U29550 (.A1(n27406), .A2(n26395), .ZN(N42422));
    INVX1 U29551 (.I(N12856), .ZN(N42423));
    NANDX1 U29552 (.A1(n18040), .A2(N2859), .ZN(n42424));
    NANDX1 U29553 (.A1(N3240), .A2(N9712), .ZN(n42425));
    NOR2X1 U29554 (.A1(n24042), .A2(N4665), .ZN(N42426));
    INVX1 U29555 (.I(N8456), .ZN(N42427));
    INVX1 U29556 (.I(N8124), .ZN(N42428));
    INVX1 U29557 (.I(N5395), .ZN(n42429));
    INVX1 U29558 (.I(n20236), .ZN(N42430));
    NANDX1 U29559 (.A1(n27044), .A2(n29245), .ZN(N42431));
    NANDX1 U29560 (.A1(n14569), .A2(n29278), .ZN(N42432));
    NOR2X1 U29561 (.A1(n17326), .A2(N11351), .ZN(N42433));
    NANDX1 U29562 (.A1(N3155), .A2(N7608), .ZN(N42434));
    NOR2X1 U29563 (.A1(N4571), .A2(N4637), .ZN(n42435));
    NOR2X1 U29564 (.A1(N7430), .A2(N6540), .ZN(N42436));
    NOR2X1 U29565 (.A1(N5702), .A2(n26257), .ZN(n42437));
    INVX1 U29566 (.I(N10366), .ZN(N42438));
    NANDX1 U29567 (.A1(n24571), .A2(n23790), .ZN(N42439));
    NOR2X1 U29568 (.A1(n16691), .A2(n29185), .ZN(N42440));
    INVX1 U29569 (.I(n25487), .ZN(N42441));
    INVX1 U29570 (.I(N55), .ZN(n42442));
    NANDX1 U29571 (.A1(n22663), .A2(N3184), .ZN(n42443));
    NOR2X1 U29572 (.A1(n13254), .A2(N9070), .ZN(n42444));
    NOR2X1 U29573 (.A1(N5347), .A2(N12224), .ZN(n42445));
    NANDX1 U29574 (.A1(n29158), .A2(n16795), .ZN(N42446));
    INVX1 U29575 (.I(n29432), .ZN(n42447));
    NANDX1 U29576 (.A1(n19551), .A2(N2808), .ZN(N42448));
    NOR2X1 U29577 (.A1(N4232), .A2(n18923), .ZN(N42449));
    INVX1 U29578 (.I(n24758), .ZN(N42450));
    NOR2X1 U29579 (.A1(N11065), .A2(N11832), .ZN(N42451));
    INVX1 U29580 (.I(n28810), .ZN(n42452));
    NANDX1 U29581 (.A1(N2518), .A2(n23094), .ZN(N42453));
    NANDX1 U29582 (.A1(n27112), .A2(n15619), .ZN(n42454));
    INVX1 U29583 (.I(N9270), .ZN(n42455));
    NOR2X1 U29584 (.A1(N4408), .A2(N2778), .ZN(n42456));
    NANDX1 U29585 (.A1(N5193), .A2(N11153), .ZN(N42457));
    NOR2X1 U29586 (.A1(N10548), .A2(N5467), .ZN(N42458));
    NANDX1 U29587 (.A1(N11893), .A2(n13578), .ZN(N42459));
    NANDX1 U29588 (.A1(N241), .A2(n17809), .ZN(N42460));
    NANDX1 U29589 (.A1(n17652), .A2(N12430), .ZN(N42461));
    NANDX1 U29590 (.A1(n17277), .A2(N12822), .ZN(N42462));
    NOR2X1 U29591 (.A1(N4510), .A2(n27800), .ZN(N42463));
    NANDX1 U29592 (.A1(n27604), .A2(n19955), .ZN(N42464));
    INVX1 U29593 (.I(n13085), .ZN(N42465));
    INVX1 U29594 (.I(n14913), .ZN(N42466));
    INVX1 U29595 (.I(N8261), .ZN(n42467));
    INVX1 U29596 (.I(n23161), .ZN(N42468));
    NANDX1 U29597 (.A1(n17404), .A2(N3384), .ZN(N42469));
    INVX1 U29598 (.I(N11431), .ZN(N42470));
    NANDX1 U29599 (.A1(n24453), .A2(n25009), .ZN(N42471));
    INVX1 U29600 (.I(n13254), .ZN(N42472));
    INVX1 U29601 (.I(N3869), .ZN(N42473));
    NANDX1 U29602 (.A1(n13670), .A2(N2853), .ZN(n42474));
    NANDX1 U29603 (.A1(n26491), .A2(n20444), .ZN(N42475));
    INVX1 U29604 (.I(N12715), .ZN(N42476));
    NANDX1 U29605 (.A1(n15841), .A2(N2532), .ZN(N42477));
    NOR2X1 U29606 (.A1(n28925), .A2(n17824), .ZN(n42478));
    NOR2X1 U29607 (.A1(n17867), .A2(n26084), .ZN(n42479));
    NOR2X1 U29608 (.A1(N10890), .A2(n28098), .ZN(N42480));
    NOR2X1 U29609 (.A1(N2834), .A2(n29219), .ZN(n42481));
    INVX1 U29610 (.I(n15872), .ZN(N42482));
    INVX1 U29611 (.I(n15172), .ZN(N42483));
    NOR2X1 U29612 (.A1(n25349), .A2(n27851), .ZN(N42484));
    NANDX1 U29613 (.A1(n14678), .A2(N11384), .ZN(n42485));
    NOR2X1 U29614 (.A1(N9845), .A2(N7737), .ZN(n42486));
    NOR2X1 U29615 (.A1(n28219), .A2(n20451), .ZN(N42487));
    NANDX1 U29616 (.A1(n13922), .A2(N11543), .ZN(N42488));
    NANDX1 U29617 (.A1(N1270), .A2(n29366), .ZN(n42489));
    INVX1 U29618 (.I(N7697), .ZN(n42490));
    NANDX1 U29619 (.A1(n18676), .A2(N7147), .ZN(N42491));
    NOR2X1 U29620 (.A1(n27545), .A2(N9981), .ZN(N42492));
    INVX1 U29621 (.I(n17708), .ZN(N42493));
    NOR2X1 U29622 (.A1(N11571), .A2(N2742), .ZN(N42494));
    NOR2X1 U29623 (.A1(n25481), .A2(N456), .ZN(n42495));
    NOR2X1 U29624 (.A1(n28719), .A2(N400), .ZN(N42496));
    NOR2X1 U29625 (.A1(n27124), .A2(n26834), .ZN(n42497));
    NANDX1 U29626 (.A1(n25205), .A2(N5709), .ZN(N42498));
    INVX1 U29627 (.I(n27687), .ZN(N42499));
    INVX1 U29628 (.I(N12146), .ZN(N42500));
    INVX1 U29629 (.I(N5041), .ZN(n42501));
    INVX1 U29630 (.I(n25214), .ZN(N42502));
    NOR2X1 U29631 (.A1(N5015), .A2(N2224), .ZN(N42503));
    NOR2X1 U29632 (.A1(n21120), .A2(N765), .ZN(n42504));
    INVX1 U29633 (.I(N8691), .ZN(N42505));
    NANDX1 U29634 (.A1(n26174), .A2(n30130), .ZN(n42506));
    NOR2X1 U29635 (.A1(n21517), .A2(N448), .ZN(n42507));
    NANDX1 U29636 (.A1(n20098), .A2(n19545), .ZN(N42508));
    INVX1 U29637 (.I(N5646), .ZN(n42509));
    INVX1 U29638 (.I(N4419), .ZN(n42510));
    INVX1 U29639 (.I(n21950), .ZN(n42511));
    NOR2X1 U29640 (.A1(n16961), .A2(n27761), .ZN(N42512));
    NANDX1 U29641 (.A1(N4341), .A2(N2664), .ZN(N42513));
    NOR2X1 U29642 (.A1(n18115), .A2(N10138), .ZN(n42514));
    NOR2X1 U29643 (.A1(n20338), .A2(n18006), .ZN(N42515));
    NOR2X1 U29644 (.A1(n21102), .A2(n13911), .ZN(N42516));
    INVX1 U29645 (.I(N6142), .ZN(N42517));
    NANDX1 U29646 (.A1(n19309), .A2(n24087), .ZN(n42518));
    INVX1 U29647 (.I(N8318), .ZN(N42519));
    NANDX1 U29648 (.A1(n28682), .A2(n27862), .ZN(n42520));
    NOR2X1 U29649 (.A1(N4190), .A2(N2527), .ZN(n42521));
    NANDX1 U29650 (.A1(n23601), .A2(n13037), .ZN(N42522));
    NOR2X1 U29651 (.A1(N10424), .A2(N10661), .ZN(N42523));
    NANDX1 U29652 (.A1(N3325), .A2(n13324), .ZN(N42524));
    NANDX1 U29653 (.A1(n21439), .A2(n23462), .ZN(n42525));
    NANDX1 U29654 (.A1(N201), .A2(n30028), .ZN(n42526));
    INVX1 U29655 (.I(N9863), .ZN(N42527));
    INVX1 U29656 (.I(n22216), .ZN(N42528));
    NANDX1 U29657 (.A1(N12308), .A2(n30086), .ZN(N42529));
    NANDX1 U29658 (.A1(n20892), .A2(N8266), .ZN(n42530));
    NOR2X1 U29659 (.A1(n19437), .A2(N5990), .ZN(N42531));
    NANDX1 U29660 (.A1(n23626), .A2(n27215), .ZN(N42532));
    NANDX1 U29661 (.A1(N5650), .A2(N10114), .ZN(n42533));
    INVX1 U29662 (.I(N4634), .ZN(N42534));
    INVX1 U29663 (.I(N9709), .ZN(N42535));
    NANDX1 U29664 (.A1(N3961), .A2(n19735), .ZN(n42536));
    INVX1 U29665 (.I(n15983), .ZN(n42537));
    NOR2X1 U29666 (.A1(n18158), .A2(n15873), .ZN(n42538));
    NOR2X1 U29667 (.A1(n28020), .A2(n18235), .ZN(n42539));
    NANDX1 U29668 (.A1(N2448), .A2(N405), .ZN(n42540));
    NANDX1 U29669 (.A1(N961), .A2(n21297), .ZN(N42541));
    NOR2X1 U29670 (.A1(n25060), .A2(n29294), .ZN(N42542));
    INVX1 U29671 (.I(n28916), .ZN(n42543));
    NANDX1 U29672 (.A1(N2647), .A2(n24208), .ZN(n42544));
    INVX1 U29673 (.I(N1322), .ZN(N42545));
    INVX1 U29674 (.I(n21626), .ZN(n42546));
    NANDX1 U29675 (.A1(n29531), .A2(n18145), .ZN(N42547));
    NOR2X1 U29676 (.A1(N7689), .A2(N5965), .ZN(N42548));
    NOR2X1 U29677 (.A1(n26956), .A2(N12683), .ZN(N42549));
    NOR2X1 U29678 (.A1(N7547), .A2(n29263), .ZN(n42550));
    NOR2X1 U29679 (.A1(N10353), .A2(N1573), .ZN(N42551));
    NOR2X1 U29680 (.A1(N1668), .A2(n21232), .ZN(N42552));
    INVX1 U29681 (.I(N1248), .ZN(N42553));
    NOR2X1 U29682 (.A1(n21107), .A2(n25515), .ZN(N42554));
    NANDX1 U29683 (.A1(N2313), .A2(n16723), .ZN(n42555));
    NOR2X1 U29684 (.A1(N7866), .A2(n18044), .ZN(N42556));
    NOR2X1 U29685 (.A1(n18052), .A2(N10001), .ZN(n42557));
    NOR2X1 U29686 (.A1(N6059), .A2(n13178), .ZN(n42558));
    INVX1 U29687 (.I(N584), .ZN(N42559));
    NANDX1 U29688 (.A1(n17105), .A2(n13266), .ZN(n42560));
    INVX1 U29689 (.I(n13212), .ZN(N42561));
    INVX1 U29690 (.I(N84), .ZN(N42562));
    NOR2X1 U29691 (.A1(N2525), .A2(N739), .ZN(N42563));
    NANDX1 U29692 (.A1(n23756), .A2(n22689), .ZN(N42564));
    NANDX1 U29693 (.A1(N9772), .A2(n13659), .ZN(N42565));
    NOR2X1 U29694 (.A1(N1826), .A2(N4532), .ZN(n42566));
    INVX1 U29695 (.I(n18087), .ZN(n42567));
    NANDX1 U29696 (.A1(N3606), .A2(N12593), .ZN(n42568));
    INVX1 U29697 (.I(N2167), .ZN(N42569));
    NOR2X1 U29698 (.A1(n25068), .A2(n15344), .ZN(n42570));
    NOR2X1 U29699 (.A1(n25651), .A2(n17543), .ZN(N42571));
    NANDX1 U29700 (.A1(n27478), .A2(n24635), .ZN(N42572));
    NANDX1 U29701 (.A1(N9732), .A2(n13280), .ZN(N42573));
    INVX1 U29702 (.I(N12256), .ZN(n42574));
    NOR2X1 U29703 (.A1(n18557), .A2(n24573), .ZN(N42575));
    NOR2X1 U29704 (.A1(n22156), .A2(n22905), .ZN(n42576));
    INVX1 U29705 (.I(n21133), .ZN(N42577));
    NOR2X1 U29706 (.A1(N1880), .A2(N6695), .ZN(N42578));
    NANDX1 U29707 (.A1(N2837), .A2(n28998), .ZN(N42579));
    NOR2X1 U29708 (.A1(n21846), .A2(N1028), .ZN(n42580));
    NANDX1 U29709 (.A1(N5337), .A2(n16371), .ZN(N42581));
    NANDX1 U29710 (.A1(n19548), .A2(n22474), .ZN(N42582));
    INVX1 U29711 (.I(n16888), .ZN(n42583));
    NOR2X1 U29712 (.A1(N473), .A2(n26619), .ZN(N42584));
    NANDX1 U29713 (.A1(N5238), .A2(n27436), .ZN(N42585));
    INVX1 U29714 (.I(n23794), .ZN(N42586));
    NANDX1 U29715 (.A1(N5080), .A2(N4373), .ZN(N42587));
    INVX1 U29716 (.I(n21127), .ZN(N42588));
    INVX1 U29717 (.I(n27929), .ZN(N42589));
    INVX1 U29718 (.I(n20761), .ZN(N42590));
    INVX1 U29719 (.I(n14404), .ZN(N42591));
    NOR2X1 U29720 (.A1(N12863), .A2(n24810), .ZN(N42592));
    NANDX1 U29721 (.A1(N3050), .A2(N9), .ZN(n42593));
    NANDX1 U29722 (.A1(n27274), .A2(n19556), .ZN(n42594));
    NOR2X1 U29723 (.A1(n23668), .A2(N6307), .ZN(n42595));
    NOR2X1 U29724 (.A1(N12701), .A2(n21486), .ZN(N42596));
    INVX1 U29725 (.I(N6499), .ZN(n42597));
    INVX1 U29726 (.I(N6454), .ZN(n42598));
    NANDX1 U29727 (.A1(n17776), .A2(N11533), .ZN(N42599));
    NANDX1 U29728 (.A1(n20975), .A2(N2522), .ZN(n42600));
    NOR2X1 U29729 (.A1(n18766), .A2(n14089), .ZN(N42601));
    INVX1 U29730 (.I(n17796), .ZN(N42602));
    NANDX1 U29731 (.A1(N5960), .A2(N522), .ZN(N42603));
    NANDX1 U29732 (.A1(N3730), .A2(n22269), .ZN(n42604));
    NOR2X1 U29733 (.A1(n17871), .A2(n19406), .ZN(N42605));
    NANDX1 U29734 (.A1(n12909), .A2(N1497), .ZN(N42606));
    INVX1 U29735 (.I(n13479), .ZN(N42607));
    NANDX1 U29736 (.A1(n24763), .A2(N9982), .ZN(n42608));
    NOR2X1 U29737 (.A1(N1970), .A2(n16435), .ZN(N42609));
    INVX1 U29738 (.I(N8307), .ZN(N42610));
    INVX1 U29739 (.I(N9758), .ZN(N42611));
    INVX1 U29740 (.I(n19050), .ZN(N42612));
    NANDX1 U29741 (.A1(N6470), .A2(n21699), .ZN(n42613));
    INVX1 U29742 (.I(n24265), .ZN(N42614));
    NANDX1 U29743 (.A1(n27908), .A2(n13347), .ZN(N42615));
    INVX1 U29744 (.I(N1501), .ZN(N42616));
    INVX1 U29745 (.I(N9192), .ZN(n42617));
    INVX1 U29746 (.I(n13445), .ZN(n42618));
    NANDX1 U29747 (.A1(n20840), .A2(N3502), .ZN(N42619));
    NOR2X1 U29748 (.A1(N4181), .A2(N6259), .ZN(N42620));
    NANDX1 U29749 (.A1(N2723), .A2(N4076), .ZN(n42621));
    INVX1 U29750 (.I(n19157), .ZN(N42622));
    INVX1 U29751 (.I(n14339), .ZN(n42623));
    NOR2X1 U29752 (.A1(N366), .A2(N2043), .ZN(N42624));
    NOR2X1 U29753 (.A1(N5839), .A2(N8512), .ZN(n42625));
    NOR2X1 U29754 (.A1(N9089), .A2(N2640), .ZN(n42626));
    NANDX1 U29755 (.A1(n25557), .A2(N4547), .ZN(n42627));
    NOR2X1 U29756 (.A1(n27057), .A2(N10025), .ZN(N42628));
    NANDX1 U29757 (.A1(N4851), .A2(n23469), .ZN(N42629));
    NANDX1 U29758 (.A1(n14251), .A2(n26970), .ZN(N42630));
    NANDX1 U29759 (.A1(N6992), .A2(n21790), .ZN(N42631));
    NOR2X1 U29760 (.A1(N9714), .A2(n25865), .ZN(N42632));
    NOR2X1 U29761 (.A1(n28870), .A2(N5034), .ZN(n42633));
    INVX1 U29762 (.I(N4280), .ZN(n42634));
    INVX1 U29763 (.I(N1783), .ZN(N42635));
    NANDX1 U29764 (.A1(N11238), .A2(n28993), .ZN(N42636));
    NOR2X1 U29765 (.A1(N8887), .A2(N1495), .ZN(n42637));
    NANDX1 U29766 (.A1(N4306), .A2(N6041), .ZN(N42638));
    NANDX1 U29767 (.A1(n19924), .A2(N4627), .ZN(N42639));
    INVX1 U29768 (.I(n13335), .ZN(n42640));
    INVX1 U29769 (.I(N884), .ZN(n42641));
    INVX1 U29770 (.I(N2050), .ZN(N42642));
    INVX1 U29771 (.I(N4440), .ZN(n42643));
    NANDX1 U29772 (.A1(n27272), .A2(n14154), .ZN(n42644));
    NANDX1 U29773 (.A1(N12674), .A2(N1447), .ZN(N42645));
    INVX1 U29774 (.I(N975), .ZN(N42646));
    INVX1 U29775 (.I(N7121), .ZN(n42647));
    NANDX1 U29776 (.A1(N11723), .A2(N6919), .ZN(n42648));
    NANDX1 U29777 (.A1(N10998), .A2(N4366), .ZN(N42649));
    NANDX1 U29778 (.A1(N12164), .A2(N8671), .ZN(N42650));
    NANDX1 U29779 (.A1(N1242), .A2(n17155), .ZN(N42651));
    INVX1 U29780 (.I(n17560), .ZN(n42652));
    NANDX1 U29781 (.A1(n26248), .A2(n18443), .ZN(N42653));
    NOR2X1 U29782 (.A1(n16858), .A2(n24770), .ZN(n42654));
    NOR2X1 U29783 (.A1(n29257), .A2(N10465), .ZN(N42655));
    NANDX1 U29784 (.A1(N7247), .A2(N11699), .ZN(n42656));
    INVX1 U29785 (.I(N8968), .ZN(N42657));
    NANDX1 U29786 (.A1(n19385), .A2(N4649), .ZN(n42658));
    NANDX1 U29787 (.A1(N970), .A2(N128), .ZN(N42659));
    NOR2X1 U29788 (.A1(N11967), .A2(N4493), .ZN(n42660));
    NANDX1 U29789 (.A1(N12692), .A2(N1724), .ZN(n42661));
    INVX1 U29790 (.I(n13933), .ZN(N42662));
    NOR2X1 U29791 (.A1(n19086), .A2(n20053), .ZN(n42663));
    NANDX1 U29792 (.A1(N3757), .A2(N8359), .ZN(N42664));
    INVX1 U29793 (.I(N9176), .ZN(N42665));
    INVX1 U29794 (.I(N3651), .ZN(n42666));
    NANDX1 U29795 (.A1(N2016), .A2(n15864), .ZN(N42667));
    NANDX1 U29796 (.A1(n13715), .A2(N10825), .ZN(n42668));
    INVX1 U29797 (.I(n14948), .ZN(n42669));
    NOR2X1 U29798 (.A1(N6278), .A2(n18938), .ZN(n42670));
    NOR2X1 U29799 (.A1(N6405), .A2(N1662), .ZN(N42671));
    INVX1 U29800 (.I(n29595), .ZN(N42672));
    NOR2X1 U29801 (.A1(n21519), .A2(N1182), .ZN(N42673));
    INVX1 U29802 (.I(N5315), .ZN(n42674));
    NANDX1 U29803 (.A1(N11889), .A2(n25367), .ZN(n42675));
    NOR2X1 U29804 (.A1(n15645), .A2(n22286), .ZN(n42676));
    INVX1 U29805 (.I(n24820), .ZN(n42677));
    INVX1 U29806 (.I(n21473), .ZN(n42678));
    NOR2X1 U29807 (.A1(n15853), .A2(N7199), .ZN(N42679));
    INVX1 U29808 (.I(n18128), .ZN(n42680));
    NOR2X1 U29809 (.A1(N8709), .A2(N2938), .ZN(N42681));
    NOR2X1 U29810 (.A1(N3547), .A2(N10437), .ZN(N42682));
    NANDX1 U29811 (.A1(n28650), .A2(N12098), .ZN(N42683));
    NOR2X1 U29812 (.A1(n28107), .A2(N6847), .ZN(N42684));
    NOR2X1 U29813 (.A1(n17849), .A2(N11089), .ZN(N42685));
    NANDX1 U29814 (.A1(n26469), .A2(n22977), .ZN(N42686));
    NANDX1 U29815 (.A1(N1304), .A2(n27182), .ZN(N42687));
    NOR2X1 U29816 (.A1(n19126), .A2(n21865), .ZN(N42688));
    INVX1 U29817 (.I(N10462), .ZN(n42689));
    NOR2X1 U29818 (.A1(N10487), .A2(N6221), .ZN(n42690));
    INVX1 U29819 (.I(n28614), .ZN(N42691));
    NOR2X1 U29820 (.A1(N6311), .A2(n20113), .ZN(n42692));
    NOR2X1 U29821 (.A1(n28556), .A2(n19110), .ZN(N42693));
    INVX1 U29822 (.I(n27068), .ZN(n42694));
    NANDX1 U29823 (.A1(N1002), .A2(n13598), .ZN(n42695));
    NOR2X1 U29824 (.A1(N4727), .A2(n20008), .ZN(n42696));
    NOR2X1 U29825 (.A1(n21025), .A2(n16339), .ZN(n42697));
    INVX1 U29826 (.I(N2416), .ZN(N42698));
    INVX1 U29827 (.I(n27585), .ZN(N42699));
    INVX1 U29828 (.I(n13890), .ZN(N42700));
    NANDX1 U29829 (.A1(n19424), .A2(n24351), .ZN(N42701));
    NANDX1 U29830 (.A1(n29911), .A2(N435), .ZN(N42702));
    INVX1 U29831 (.I(n16948), .ZN(N42703));
    NOR2X1 U29832 (.A1(N2310), .A2(n25621), .ZN(N42704));
    NANDX1 U29833 (.A1(N728), .A2(n14593), .ZN(n42705));
    NOR2X1 U29834 (.A1(n16356), .A2(N4223), .ZN(n42706));
    NOR2X1 U29835 (.A1(n18515), .A2(N699), .ZN(n42707));
    INVX1 U29836 (.I(N8385), .ZN(N42708));
    NANDX1 U29837 (.A1(N2352), .A2(n13284), .ZN(n42709));
    NANDX1 U29838 (.A1(n23465), .A2(n19487), .ZN(N42710));
    NANDX1 U29839 (.A1(N6678), .A2(N3240), .ZN(N42711));
    INVX1 U29840 (.I(n26102), .ZN(n42712));
    INVX1 U29841 (.I(n19642), .ZN(N42713));
    NOR2X1 U29842 (.A1(N5146), .A2(n15641), .ZN(N42714));
    NOR2X1 U29843 (.A1(N6945), .A2(n17950), .ZN(n42715));
    INVX1 U29844 (.I(N5325), .ZN(n42716));
    NANDX1 U29845 (.A1(N11322), .A2(n22500), .ZN(N42717));
    INVX1 U29846 (.I(N4106), .ZN(N42718));
    INVX1 U29847 (.I(N532), .ZN(N42719));
    NOR2X1 U29848 (.A1(N10565), .A2(N8916), .ZN(n42720));
    NOR2X1 U29849 (.A1(N1477), .A2(N10761), .ZN(N42721));
    INVX1 U29850 (.I(n24942), .ZN(n42722));
    INVX1 U29851 (.I(n19485), .ZN(N42723));
    INVX1 U29852 (.I(n22047), .ZN(N42724));
    INVX1 U29853 (.I(n16144), .ZN(N42725));
    INVX1 U29854 (.I(n18795), .ZN(N42726));
    NOR2X1 U29855 (.A1(N1767), .A2(n22996), .ZN(N42727));
    NOR2X1 U29856 (.A1(N8712), .A2(N10808), .ZN(n42728));
    INVX1 U29857 (.I(N2597), .ZN(N42729));
    INVX1 U29858 (.I(N9738), .ZN(N42730));
    NOR2X1 U29859 (.A1(n18762), .A2(n13843), .ZN(N42731));
    INVX1 U29860 (.I(N7854), .ZN(N42732));
    NOR2X1 U29861 (.A1(N11883), .A2(N5331), .ZN(N42733));
    NOR2X1 U29862 (.A1(N1920), .A2(n16091), .ZN(N42734));
    NOR2X1 U29863 (.A1(n26861), .A2(N4761), .ZN(n42735));
    NOR2X1 U29864 (.A1(n16904), .A2(n15369), .ZN(n42736));
    NOR2X1 U29865 (.A1(n21608), .A2(N11990), .ZN(N42737));
    NOR2X1 U29866 (.A1(n22050), .A2(n13756), .ZN(n42738));
    NOR2X1 U29867 (.A1(n23737), .A2(N11028), .ZN(N42739));
    NANDX1 U29868 (.A1(n22153), .A2(N2186), .ZN(N42740));
    NOR2X1 U29869 (.A1(N1753), .A2(N4404), .ZN(N42741));
    NANDX1 U29870 (.A1(N4157), .A2(N5722), .ZN(N42742));
    INVX1 U29871 (.I(n30062), .ZN(n42743));
    NOR2X1 U29872 (.A1(N7263), .A2(n16018), .ZN(n42744));
    NOR2X1 U29873 (.A1(n23353), .A2(N8086), .ZN(N42745));
    INVX1 U29874 (.I(n28114), .ZN(N42746));
    NOR2X1 U29875 (.A1(n28970), .A2(N1906), .ZN(N42747));
    NOR2X1 U29876 (.A1(n20440), .A2(n13895), .ZN(N42748));
    NANDX1 U29877 (.A1(N12352), .A2(n16211), .ZN(n42749));
    INVX1 U29878 (.I(N5951), .ZN(n42750));
    NOR2X1 U29879 (.A1(N2080), .A2(n28103), .ZN(n42751));
    NANDX1 U29880 (.A1(N276), .A2(n18417), .ZN(n42752));
    NOR2X1 U29881 (.A1(n24492), .A2(N11134), .ZN(N42753));
    NANDX1 U29882 (.A1(n26424), .A2(n29756), .ZN(N42754));
    NANDX1 U29883 (.A1(N3550), .A2(N4197), .ZN(N42755));
    NANDX1 U29884 (.A1(n26902), .A2(N12282), .ZN(N42756));
    NANDX1 U29885 (.A1(n13439), .A2(n20482), .ZN(N42757));
    NOR2X1 U29886 (.A1(n15344), .A2(n20689), .ZN(N42758));
    NOR2X1 U29887 (.A1(n17799), .A2(n20260), .ZN(n42759));
    NANDX1 U29888 (.A1(N3873), .A2(N612), .ZN(N42760));
    NANDX1 U29889 (.A1(N8233), .A2(N2691), .ZN(n42761));
    NOR2X1 U29890 (.A1(n14778), .A2(n21664), .ZN(n42762));
    INVX1 U29891 (.I(n14287), .ZN(N42763));
    INVX1 U29892 (.I(n27998), .ZN(N42764));
    NOR2X1 U29893 (.A1(N866), .A2(n27616), .ZN(N42765));
    NANDX1 U29894 (.A1(N4415), .A2(n20373), .ZN(N42766));
    NOR2X1 U29895 (.A1(n19877), .A2(n21216), .ZN(n42767));
    NOR2X1 U29896 (.A1(N3179), .A2(N11560), .ZN(N42768));
    NOR2X1 U29897 (.A1(N7083), .A2(N2111), .ZN(N42769));
    NANDX1 U29898 (.A1(n24882), .A2(N10931), .ZN(n42770));
    INVX1 U29899 (.I(n28754), .ZN(N42771));
    NANDX1 U29900 (.A1(N10532), .A2(n25547), .ZN(n42772));
    INVX1 U29901 (.I(n20419), .ZN(N42773));
    INVX1 U29902 (.I(n13019), .ZN(N42774));
    INVX1 U29903 (.I(n24473), .ZN(N42775));
    NANDX1 U29904 (.A1(N5007), .A2(N2413), .ZN(N42776));
    NANDX1 U29905 (.A1(n21184), .A2(N10445), .ZN(N42777));
    NOR2X1 U29906 (.A1(n30117), .A2(n15076), .ZN(N42778));
    INVX1 U29907 (.I(n21195), .ZN(N42779));
    INVX1 U29908 (.I(n23053), .ZN(N42780));
    NOR2X1 U29909 (.A1(n19031), .A2(n18696), .ZN(N42781));
    NOR2X1 U29910 (.A1(n26186), .A2(n13440), .ZN(N42782));
    NANDX1 U29911 (.A1(N1917), .A2(N617), .ZN(n42783));
    INVX1 U29912 (.I(N12448), .ZN(N42784));
    NANDX1 U29913 (.A1(n25814), .A2(n21428), .ZN(N42785));
    NANDX1 U29914 (.A1(n27393), .A2(n17135), .ZN(N42786));
    INVX1 U29915 (.I(N3413), .ZN(N42787));
    NOR2X1 U29916 (.A1(n21657), .A2(n29134), .ZN(n42788));
    NOR2X1 U29917 (.A1(n20662), .A2(n29131), .ZN(N42789));
    NANDX1 U29918 (.A1(N5601), .A2(n18868), .ZN(n42790));
    INVX1 U29919 (.I(n22534), .ZN(N42791));
    NOR2X1 U29920 (.A1(N2661), .A2(n30125), .ZN(n42792));
    NOR2X1 U29921 (.A1(n14647), .A2(n14735), .ZN(n42793));
    INVX1 U29922 (.I(N7426), .ZN(N42794));
    INVX1 U29923 (.I(N10218), .ZN(N42795));
    NANDX1 U29924 (.A1(n17660), .A2(N6243), .ZN(N42796));
    NANDX1 U29925 (.A1(N8950), .A2(N1016), .ZN(N42797));
    NOR2X1 U29926 (.A1(n14645), .A2(N8821), .ZN(n42798));
    INVX1 U29927 (.I(n25346), .ZN(N42799));
    NOR2X1 U29928 (.A1(n14346), .A2(n15655), .ZN(n42800));
    INVX1 U29929 (.I(N1901), .ZN(N42801));
    NANDX1 U29930 (.A1(n15163), .A2(n20768), .ZN(N42802));
    NOR2X1 U29931 (.A1(n26258), .A2(n21112), .ZN(N42803));
    NANDX1 U29932 (.A1(n14806), .A2(n28712), .ZN(N42804));
    NOR2X1 U29933 (.A1(n29540), .A2(n19614), .ZN(N42805));
    NANDX1 U29934 (.A1(n16054), .A2(n29831), .ZN(n42806));
    INVX1 U29935 (.I(N3576), .ZN(n42807));
    NOR2X1 U29936 (.A1(N4132), .A2(N1086), .ZN(N42808));
    NOR2X1 U29937 (.A1(n16069), .A2(n15730), .ZN(N42809));
    NOR2X1 U29938 (.A1(n19979), .A2(n29636), .ZN(N42810));
    NANDX1 U29939 (.A1(n22886), .A2(n15153), .ZN(N42811));
    INVX1 U29940 (.I(n24786), .ZN(n42812));
    NOR2X1 U29941 (.A1(n17959), .A2(N3977), .ZN(N42813));
    INVX1 U29942 (.I(N2640), .ZN(N42814));
    INVX1 U29943 (.I(n20107), .ZN(N42815));
    NOR2X1 U29944 (.A1(N12223), .A2(n20521), .ZN(N42816));
    INVX1 U29945 (.I(n20398), .ZN(N42817));
    NANDX1 U29946 (.A1(N2764), .A2(N8652), .ZN(N42818));
    NANDX1 U29947 (.A1(n25037), .A2(N3149), .ZN(n42819));
    INVX1 U29948 (.I(n14683), .ZN(N42820));
    INVX1 U29949 (.I(n15130), .ZN(N42821));
    NANDX1 U29950 (.A1(n28951), .A2(n23669), .ZN(N42822));
    NOR2X1 U29951 (.A1(n22184), .A2(N4978), .ZN(N42823));
    NOR2X1 U29952 (.A1(n13541), .A2(n18324), .ZN(N42824));
    INVX1 U29953 (.I(n20061), .ZN(N42825));
    INVX1 U29954 (.I(N5906), .ZN(N42826));
    NOR2X1 U29955 (.A1(n24510), .A2(n26012), .ZN(n42827));
    NOR2X1 U29956 (.A1(N6596), .A2(N4956), .ZN(n42828));
    INVX1 U29957 (.I(n15554), .ZN(n42829));
    NANDX1 U29958 (.A1(N6741), .A2(n24205), .ZN(N42830));
    NOR2X1 U29959 (.A1(n20339), .A2(n15915), .ZN(N42831));
    NOR2X1 U29960 (.A1(N4884), .A2(n21834), .ZN(n42832));
    INVX1 U29961 (.I(n23857), .ZN(N42833));
    NOR2X1 U29962 (.A1(n24528), .A2(N12191), .ZN(n42834));
    NOR2X1 U29963 (.A1(n29505), .A2(N4238), .ZN(n42835));
    NOR2X1 U29964 (.A1(N6253), .A2(N5941), .ZN(n42836));
    NANDX1 U29965 (.A1(n17114), .A2(N407), .ZN(N42837));
    NOR2X1 U29966 (.A1(N11486), .A2(n14980), .ZN(N42838));
    NANDX1 U29967 (.A1(N6642), .A2(n19935), .ZN(n42839));
    NOR2X1 U29968 (.A1(n22195), .A2(n23113), .ZN(n42840));
    INVX1 U29969 (.I(N4824), .ZN(n42841));
    NANDX1 U29970 (.A1(n22725), .A2(n20738), .ZN(N42842));
    NANDX1 U29971 (.A1(n27608), .A2(N995), .ZN(N42843));
    NOR2X1 U29972 (.A1(N9888), .A2(N10203), .ZN(n42844));
    INVX1 U29973 (.I(n22078), .ZN(N42845));
    NANDX1 U29974 (.A1(n13005), .A2(n14877), .ZN(N42846));
    INVX1 U29975 (.I(N7818), .ZN(N42847));
    INVX1 U29976 (.I(n15350), .ZN(N42848));
    NOR2X1 U29977 (.A1(N9785), .A2(n19889), .ZN(N42849));
    NOR2X1 U29978 (.A1(n13325), .A2(N11557), .ZN(N42850));
    INVX1 U29979 (.I(n21820), .ZN(n42851));
    NANDX1 U29980 (.A1(n23676), .A2(n14795), .ZN(N42852));
    NOR2X1 U29981 (.A1(n28499), .A2(n24576), .ZN(N42853));
    NANDX1 U29982 (.A1(N7660), .A2(N12827), .ZN(N42854));
    INVX1 U29983 (.I(N8655), .ZN(N42855));
    NANDX1 U29984 (.A1(N9534), .A2(N7418), .ZN(n42856));
    INVX1 U29985 (.I(n20172), .ZN(N42857));
    INVX1 U29986 (.I(n28577), .ZN(n42858));
    NANDX1 U29987 (.A1(n29505), .A2(N6257), .ZN(N42859));
    NOR2X1 U29988 (.A1(n14717), .A2(N1050), .ZN(N42860));
    NOR2X1 U29989 (.A1(n23166), .A2(n26026), .ZN(n42861));
    NANDX1 U29990 (.A1(N4586), .A2(N8809), .ZN(n42862));
    INVX1 U29991 (.I(N11788), .ZN(N42863));
    NOR2X1 U29992 (.A1(n20996), .A2(N2678), .ZN(N42864));
    NANDX1 U29993 (.A1(N3995), .A2(N4853), .ZN(n42865));
    NANDX1 U29994 (.A1(n16821), .A2(N4498), .ZN(N42866));
    NOR2X1 U29995 (.A1(n18756), .A2(n14031), .ZN(n42867));
    NANDX1 U29996 (.A1(N4191), .A2(N4066), .ZN(N42868));
    NOR2X1 U29997 (.A1(N2630), .A2(n27674), .ZN(N42869));
    NANDX1 U29998 (.A1(n27584), .A2(N11825), .ZN(n42870));
    NANDX1 U29999 (.A1(n17194), .A2(n13019), .ZN(N42871));
    NOR2X1 U30000 (.A1(n13083), .A2(n27537), .ZN(N42872));
    INVX1 U30001 (.I(N10452), .ZN(n42873));
    NOR2X1 U30002 (.A1(N5422), .A2(N1360), .ZN(N42874));
    NOR2X1 U30003 (.A1(n26797), .A2(n20767), .ZN(N42875));
    NOR2X1 U30004 (.A1(N1512), .A2(n17696), .ZN(N42876));
    NOR2X1 U30005 (.A1(N6010), .A2(N11840), .ZN(n42877));
    INVX1 U30006 (.I(N8601), .ZN(n42878));
    NOR2X1 U30007 (.A1(n26780), .A2(N1227), .ZN(n42879));
    NOR2X1 U30008 (.A1(n17970), .A2(n28901), .ZN(N42880));
    INVX1 U30009 (.I(n15417), .ZN(n42881));
    NANDX1 U30010 (.A1(n22599), .A2(N2473), .ZN(N42882));
    NOR2X1 U30011 (.A1(n23088), .A2(N4116), .ZN(n42883));
    INVX1 U30012 (.I(n16722), .ZN(N42884));
    INVX1 U30013 (.I(n13167), .ZN(N42885));
    NANDX1 U30014 (.A1(n15927), .A2(N7625), .ZN(n42886));
    INVX1 U30015 (.I(n25254), .ZN(N42887));
    NOR2X1 U30016 (.A1(N8876), .A2(N1373), .ZN(N42888));
    NOR2X1 U30017 (.A1(n14885), .A2(n13212), .ZN(N42889));
    INVX1 U30018 (.I(n23485), .ZN(n42890));
    NANDX1 U30019 (.A1(n24961), .A2(n24712), .ZN(n42891));
    INVX1 U30020 (.I(N12793), .ZN(N42892));
    NOR2X1 U30021 (.A1(n14210), .A2(n16770), .ZN(N42893));
    NANDX1 U30022 (.A1(N6671), .A2(N7804), .ZN(N42894));
    INVX1 U30023 (.I(n18319), .ZN(n42895));
    INVX1 U30024 (.I(N2781), .ZN(N42896));
    NANDX1 U30025 (.A1(n15047), .A2(n15947), .ZN(N42897));
    INVX1 U30026 (.I(n19535), .ZN(N42898));
    NOR2X1 U30027 (.A1(n22971), .A2(n14651), .ZN(n42899));
    NOR2X1 U30028 (.A1(N1709), .A2(n16024), .ZN(N42900));
    NOR2X1 U30029 (.A1(n16593), .A2(n17796), .ZN(n42901));
    INVX1 U30030 (.I(n28639), .ZN(N42902));
    NANDX1 U30031 (.A1(n24202), .A2(N11774), .ZN(N42903));
    NOR2X1 U30032 (.A1(n25555), .A2(N12370), .ZN(N42904));
    NANDX1 U30033 (.A1(N12188), .A2(n23553), .ZN(N42905));
    INVX1 U30034 (.I(N8552), .ZN(N42906));
    NANDX1 U30035 (.A1(N6783), .A2(N9031), .ZN(n42907));
    INVX1 U30036 (.I(N11686), .ZN(N42908));
    INVX1 U30037 (.I(n24054), .ZN(N42909));
    INVX1 U30038 (.I(N2036), .ZN(N42910));
    NANDX1 U30039 (.A1(N8688), .A2(N5247), .ZN(N42911));
    NANDX1 U30040 (.A1(n29094), .A2(N9831), .ZN(N42912));
    NANDX1 U30041 (.A1(N4111), .A2(n16188), .ZN(N42913));
    NOR2X1 U30042 (.A1(n21310), .A2(n26278), .ZN(N42914));
    NANDX1 U30043 (.A1(N2946), .A2(N5301), .ZN(N42915));
    NOR2X1 U30044 (.A1(n15315), .A2(N9973), .ZN(n42916));
    NOR2X1 U30045 (.A1(n27428), .A2(n28574), .ZN(N42917));
    INVX1 U30046 (.I(n14057), .ZN(N42918));
    NOR2X1 U30047 (.A1(n16751), .A2(n22164), .ZN(N42919));
    INVX1 U30048 (.I(n29389), .ZN(N42920));
    NANDX1 U30049 (.A1(N9880), .A2(N1287), .ZN(N42921));
    NOR2X1 U30050 (.A1(n18567), .A2(n25231), .ZN(N42922));
    NANDX1 U30051 (.A1(N6085), .A2(N4925), .ZN(N42923));
    INVX1 U30052 (.I(N10195), .ZN(N42924));
    NANDX1 U30053 (.A1(n26526), .A2(N1367), .ZN(N42925));
    INVX1 U30054 (.I(N10831), .ZN(N42926));
    NANDX1 U30055 (.A1(N11113), .A2(N9252), .ZN(N42927));
    NANDX1 U30056 (.A1(N9646), .A2(N8420), .ZN(N42928));
    NANDX1 U30057 (.A1(n26780), .A2(N4701), .ZN(N42929));
    INVX1 U30058 (.I(N1862), .ZN(n42930));
    NOR2X1 U30059 (.A1(n18819), .A2(n26025), .ZN(n42931));
    NOR2X1 U30060 (.A1(n23460), .A2(N5767), .ZN(N42932));
    NOR2X1 U30061 (.A1(N11272), .A2(n12895), .ZN(n42933));
    NOR2X1 U30062 (.A1(N7721), .A2(n18979), .ZN(n42934));
    NANDX1 U30063 (.A1(n25308), .A2(n29173), .ZN(n42935));
    INVX1 U30064 (.I(N10257), .ZN(N42936));
    NOR2X1 U30065 (.A1(n14611), .A2(n21088), .ZN(n42937));
    NANDX1 U30066 (.A1(n14285), .A2(n18900), .ZN(N42938));
    NOR2X1 U30067 (.A1(n23930), .A2(n15880), .ZN(N42939));
    INVX1 U30068 (.I(N9134), .ZN(N42940));
    NOR2X1 U30069 (.A1(n29548), .A2(N10995), .ZN(N42941));
    NOR2X1 U30070 (.A1(n18230), .A2(n25580), .ZN(N42942));
    NANDX1 U30071 (.A1(N113), .A2(n19907), .ZN(n42943));
    NANDX1 U30072 (.A1(n30082), .A2(N2664), .ZN(N42944));
    NOR2X1 U30073 (.A1(N7666), .A2(N10203), .ZN(n42945));
    INVX1 U30074 (.I(n21534), .ZN(N42946));
    NANDX1 U30075 (.A1(n22392), .A2(N1653), .ZN(N42947));
    NANDX1 U30076 (.A1(N6865), .A2(N11301), .ZN(n42948));
    NOR2X1 U30077 (.A1(N9710), .A2(n18761), .ZN(N42949));
    NANDX1 U30078 (.A1(n22201), .A2(n23202), .ZN(N42950));
    NOR2X1 U30079 (.A1(N1197), .A2(n13644), .ZN(N42951));
    INVX1 U30080 (.I(N752), .ZN(N42952));
    INVX1 U30081 (.I(n16406), .ZN(N42953));
    INVX1 U30082 (.I(n23813), .ZN(n42954));
    INVX1 U30083 (.I(n16100), .ZN(n42955));
    NOR2X1 U30084 (.A1(N5024), .A2(N7325), .ZN(N42956));
    NANDX1 U30085 (.A1(N1250), .A2(n17527), .ZN(N42957));
    NANDX1 U30086 (.A1(N11344), .A2(N3887), .ZN(N42958));
    NOR2X1 U30087 (.A1(N1558), .A2(n20784), .ZN(N42959));
    NOR2X1 U30088 (.A1(N12858), .A2(n19516), .ZN(n42960));
    NANDX1 U30089 (.A1(n20180), .A2(n15526), .ZN(n42961));
    NOR2X1 U30090 (.A1(n13244), .A2(n14292), .ZN(n42962));
    NANDX1 U30091 (.A1(n15448), .A2(N12469), .ZN(N42963));
    NANDX1 U30092 (.A1(n18106), .A2(n28874), .ZN(N42964));
    NOR2X1 U30093 (.A1(N11782), .A2(n22514), .ZN(N42965));
    NOR2X1 U30094 (.A1(n14282), .A2(n27538), .ZN(N42966));
    NOR2X1 U30095 (.A1(N1111), .A2(n17348), .ZN(n42967));
    NANDX1 U30096 (.A1(n20230), .A2(n28692), .ZN(n42968));
    NOR2X1 U30097 (.A1(N1467), .A2(n18810), .ZN(N42969));
    INVX1 U30098 (.I(n19705), .ZN(n42970));
    NANDX1 U30099 (.A1(N4515), .A2(N6076), .ZN(N42971));
    NANDX1 U30100 (.A1(n20040), .A2(n14648), .ZN(N42972));
    INVX1 U30101 (.I(N4195), .ZN(N42973));
    INVX1 U30102 (.I(n27522), .ZN(N42974));
    INVX1 U30103 (.I(N12056), .ZN(n42975));
    INVX1 U30104 (.I(N3960), .ZN(n42976));
    NOR2X1 U30105 (.A1(n15832), .A2(n26474), .ZN(N42977));
    NOR2X1 U30106 (.A1(n18674), .A2(N12435), .ZN(n42978));
    NANDX1 U30107 (.A1(n19784), .A2(n29782), .ZN(N42979));
    NANDX1 U30108 (.A1(n28575), .A2(n16897), .ZN(n42980));
    NANDX1 U30109 (.A1(n30041), .A2(n24267), .ZN(n42981));
    NANDX1 U30110 (.A1(n19608), .A2(n14358), .ZN(n42982));
    NANDX1 U30111 (.A1(n14244), .A2(n13188), .ZN(N42983));
    NANDX1 U30112 (.A1(n17452), .A2(n25262), .ZN(N42984));
    NANDX1 U30113 (.A1(n18989), .A2(N11207), .ZN(N42985));
    NOR2X1 U30114 (.A1(N907), .A2(n26696), .ZN(N42986));
    NOR2X1 U30115 (.A1(n26932), .A2(N952), .ZN(N42987));
    INVX1 U30116 (.I(n22754), .ZN(N42988));
    INVX1 U30117 (.I(N899), .ZN(N42989));
    INVX1 U30118 (.I(n27970), .ZN(N42990));
    INVX1 U30119 (.I(n19377), .ZN(N42991));
    NOR2X1 U30120 (.A1(N6001), .A2(N16), .ZN(n42992));
    NANDX1 U30121 (.A1(n18829), .A2(n25927), .ZN(N42993));
    INVX1 U30122 (.I(N3049), .ZN(N42994));
    NANDX1 U30123 (.A1(N7145), .A2(n16236), .ZN(N42995));
    INVX1 U30124 (.I(n13158), .ZN(N42996));
    NOR2X1 U30125 (.A1(N10792), .A2(N2009), .ZN(N42997));
    NOR2X1 U30126 (.A1(n29098), .A2(N2915), .ZN(n42998));
    NOR2X1 U30127 (.A1(N2528), .A2(n18407), .ZN(N42999));
    NANDX1 U30128 (.A1(n21130), .A2(N11023), .ZN(n43000));
    NOR2X1 U30129 (.A1(n22028), .A2(n13977), .ZN(N43001));
    NOR2X1 U30130 (.A1(n29830), .A2(N3216), .ZN(N43002));
    NANDX1 U30131 (.A1(N5694), .A2(n21929), .ZN(N43003));
    INVX1 U30132 (.I(n13083), .ZN(N43004));
    NOR2X1 U30133 (.A1(n18694), .A2(n16131), .ZN(N43005));
    NANDX1 U30134 (.A1(n25839), .A2(n20927), .ZN(N43006));
    NANDX1 U30135 (.A1(N8859), .A2(n20848), .ZN(n43007));
    INVX1 U30136 (.I(N10867), .ZN(N43008));
    INVX1 U30137 (.I(n28515), .ZN(N43009));
    NANDX1 U30138 (.A1(N9522), .A2(n19603), .ZN(N43010));
    NOR2X1 U30139 (.A1(N6719), .A2(n29293), .ZN(N43011));
    NOR2X1 U30140 (.A1(N12102), .A2(N9745), .ZN(N43012));
    NOR2X1 U30141 (.A1(n26755), .A2(N9437), .ZN(N43013));
    INVX1 U30142 (.I(n26239), .ZN(N43014));
    NANDX1 U30143 (.A1(N6437), .A2(n21894), .ZN(n43015));
    NANDX1 U30144 (.A1(n24155), .A2(N10451), .ZN(N43016));
    NOR2X1 U30145 (.A1(n26512), .A2(n24850), .ZN(n43017));
    INVX1 U30146 (.I(n15138), .ZN(N43018));
    INVX1 U30147 (.I(n14403), .ZN(N43019));
    NOR2X1 U30148 (.A1(N2998), .A2(n16239), .ZN(N43020));
    NANDX1 U30149 (.A1(n24037), .A2(n14322), .ZN(N43021));
    INVX1 U30150 (.I(N3208), .ZN(N43022));
    NANDX1 U30151 (.A1(n27510), .A2(N12100), .ZN(n43023));
    INVX1 U30152 (.I(N7117), .ZN(N43024));
    INVX1 U30153 (.I(N6881), .ZN(n43025));
    NANDX1 U30154 (.A1(n19476), .A2(N2982), .ZN(N43026));
    INVX1 U30155 (.I(n14473), .ZN(N43027));
    INVX1 U30156 (.I(N6879), .ZN(N43028));
    INVX1 U30157 (.I(N12447), .ZN(N43029));
    NOR2X1 U30158 (.A1(n23562), .A2(N7159), .ZN(N43030));
    INVX1 U30159 (.I(N8562), .ZN(N43031));
    INVX1 U30160 (.I(n13422), .ZN(n43032));
    INVX1 U30161 (.I(n20985), .ZN(N43033));
    NANDX1 U30162 (.A1(n20428), .A2(N3445), .ZN(N43034));
    NANDX1 U30163 (.A1(n30083), .A2(N6653), .ZN(N43035));
    INVX1 U30164 (.I(n27455), .ZN(N43036));
    NANDX1 U30165 (.A1(N10829), .A2(n23132), .ZN(N43037));
    NOR2X1 U30166 (.A1(N6270), .A2(N9548), .ZN(N43038));
    NANDX1 U30167 (.A1(N9251), .A2(n29791), .ZN(N43039));
    NANDX1 U30168 (.A1(N11248), .A2(n25230), .ZN(N43040));
    NOR2X1 U30169 (.A1(N12255), .A2(N11996), .ZN(N43041));
    INVX1 U30170 (.I(N7975), .ZN(N43042));
    NOR2X1 U30171 (.A1(N10809), .A2(n25962), .ZN(N43043));
    NANDX1 U30172 (.A1(N11046), .A2(n16810), .ZN(N43044));
    NANDX1 U30173 (.A1(n20034), .A2(n20254), .ZN(n43045));
    NOR2X1 U30174 (.A1(n19979), .A2(n15467), .ZN(n43046));
    INVX1 U30175 (.I(N5858), .ZN(N43047));
    NANDX1 U30176 (.A1(n22139), .A2(n28989), .ZN(N43048));
    NANDX1 U30177 (.A1(n28408), .A2(n27097), .ZN(N43049));
    INVX1 U30178 (.I(n26220), .ZN(N43050));
    INVX1 U30179 (.I(N9680), .ZN(N43051));
    INVX1 U30180 (.I(N10404), .ZN(N43052));
    NANDX1 U30181 (.A1(N8145), .A2(N10960), .ZN(n43053));
    NANDX1 U30182 (.A1(n16119), .A2(N3277), .ZN(N43054));
    INVX1 U30183 (.I(N11944), .ZN(n43055));
    NOR2X1 U30184 (.A1(N1027), .A2(n17314), .ZN(n43056));
    INVX1 U30185 (.I(n21060), .ZN(N43057));
    NOR2X1 U30186 (.A1(N2140), .A2(n29599), .ZN(N43058));
    NOR2X1 U30187 (.A1(n24888), .A2(n24017), .ZN(N43059));
    NANDX1 U30188 (.A1(n16889), .A2(N11430), .ZN(N43060));
    NOR2X1 U30189 (.A1(n15160), .A2(N8389), .ZN(N43061));
    INVX1 U30190 (.I(N11242), .ZN(N43062));
    NOR2X1 U30191 (.A1(N8110), .A2(N7132), .ZN(N43063));
    INVX1 U30192 (.I(n26612), .ZN(N43064));
    NOR2X1 U30193 (.A1(N3486), .A2(n17224), .ZN(N43065));
    NOR2X1 U30194 (.A1(n25460), .A2(N7205), .ZN(N43066));
    NANDX1 U30195 (.A1(n23035), .A2(N8231), .ZN(n43067));
    INVX1 U30196 (.I(n21689), .ZN(N43068));
    NANDX1 U30197 (.A1(n15065), .A2(n23828), .ZN(N43069));
    INVX1 U30198 (.I(n15083), .ZN(N43070));
    NOR2X1 U30199 (.A1(n18451), .A2(n26441), .ZN(N43071));
    NANDX1 U30200 (.A1(n29880), .A2(n26965), .ZN(N43072));
    NOR2X1 U30201 (.A1(n26829), .A2(n25395), .ZN(n43073));
    NOR2X1 U30202 (.A1(N8952), .A2(n22065), .ZN(n43074));
    INVX1 U30203 (.I(n20176), .ZN(N43075));
    NOR2X1 U30204 (.A1(N8381), .A2(n23662), .ZN(n43076));
    NOR2X1 U30205 (.A1(n28336), .A2(N7545), .ZN(n43077));
    INVX1 U30206 (.I(n18658), .ZN(n43078));
    NOR2X1 U30207 (.A1(N9620), .A2(N7595), .ZN(N43079));
    NOR2X1 U30208 (.A1(n16031), .A2(N11220), .ZN(N43080));
    INVX1 U30209 (.I(N10465), .ZN(N43081));
    NANDX1 U30210 (.A1(N82), .A2(n28915), .ZN(N43082));
    INVX1 U30211 (.I(n24110), .ZN(N43083));
    NOR2X1 U30212 (.A1(n26693), .A2(n21720), .ZN(N43084));
    NANDX1 U30213 (.A1(N10511), .A2(N435), .ZN(n43085));
    NANDX1 U30214 (.A1(N2439), .A2(n23676), .ZN(n43086));
    NANDX1 U30215 (.A1(n20977), .A2(N1919), .ZN(n43087));
    INVX1 U30216 (.I(n15163), .ZN(N43088));
    NOR2X1 U30217 (.A1(N2529), .A2(n27991), .ZN(N43089));
    NANDX1 U30218 (.A1(N10229), .A2(n26172), .ZN(n43090));
    NANDX1 U30219 (.A1(n20920), .A2(N12065), .ZN(N43091));
    NOR2X1 U30220 (.A1(N2424), .A2(n22529), .ZN(n43092));
    NANDX1 U30221 (.A1(N2505), .A2(N9867), .ZN(N43093));
    NANDX1 U30222 (.A1(n26614), .A2(n27084), .ZN(N43094));
    NANDX1 U30223 (.A1(N6758), .A2(N10856), .ZN(N43095));
    NOR2X1 U30224 (.A1(n25890), .A2(n22277), .ZN(n43096));
    INVX1 U30225 (.I(n19428), .ZN(n43097));
    NANDX1 U30226 (.A1(n18204), .A2(N9908), .ZN(N43098));
    INVX1 U30227 (.I(N3229), .ZN(n43099));
    NANDX1 U30228 (.A1(n28507), .A2(n19781), .ZN(n43100));
    INVX1 U30229 (.I(N8598), .ZN(n43101));
    NOR2X1 U30230 (.A1(N9409), .A2(n18079), .ZN(n43102));
    NOR2X1 U30231 (.A1(N12679), .A2(n20502), .ZN(n43103));
    NANDX1 U30232 (.A1(N12114), .A2(n23006), .ZN(n43104));
    INVX1 U30233 (.I(n22716), .ZN(N43105));
    INVX1 U30234 (.I(n22904), .ZN(N43106));
    INVX1 U30235 (.I(n14801), .ZN(N43107));
    NANDX1 U30236 (.A1(n24661), .A2(N10553), .ZN(N43108));
    NANDX1 U30237 (.A1(n21888), .A2(n18541), .ZN(n43109));
    NOR2X1 U30238 (.A1(N9955), .A2(n28448), .ZN(N43110));
    NOR2X1 U30239 (.A1(N1744), .A2(n27033), .ZN(N43111));
    NOR2X1 U30240 (.A1(N10085), .A2(n21513), .ZN(N43112));
    INVX1 U30241 (.I(n14460), .ZN(N43113));
    NANDX1 U30242 (.A1(n17504), .A2(n19461), .ZN(N43114));
    NANDX1 U30243 (.A1(N7868), .A2(n16853), .ZN(N43115));
    INVX1 U30244 (.I(n19434), .ZN(N43116));
    NANDX1 U30245 (.A1(n25413), .A2(n16038), .ZN(N43117));
    NOR2X1 U30246 (.A1(N2270), .A2(N701), .ZN(N43118));
    INVX1 U30247 (.I(n15491), .ZN(N43119));
    INVX1 U30248 (.I(n19337), .ZN(n43120));
    NOR2X1 U30249 (.A1(n18355), .A2(N4516), .ZN(N43121));
    NOR2X1 U30250 (.A1(N5226), .A2(n27111), .ZN(N43122));
    NANDX1 U30251 (.A1(N2121), .A2(n17939), .ZN(N43123));
    NANDX1 U30252 (.A1(n23633), .A2(n17364), .ZN(N43124));
    INVX1 U30253 (.I(n12978), .ZN(N43125));
    NOR2X1 U30254 (.A1(N9928), .A2(n15001), .ZN(N43126));
    INVX1 U30255 (.I(n15341), .ZN(N43127));
    NANDX1 U30256 (.A1(N9152), .A2(n16574), .ZN(n43128));
    NOR2X1 U30257 (.A1(n13751), .A2(N10572), .ZN(n43129));
    INVX1 U30258 (.I(N3012), .ZN(N43130));
    NANDX1 U30259 (.A1(n19294), .A2(N2826), .ZN(N43131));
    INVX1 U30260 (.I(n15096), .ZN(N43132));
    NOR2X1 U30261 (.A1(n27863), .A2(n20852), .ZN(n43133));
    NOR2X1 U30262 (.A1(n24837), .A2(n28352), .ZN(N43134));
    INVX1 U30263 (.I(N1199), .ZN(N43135));
    NANDX1 U30264 (.A1(n17841), .A2(n18562), .ZN(n43136));
    NOR2X1 U30265 (.A1(N681), .A2(N413), .ZN(N43137));
    NOR2X1 U30266 (.A1(N4242), .A2(n20268), .ZN(n43138));
    INVX1 U30267 (.I(N10501), .ZN(N43139));
    INVX1 U30268 (.I(n13790), .ZN(N43140));
    NOR2X1 U30269 (.A1(N1593), .A2(n12923), .ZN(N43141));
    NOR2X1 U30270 (.A1(n23303), .A2(n16934), .ZN(N43142));
    NANDX1 U30271 (.A1(n26128), .A2(N10144), .ZN(N43143));
    INVX1 U30272 (.I(n24429), .ZN(N43144));
    INVX1 U30273 (.I(n29502), .ZN(N43145));
    NANDX1 U30274 (.A1(n21267), .A2(n16277), .ZN(N43146));
    NANDX1 U30275 (.A1(n22465), .A2(N9197), .ZN(N43147));
    NOR2X1 U30276 (.A1(n29587), .A2(n22722), .ZN(N43148));
    NOR2X1 U30277 (.A1(n29999), .A2(N4598), .ZN(n43149));
    NANDX1 U30278 (.A1(N8690), .A2(N1814), .ZN(N43150));
    NANDX1 U30279 (.A1(n26669), .A2(N4165), .ZN(N43151));
    INVX1 U30280 (.I(n16823), .ZN(N43152));
    INVX1 U30281 (.I(N145), .ZN(N43153));
    NANDX1 U30282 (.A1(n22581), .A2(n23836), .ZN(N43154));
    INVX1 U30283 (.I(N2587), .ZN(n43155));
    NANDX1 U30284 (.A1(N7528), .A2(n29154), .ZN(N43156));
    INVX1 U30285 (.I(N5345), .ZN(N43157));
    NANDX1 U30286 (.A1(N6551), .A2(n27508), .ZN(N43158));
    NANDX1 U30287 (.A1(N4309), .A2(N7237), .ZN(N43159));
    NOR2X1 U30288 (.A1(n27030), .A2(n17783), .ZN(n43160));
    NOR2X1 U30289 (.A1(N1490), .A2(n21132), .ZN(N43161));
    INVX1 U30290 (.I(n22001), .ZN(N43162));
    NOR2X1 U30291 (.A1(n12961), .A2(n26165), .ZN(N43163));
    NOR2X1 U30292 (.A1(n18344), .A2(N1675), .ZN(N43164));
    INVX1 U30293 (.I(n16892), .ZN(N43165));
    INVX1 U30294 (.I(N1692), .ZN(N43166));
    INVX1 U30295 (.I(n26842), .ZN(n43167));
    NANDX1 U30296 (.A1(N7518), .A2(n14419), .ZN(N43168));
    NOR2X1 U30297 (.A1(N1423), .A2(N4565), .ZN(N43169));
    INVX1 U30298 (.I(n17491), .ZN(N43170));
    INVX1 U30299 (.I(N12432), .ZN(n43171));
    NANDX1 U30300 (.A1(n25053), .A2(n28022), .ZN(n43172));
    NOR2X1 U30301 (.A1(n14094), .A2(n29511), .ZN(N43173));
    NOR2X1 U30302 (.A1(N386), .A2(n21374), .ZN(N43174));
    NOR2X1 U30303 (.A1(N1907), .A2(N5963), .ZN(N43175));
    NOR2X1 U30304 (.A1(N8811), .A2(N7637), .ZN(n43176));
    INVX1 U30305 (.I(n25702), .ZN(n43177));
    NANDX1 U30306 (.A1(n21563), .A2(n25692), .ZN(n43178));
    INVX1 U30307 (.I(N2724), .ZN(N43179));
    INVX1 U30308 (.I(n20136), .ZN(N43180));
    NOR2X1 U30309 (.A1(N11753), .A2(n13261), .ZN(N43181));
    INVX1 U30310 (.I(n29244), .ZN(n43182));
    NANDX1 U30311 (.A1(N1973), .A2(n23833), .ZN(N43183));
    INVX1 U30312 (.I(n29994), .ZN(n43184));
    INVX1 U30313 (.I(N5126), .ZN(n43185));
    INVX1 U30314 (.I(N5255), .ZN(n43186));
    NANDX1 U30315 (.A1(n27862), .A2(N9285), .ZN(N43187));
    NANDX1 U30316 (.A1(N3687), .A2(n21163), .ZN(N43188));
    NOR2X1 U30317 (.A1(n30022), .A2(N10897), .ZN(N43189));
    INVX1 U30318 (.I(n20337), .ZN(N43190));
    NOR2X1 U30319 (.A1(N3165), .A2(n26054), .ZN(N43191));
    NOR2X1 U30320 (.A1(n13495), .A2(n16052), .ZN(N43192));
    NANDX1 U30321 (.A1(n25248), .A2(n29313), .ZN(N43193));
    NOR2X1 U30322 (.A1(n24354), .A2(N6732), .ZN(N43194));
    NANDX1 U30323 (.A1(N6610), .A2(n27901), .ZN(n43195));
    NOR2X1 U30324 (.A1(N1239), .A2(N2889), .ZN(N43196));
    NOR2X1 U30325 (.A1(n25191), .A2(n27098), .ZN(N43197));
    INVX1 U30326 (.I(N4338), .ZN(n43198));
    NOR2X1 U30327 (.A1(N8610), .A2(n14061), .ZN(n43199));
    INVX1 U30328 (.I(N8494), .ZN(N43200));
    INVX1 U30329 (.I(n24034), .ZN(n43201));
    NOR2X1 U30330 (.A1(n27279), .A2(n15760), .ZN(n43202));
    NOR2X1 U30331 (.A1(n20885), .A2(n29254), .ZN(N43203));
    NOR2X1 U30332 (.A1(n18787), .A2(n24364), .ZN(N43204));
    INVX1 U30333 (.I(n17669), .ZN(n43205));
    NOR2X1 U30334 (.A1(N947), .A2(n18523), .ZN(N43206));
    INVX1 U30335 (.I(n28847), .ZN(N43207));
    NANDX1 U30336 (.A1(N3550), .A2(n20297), .ZN(n43208));
    INVX1 U30337 (.I(n28740), .ZN(n43209));
    INVX1 U30338 (.I(N1217), .ZN(N43210));
    NANDX1 U30339 (.A1(n17453), .A2(N9826), .ZN(N43211));
    NANDX1 U30340 (.A1(n22437), .A2(N6880), .ZN(N43212));
    NANDX1 U30341 (.A1(N4895), .A2(n24270), .ZN(n43213));
    NOR2X1 U30342 (.A1(n20654), .A2(N7439), .ZN(N43214));
    NANDX1 U30343 (.A1(n19770), .A2(n25357), .ZN(N43215));
    INVX1 U30344 (.I(n13997), .ZN(N43216));
    NOR2X1 U30345 (.A1(N1847), .A2(n21137), .ZN(n43217));
    NOR2X1 U30346 (.A1(n20370), .A2(n23448), .ZN(n43218));
    INVX1 U30347 (.I(n28163), .ZN(N43219));
    NANDX1 U30348 (.A1(N9388), .A2(n13018), .ZN(n43220));
    NANDX1 U30349 (.A1(n15205), .A2(N2795), .ZN(n43221));
    NOR2X1 U30350 (.A1(N2520), .A2(N1181), .ZN(N43222));
    NOR2X1 U30351 (.A1(n13518), .A2(N8060), .ZN(N43223));
    NANDX1 U30352 (.A1(n18412), .A2(N2192), .ZN(n43224));
    INVX1 U30353 (.I(N8928), .ZN(N43225));
    NANDX1 U30354 (.A1(N11911), .A2(n28697), .ZN(N43226));
    NOR2X1 U30355 (.A1(n26226), .A2(N1117), .ZN(n43227));
    NOR2X1 U30356 (.A1(n16633), .A2(N10815), .ZN(n43228));
    NOR2X1 U30357 (.A1(N6865), .A2(N4125), .ZN(n43229));
    INVX1 U30358 (.I(n23589), .ZN(N43230));
    NANDX1 U30359 (.A1(n27799), .A2(n25167), .ZN(n43231));
    NOR2X1 U30360 (.A1(N1427), .A2(n27961), .ZN(N43232));
    INVX1 U30361 (.I(n22644), .ZN(N43233));
    NOR2X1 U30362 (.A1(n16405), .A2(N6024), .ZN(N43234));
    NANDX1 U30363 (.A1(N5127), .A2(n24435), .ZN(n43235));
    NANDX1 U30364 (.A1(N10070), .A2(n21923), .ZN(N43236));
    INVX1 U30365 (.I(N10541), .ZN(N43237));
    NANDX1 U30366 (.A1(N8112), .A2(n25327), .ZN(N43238));
    INVX1 U30367 (.I(N9655), .ZN(n43239));
    NOR2X1 U30368 (.A1(N9535), .A2(N1579), .ZN(N43240));
    INVX1 U30369 (.I(n13660), .ZN(N43241));
    INVX1 U30370 (.I(N699), .ZN(N43242));
    NANDX1 U30371 (.A1(n17651), .A2(n14426), .ZN(N43243));
    NANDX1 U30372 (.A1(n19077), .A2(N12249), .ZN(N43244));
    NANDX1 U30373 (.A1(N11583), .A2(n29950), .ZN(N43245));
    NANDX1 U30374 (.A1(n17607), .A2(n25573), .ZN(N43246));
    NANDX1 U30375 (.A1(N465), .A2(n23387), .ZN(N43247));
    INVX1 U30376 (.I(n22388), .ZN(N43248));
    INVX1 U30377 (.I(N1218), .ZN(n43249));
    NANDX1 U30378 (.A1(n16063), .A2(n26544), .ZN(N43250));
    NOR2X1 U30379 (.A1(n25717), .A2(n26926), .ZN(n43251));
    INVX1 U30380 (.I(n15856), .ZN(N43252));
    INVX1 U30381 (.I(N11769), .ZN(N43253));
    INVX1 U30382 (.I(n23432), .ZN(n43254));
    NANDX1 U30383 (.A1(N11919), .A2(N7720), .ZN(N43255));
    NOR2X1 U30384 (.A1(N858), .A2(N8529), .ZN(N43256));
    NOR2X1 U30385 (.A1(N1002), .A2(N8341), .ZN(n43257));
    NANDX1 U30386 (.A1(N7169), .A2(n22474), .ZN(N43258));
    NOR2X1 U30387 (.A1(N7633), .A2(N4284), .ZN(N43259));
    INVX1 U30388 (.I(n18581), .ZN(N43260));
    INVX1 U30389 (.I(n19353), .ZN(n43261));
    NOR2X1 U30390 (.A1(n16859), .A2(N4320), .ZN(N43262));
    INVX1 U30391 (.I(N999), .ZN(N43263));
    NOR2X1 U30392 (.A1(N6558), .A2(n16855), .ZN(n43264));
    INVX1 U30393 (.I(N6887), .ZN(n43265));
    NOR2X1 U30394 (.A1(n17137), .A2(n29118), .ZN(N43266));
    NOR2X1 U30395 (.A1(n13417), .A2(N5242), .ZN(N43267));
    INVX1 U30396 (.I(n21946), .ZN(n43268));
    INVX1 U30397 (.I(N2022), .ZN(n43269));
    INVX1 U30398 (.I(n17432), .ZN(N43270));
    INVX1 U30399 (.I(n29882), .ZN(n43271));
    NANDX1 U30400 (.A1(N5384), .A2(N4028), .ZN(n43272));
    INVX1 U30401 (.I(N12525), .ZN(n43273));
    NANDX1 U30402 (.A1(N10665), .A2(n20960), .ZN(N43274));
    INVX1 U30403 (.I(N3546), .ZN(N43275));
    NOR2X1 U30404 (.A1(n22680), .A2(n23352), .ZN(n43276));
    INVX1 U30405 (.I(n28095), .ZN(N43277));
    INVX1 U30406 (.I(N8534), .ZN(n43278));
    INVX1 U30407 (.I(n22753), .ZN(N43279));
    NOR2X1 U30408 (.A1(n20683), .A2(N6033), .ZN(N43280));
    INVX1 U30409 (.I(n21703), .ZN(N43281));
    NANDX1 U30410 (.A1(n13473), .A2(n23725), .ZN(n43282));
    NOR2X1 U30411 (.A1(N767), .A2(n21475), .ZN(N43283));
    NANDX1 U30412 (.A1(N4080), .A2(n26858), .ZN(N43284));
    NOR2X1 U30413 (.A1(n25529), .A2(N9246), .ZN(N43285));
    INVX1 U30414 (.I(n24755), .ZN(n43286));
    NOR2X1 U30415 (.A1(N1207), .A2(n16861), .ZN(N43287));
    NOR2X1 U30416 (.A1(n23886), .A2(N10075), .ZN(N43288));
    INVX1 U30417 (.I(N10405), .ZN(N43289));
    NOR2X1 U30418 (.A1(N5338), .A2(N8046), .ZN(N43290));
    NOR2X1 U30419 (.A1(N12851), .A2(n17289), .ZN(n43291));
    NOR2X1 U30420 (.A1(N2727), .A2(N8854), .ZN(n43292));
    NANDX1 U30421 (.A1(n16199), .A2(n21139), .ZN(n43293));
    INVX1 U30422 (.I(N5526), .ZN(N43294));
    NANDX1 U30423 (.A1(n25497), .A2(N9606), .ZN(N43295));
    NANDX1 U30424 (.A1(N199), .A2(n23695), .ZN(n43296));
    NANDX1 U30425 (.A1(n21300), .A2(N6873), .ZN(N43297));
    NANDX1 U30426 (.A1(n22506), .A2(n23733), .ZN(N43298));
    NANDX1 U30427 (.A1(N4815), .A2(N3670), .ZN(N43299));
    NOR2X1 U30428 (.A1(n15219), .A2(n19361), .ZN(N43300));
    NOR2X1 U30429 (.A1(N11825), .A2(n27667), .ZN(N43301));
    NOR2X1 U30430 (.A1(n29113), .A2(N11868), .ZN(N43302));
    INVX1 U30431 (.I(N7830), .ZN(n43303));
    INVX1 U30432 (.I(n24704), .ZN(n43304));
    INVX1 U30433 (.I(N2974), .ZN(N43305));
    NANDX1 U30434 (.A1(n30005), .A2(n17031), .ZN(N43306));
    NANDX1 U30435 (.A1(n27763), .A2(n17229), .ZN(N43307));
    NANDX1 U30436 (.A1(N4628), .A2(n27089), .ZN(N43308));
    INVX1 U30437 (.I(N259), .ZN(n43309));
    NOR2X1 U30438 (.A1(n29680), .A2(n21183), .ZN(N43310));
    INVX1 U30439 (.I(N3213), .ZN(n43311));
    NOR2X1 U30440 (.A1(n16612), .A2(N11134), .ZN(n43312));
    NOR2X1 U30441 (.A1(n28437), .A2(N8663), .ZN(N43313));
    NOR2X1 U30442 (.A1(n27412), .A2(n20530), .ZN(n43314));
    INVX1 U30443 (.I(n23802), .ZN(n43315));
    NOR2X1 U30444 (.A1(n29251), .A2(n29892), .ZN(N43316));
    NANDX1 U30445 (.A1(n17904), .A2(n29759), .ZN(N43317));
    NANDX1 U30446 (.A1(n16162), .A2(n15945), .ZN(N43318));
    NANDX1 U30447 (.A1(n15237), .A2(n20573), .ZN(N43319));
    NOR2X1 U30448 (.A1(N2486), .A2(N9392), .ZN(N43320));
    NANDX1 U30449 (.A1(N2028), .A2(N437), .ZN(N43321));
    NOR2X1 U30450 (.A1(n23938), .A2(N9211), .ZN(N43322));
    NANDX1 U30451 (.A1(N4934), .A2(n22353), .ZN(N43323));
    NOR2X1 U30452 (.A1(n13596), .A2(n29834), .ZN(n43324));
    NANDX1 U30453 (.A1(n22686), .A2(n15683), .ZN(n43325));
    INVX1 U30454 (.I(n21504), .ZN(n43326));
    NOR2X1 U30455 (.A1(n20959), .A2(N11857), .ZN(n43327));
    NANDX1 U30456 (.A1(N9141), .A2(n19240), .ZN(N43328));
    NANDX1 U30457 (.A1(n25086), .A2(n13714), .ZN(n43329));
    INVX1 U30458 (.I(N4082), .ZN(n43330));
    NOR2X1 U30459 (.A1(n13567), .A2(n13473), .ZN(n43331));
    NANDX1 U30460 (.A1(N4156), .A2(N2470), .ZN(N43332));
    NANDX1 U30461 (.A1(n28093), .A2(N11681), .ZN(n43333));
    INVX1 U30462 (.I(n21588), .ZN(N43334));
    NANDX1 U30463 (.A1(N118), .A2(n23744), .ZN(N43335));
    NOR2X1 U30464 (.A1(n27658), .A2(N4854), .ZN(N43336));
    NOR2X1 U30465 (.A1(n18725), .A2(n14918), .ZN(N43337));
    NOR2X1 U30466 (.A1(N9546), .A2(n26774), .ZN(N43338));
    NANDX1 U30467 (.A1(n18686), .A2(n15876), .ZN(N43339));
    NANDX1 U30468 (.A1(N2195), .A2(n18151), .ZN(N43340));
    NOR2X1 U30469 (.A1(n24974), .A2(N11851), .ZN(N43341));
    INVX1 U30470 (.I(n27007), .ZN(N43342));
    NOR2X1 U30471 (.A1(n26963), .A2(n29477), .ZN(N43343));
    NOR2X1 U30472 (.A1(n13479), .A2(n29718), .ZN(n43344));
    NOR2X1 U30473 (.A1(N4929), .A2(n22174), .ZN(N43345));
    INVX1 U30474 (.I(n17234), .ZN(n43346));
    NOR2X1 U30475 (.A1(n18380), .A2(n22087), .ZN(n43347));
    NOR2X1 U30476 (.A1(N6967), .A2(N6867), .ZN(N43348));
    NANDX1 U30477 (.A1(N5073), .A2(n22202), .ZN(N43349));
    NANDX1 U30478 (.A1(N12319), .A2(n26638), .ZN(N43350));
    INVX1 U30479 (.I(n14514), .ZN(N43351));
    INVX1 U30480 (.I(N8746), .ZN(N43352));
    NANDX1 U30481 (.A1(n15063), .A2(N1416), .ZN(N43353));
    INVX1 U30482 (.I(n27316), .ZN(N43354));
    NOR2X1 U30483 (.A1(N12818), .A2(n22111), .ZN(N43355));
    NOR2X1 U30484 (.A1(N12398), .A2(n24155), .ZN(N43356));
    NOR2X1 U30485 (.A1(N4434), .A2(N3438), .ZN(N43357));
    NOR2X1 U30486 (.A1(n18759), .A2(n21817), .ZN(n43358));
    INVX1 U30487 (.I(n29479), .ZN(n43359));
    INVX1 U30488 (.I(n17078), .ZN(n43360));
    NANDX1 U30489 (.A1(n22416), .A2(N9142), .ZN(N43361));
    INVX1 U30490 (.I(N4597), .ZN(N43362));
    NOR2X1 U30491 (.A1(N10664), .A2(N7671), .ZN(n43363));
    INVX1 U30492 (.I(n19410), .ZN(N43364));
    NANDX1 U30493 (.A1(N12477), .A2(N9386), .ZN(N43365));
    NOR2X1 U30494 (.A1(N9655), .A2(n14886), .ZN(n43366));
    NOR2X1 U30495 (.A1(N1629), .A2(N3727), .ZN(n43367));
    INVX1 U30496 (.I(n14344), .ZN(N43368));
    INVX1 U30497 (.I(n18570), .ZN(N43369));
    INVX1 U30498 (.I(N4319), .ZN(n43370));
    NOR2X1 U30499 (.A1(n28158), .A2(n14529), .ZN(n43371));
    NOR2X1 U30500 (.A1(n15364), .A2(n20167), .ZN(N43372));
    NANDX1 U30501 (.A1(n26340), .A2(n17869), .ZN(N43373));
    NOR2X1 U30502 (.A1(N799), .A2(N12072), .ZN(N43374));
    INVX1 U30503 (.I(n27168), .ZN(n43375));
    INVX1 U30504 (.I(N380), .ZN(N43376));
    INVX1 U30505 (.I(n21962), .ZN(N43377));
    NOR2X1 U30506 (.A1(n21671), .A2(n20177), .ZN(N43378));
    NANDX1 U30507 (.A1(n23410), .A2(N10366), .ZN(N43379));
    NOR2X1 U30508 (.A1(n26107), .A2(n24709), .ZN(N43380));
    NOR2X1 U30509 (.A1(N3100), .A2(N913), .ZN(N43381));
    INVX1 U30510 (.I(n28988), .ZN(N43382));
    NANDX1 U30511 (.A1(n17661), .A2(N1202), .ZN(N43383));
    INVX1 U30512 (.I(n26388), .ZN(N43384));
    NANDX1 U30513 (.A1(n17757), .A2(n14120), .ZN(n43385));
    INVX1 U30514 (.I(N7117), .ZN(N43386));
    NANDX1 U30515 (.A1(n17658), .A2(N4147), .ZN(N43387));
    NANDX1 U30516 (.A1(n18037), .A2(N6758), .ZN(N43388));
    NOR2X1 U30517 (.A1(n16363), .A2(n16989), .ZN(n43389));
    NOR2X1 U30518 (.A1(n29574), .A2(n28959), .ZN(N43390));
    NOR2X1 U30519 (.A1(n23633), .A2(n24928), .ZN(N43391));
    NOR2X1 U30520 (.A1(N3749), .A2(n16588), .ZN(N43392));
    INVX1 U30521 (.I(N6880), .ZN(N43393));
    NANDX1 U30522 (.A1(n13961), .A2(n13101), .ZN(N43394));
    NOR2X1 U30523 (.A1(N5379), .A2(n28050), .ZN(n43395));
    INVX1 U30524 (.I(N11696), .ZN(n43396));
    NANDX1 U30525 (.A1(n13675), .A2(n18812), .ZN(N43397));
    NOR2X1 U30526 (.A1(N1195), .A2(n22958), .ZN(n43398));
    NANDX1 U30527 (.A1(n19231), .A2(n18276), .ZN(N43399));
    INVX1 U30528 (.I(N5457), .ZN(N43400));
    NANDX1 U30529 (.A1(N8724), .A2(n23591), .ZN(N43401));
    NANDX1 U30530 (.A1(N2311), .A2(n17087), .ZN(N43402));
    NANDX1 U30531 (.A1(N9168), .A2(n20835), .ZN(N43403));
    INVX1 U30532 (.I(n16937), .ZN(N43404));
    INVX1 U30533 (.I(n15143), .ZN(n43405));
    NOR2X1 U30534 (.A1(n17937), .A2(n20342), .ZN(n43406));
    INVX1 U30535 (.I(n15849), .ZN(N43407));
    NOR2X1 U30536 (.A1(N6395), .A2(n16441), .ZN(n43408));
    NOR2X1 U30537 (.A1(n25206), .A2(n13086), .ZN(N43409));
    INVX1 U30538 (.I(N6588), .ZN(n43410));
    NOR2X1 U30539 (.A1(n19989), .A2(n13424), .ZN(N43411));
    NOR2X1 U30540 (.A1(n25445), .A2(N7112), .ZN(N43412));
    NOR2X1 U30541 (.A1(N7460), .A2(n18318), .ZN(N43413));
    NOR2X1 U30542 (.A1(n24546), .A2(n12876), .ZN(N43414));
    NOR2X1 U30543 (.A1(N3804), .A2(n24020), .ZN(n43415));
    INVX1 U30544 (.I(N8639), .ZN(N43416));
    INVX1 U30545 (.I(n28731), .ZN(N43417));
    INVX1 U30546 (.I(n17928), .ZN(N43418));
    NANDX1 U30547 (.A1(N847), .A2(n26696), .ZN(n43419));
    NOR2X1 U30548 (.A1(n17287), .A2(n26260), .ZN(N43420));
    INVX1 U30549 (.I(n18933), .ZN(N43421));
    NANDX1 U30550 (.A1(N8601), .A2(n30021), .ZN(N43422));
    NANDX1 U30551 (.A1(n22025), .A2(n25035), .ZN(N43423));
    INVX1 U30552 (.I(n17697), .ZN(N43424));
    NANDX1 U30553 (.A1(n19636), .A2(n24575), .ZN(N43425));
    NANDX1 U30554 (.A1(N2605), .A2(n26011), .ZN(N43426));
    INVX1 U30555 (.I(N6408), .ZN(n43427));
    INVX1 U30556 (.I(n20812), .ZN(N43428));
    NOR2X1 U30557 (.A1(N6041), .A2(n19405), .ZN(n43429));
    INVX1 U30558 (.I(n23968), .ZN(N43430));
    NOR2X1 U30559 (.A1(N892), .A2(N9088), .ZN(N43431));
    NOR2X1 U30560 (.A1(N6739), .A2(N5210), .ZN(N43432));
    NANDX1 U30561 (.A1(n25672), .A2(n13530), .ZN(N43433));
    NANDX1 U30562 (.A1(n14116), .A2(N262), .ZN(N43434));
    NOR2X1 U30563 (.A1(n27712), .A2(N999), .ZN(n43435));
    NOR2X1 U30564 (.A1(N3469), .A2(N9196), .ZN(n43436));
    INVX1 U30565 (.I(n22670), .ZN(N43437));
    INVX1 U30566 (.I(N7272), .ZN(N43438));
    NANDX1 U30567 (.A1(n18208), .A2(n15726), .ZN(N43439));
    NOR2X1 U30568 (.A1(N3117), .A2(n21766), .ZN(N43440));
    NANDX1 U30569 (.A1(n21859), .A2(n15597), .ZN(n43441));
    NANDX1 U30570 (.A1(n22750), .A2(n24684), .ZN(N43442));
    NANDX1 U30571 (.A1(n29489), .A2(n29893), .ZN(N43443));
    NOR2X1 U30572 (.A1(n13584), .A2(N1846), .ZN(N43444));
    NANDX1 U30573 (.A1(n16260), .A2(n20805), .ZN(n43445));
    NANDX1 U30574 (.A1(n13834), .A2(n21804), .ZN(N43446));
    NANDX1 U30575 (.A1(N5863), .A2(n19560), .ZN(N43447));
    NOR2X1 U30576 (.A1(n17093), .A2(N1222), .ZN(N43448));
    NANDX1 U30577 (.A1(n21163), .A2(n19429), .ZN(N43449));
    NANDX1 U30578 (.A1(N4468), .A2(N11106), .ZN(N43450));
    NANDX1 U30579 (.A1(n25876), .A2(N2828), .ZN(n43451));
    NOR2X1 U30580 (.A1(N11145), .A2(n14138), .ZN(N43452));
    NANDX1 U30581 (.A1(N4616), .A2(N2050), .ZN(n43453));
    NOR2X1 U30582 (.A1(N12484), .A2(n15633), .ZN(n43454));
    NOR2X1 U30583 (.A1(n20470), .A2(n20454), .ZN(N43455));
    NANDX1 U30584 (.A1(n20461), .A2(N4150), .ZN(N43456));
    INVX1 U30585 (.I(N7276), .ZN(N43457));
    NOR2X1 U30586 (.A1(n22295), .A2(n16928), .ZN(N43458));
    NOR2X1 U30587 (.A1(n23516), .A2(n22413), .ZN(N43459));
    NOR2X1 U30588 (.A1(N1369), .A2(n24925), .ZN(N43460));
    NANDX1 U30589 (.A1(N12474), .A2(N7626), .ZN(N43461));
    NOR2X1 U30590 (.A1(N3862), .A2(N5924), .ZN(N43462));
    NANDX1 U30591 (.A1(n18000), .A2(n28904), .ZN(N43463));
    INVX1 U30592 (.I(N8610), .ZN(n43464));
    INVX1 U30593 (.I(N823), .ZN(N43465));
    INVX1 U30594 (.I(N11768), .ZN(N43466));
    NOR2X1 U30595 (.A1(N3120), .A2(N4139), .ZN(N43467));
    INVX1 U30596 (.I(n25967), .ZN(N43468));
    INVX1 U30597 (.I(N7452), .ZN(N43469));
    INVX1 U30598 (.I(n17729), .ZN(N43470));
    NANDX1 U30599 (.A1(N10069), .A2(N11107), .ZN(n43471));
    INVX1 U30600 (.I(N5321), .ZN(N43472));
    NANDX1 U30601 (.A1(n16358), .A2(n15073), .ZN(N43473));
    NANDX1 U30602 (.A1(N3102), .A2(n31902), .ZN(N43474));
    NANDX1 U30603 (.A1(n34083), .A2(n14697), .ZN(n43475));
    INVX1 U30604 (.I(n23264), .ZN(N43476));
    NANDX1 U30605 (.A1(N3005), .A2(n39785), .ZN(N43477));
    NANDX1 U30606 (.A1(n28686), .A2(n26323), .ZN(N43478));
    INVX1 U30607 (.I(N10083), .ZN(N43479));
    NANDX1 U30608 (.A1(n22546), .A2(n31758), .ZN(N43480));
    INVX1 U30609 (.I(N3871), .ZN(N43481));
    NOR2X1 U30610 (.A1(N859), .A2(n25223), .ZN(N43482));
    INVX1 U30611 (.I(N507), .ZN(N43483));
    INVX1 U30612 (.I(N7645), .ZN(N43484));
    NOR2X1 U30613 (.A1(n29725), .A2(N12397), .ZN(N43485));
    INVX1 U30614 (.I(n32826), .ZN(N43486));
    INVX1 U30615 (.I(n34632), .ZN(N43487));
    INVX1 U30616 (.I(n15523), .ZN(N43488));
    INVX1 U30617 (.I(N3228), .ZN(N43489));
    INVX1 U30618 (.I(n24019), .ZN(N43490));
    NOR2X1 U30619 (.A1(n23480), .A2(N9232), .ZN(N43491));
    NOR2X1 U30620 (.A1(N1260), .A2(N8994), .ZN(N43492));
    NANDX1 U30621 (.A1(n13485), .A2(n40751), .ZN(N43493));
    NANDX1 U30622 (.A1(N7035), .A2(n32158), .ZN(N43494));
    NOR2X1 U30623 (.A1(n21937), .A2(n16374), .ZN(N43495));
    INVX1 U30624 (.I(N2152), .ZN(N43496));
    NOR2X1 U30625 (.A1(n42560), .A2(n31877), .ZN(N43497));
    INVX1 U30626 (.I(N3233), .ZN(N43498));
    NANDX1 U30627 (.A1(n26920), .A2(n27544), .ZN(N43499));
    NANDX1 U30628 (.A1(n42442), .A2(n15406), .ZN(N43500));
    NANDX1 U30629 (.A1(N2984), .A2(n39424), .ZN(N43501));
    INVX1 U30630 (.I(n16143), .ZN(N43502));
    INVX1 U30631 (.I(n32016), .ZN(N43503));
    INVX1 U30632 (.I(N3856), .ZN(N43504));
    NOR2X1 U30633 (.A1(n20566), .A2(n34286), .ZN(N43505));
    NANDX1 U30634 (.A1(n27601), .A2(n22971), .ZN(N43506));
    INVX1 U30635 (.I(N6065), .ZN(N43507));
    INVX1 U30636 (.I(n32284), .ZN(N43508));
    NANDX1 U30637 (.A1(n42722), .A2(n21052), .ZN(N43509));
    INVX1 U30638 (.I(n25344), .ZN(N43510));
    INVX1 U30639 (.I(n30362), .ZN(N43511));
    NOR2X1 U30640 (.A1(n41507), .A2(N10916), .ZN(N43512));
    INVX1 U30641 (.I(n13441), .ZN(N43513));
    NOR2X1 U30642 (.A1(n33575), .A2(n42544), .ZN(N43514));
    INVX1 U30643 (.I(N6245), .ZN(N43515));
    INVX1 U30644 (.I(n43185), .ZN(N43516));
    NANDX1 U30645 (.A1(n20622), .A2(N9741), .ZN(N43517));
    INVX1 U30646 (.I(N1116), .ZN(N43518));
    NANDX1 U30647 (.A1(N7699), .A2(n24086), .ZN(N43519));
    NOR2X1 U30648 (.A1(N3444), .A2(n42790), .ZN(N43520));
    INVX1 U30649 (.I(n34492), .ZN(N43521));
    NOR2X1 U30650 (.A1(n39911), .A2(N10472), .ZN(N43522));
    INVX1 U30651 (.I(N10402), .ZN(n43523));
    NANDX1 U30652 (.A1(N12061), .A2(N8436), .ZN(N43524));
    NOR2X1 U30653 (.A1(n42652), .A2(N11556), .ZN(N43525));
    NOR2X1 U30654 (.A1(n22434), .A2(N308), .ZN(N43526));
    NOR2X1 U30655 (.A1(n18358), .A2(n27394), .ZN(N43527));
    INVX1 U30656 (.I(n31683), .ZN(N43528));
    INVX1 U30657 (.I(N2954), .ZN(N43529));
    NANDX1 U30658 (.A1(n38810), .A2(n19080), .ZN(N43530));
    NOR2X1 U30659 (.A1(N9104), .A2(n15976), .ZN(N43531));
    NANDX1 U30660 (.A1(N8421), .A2(n34835), .ZN(N43532));
    NANDX1 U30661 (.A1(n40140), .A2(n20953), .ZN(N43533));
    NOR2X1 U30662 (.A1(n43410), .A2(n31354), .ZN(n43534));
    INVX1 U30663 (.I(N1678), .ZN(N43535));
    INVX1 U30664 (.I(n32241), .ZN(N43536));
    NOR2X1 U30665 (.A1(n41025), .A2(n14572), .ZN(N43537));
    INVX1 U30666 (.I(n41332), .ZN(N43538));
    NANDX1 U30667 (.A1(n31327), .A2(n25253), .ZN(n43539));
    NOR2X1 U30668 (.A1(N9217), .A2(n19475), .ZN(N43540));
    NOR2X1 U30669 (.A1(n20998), .A2(N4493), .ZN(N43541));
    NOR2X1 U30670 (.A1(n19837), .A2(n13596), .ZN(N43542));
    NOR2X1 U30671 (.A1(n22119), .A2(n22016), .ZN(n43543));
    INVX1 U30672 (.I(n15420), .ZN(N43544));
    NOR2X1 U30673 (.A1(n41288), .A2(N8872), .ZN(N43545));
    NOR2X1 U30674 (.A1(n18849), .A2(n32836), .ZN(N43546));
    NANDX1 U30675 (.A1(N4845), .A2(N11284), .ZN(N43547));
    INVX1 U30676 (.I(N2397), .ZN(N43548));
    NOR2X1 U30677 (.A1(n25997), .A2(N256), .ZN(N43549));
    NANDX1 U30678 (.A1(N3531), .A2(n15188), .ZN(N43550));
    INVX1 U30679 (.I(N12748), .ZN(N43551));
    NANDX1 U30680 (.A1(n16619), .A2(n23425), .ZN(N43552));
    NOR2X1 U30681 (.A1(n39937), .A2(n43261), .ZN(N43553));
    INVX1 U30682 (.I(n25438), .ZN(n43554));
    INVX1 U30683 (.I(N10653), .ZN(N43555));
    NOR2X1 U30684 (.A1(n16686), .A2(N8696), .ZN(N43556));
    INVX1 U30685 (.I(n15237), .ZN(n43557));
    INVX1 U30686 (.I(N8644), .ZN(N43558));
    NOR2X1 U30687 (.A1(n29167), .A2(n13489), .ZN(n43559));
    INVX1 U30688 (.I(n42193), .ZN(N43560));
    NANDX1 U30689 (.A1(n21099), .A2(n14397), .ZN(n43561));
    NOR2X1 U30690 (.A1(N1234), .A2(n17928), .ZN(N43562));
    INVX1 U30691 (.I(N3294), .ZN(N43563));
    INVX1 U30692 (.I(n24710), .ZN(n43564));
    NOR2X1 U30693 (.A1(n33459), .A2(n43224), .ZN(N43565));
    INVX1 U30694 (.I(n22927), .ZN(N43566));
    NOR2X1 U30695 (.A1(n21174), .A2(n24193), .ZN(N43567));
    INVX1 U30696 (.I(n13155), .ZN(N43568));
    NANDX1 U30697 (.A1(n30569), .A2(N2950), .ZN(N43569));
    NANDX1 U30698 (.A1(n26925), .A2(N11594), .ZN(N43570));
    INVX1 U30699 (.I(N2299), .ZN(N43571));
    INVX1 U30700 (.I(N2164), .ZN(N43572));
    NOR2X1 U30701 (.A1(n20326), .A2(n12942), .ZN(N43573));
    NANDX1 U30702 (.A1(n15826), .A2(n14175), .ZN(N43574));
    NANDX1 U30703 (.A1(n16194), .A2(N7148), .ZN(n43575));
    NOR2X1 U30704 (.A1(n30583), .A2(n16740), .ZN(N43576));
    NANDX1 U30705 (.A1(n30335), .A2(N12476), .ZN(N43577));
    INVX1 U30706 (.I(N8403), .ZN(N43578));
    NANDX1 U30707 (.A1(N6049), .A2(n30276), .ZN(N43579));
    NANDX1 U30708 (.A1(N3454), .A2(n17373), .ZN(N43580));
    INVX1 U30709 (.I(N5775), .ZN(N43581));
    NANDX1 U30710 (.A1(n40706), .A2(N12696), .ZN(n43582));
    NANDX1 U30711 (.A1(N1675), .A2(N4539), .ZN(N43583));
    NANDX1 U30712 (.A1(n22000), .A2(n17481), .ZN(N43584));
    INVX1 U30713 (.I(n27506), .ZN(n43585));
    NANDX1 U30714 (.A1(N11621), .A2(N227), .ZN(N43586));
    INVX1 U30715 (.I(n34357), .ZN(N43587));
    INVX1 U30716 (.I(n34902), .ZN(N43588));
    NOR2X1 U30717 (.A1(N7351), .A2(n37057), .ZN(N43589));
    NOR2X1 U30718 (.A1(N5434), .A2(n16913), .ZN(N43590));
    NOR2X1 U30719 (.A1(n35709), .A2(n43076), .ZN(N43591));
    INVX1 U30720 (.I(n42761), .ZN(N43592));
    NOR2X1 U30721 (.A1(n33893), .A2(N114), .ZN(n43593));
    NANDX1 U30722 (.A1(n36268), .A2(n36389), .ZN(N43594));
    INVX1 U30723 (.I(n40806), .ZN(N43595));
    INVX1 U30724 (.I(n28982), .ZN(N43596));
    INVX1 U30725 (.I(n18808), .ZN(N43597));
    INVX1 U30726 (.I(n15509), .ZN(N43598));
    NANDX1 U30727 (.A1(N2921), .A2(n33671), .ZN(N43599));
    NOR2X1 U30728 (.A1(n23410), .A2(n25100), .ZN(N43600));
    NANDX1 U30729 (.A1(n20440), .A2(N8364), .ZN(N43601));
    NANDX1 U30730 (.A1(n25873), .A2(n14956), .ZN(N43602));
    NANDX1 U30731 (.A1(N7790), .A2(n14559), .ZN(N43603));
    NOR2X1 U30732 (.A1(N7078), .A2(n32954), .ZN(N43604));
    INVX1 U30733 (.I(n40343), .ZN(N43605));
    NOR2X1 U30734 (.A1(N5100), .A2(n22939), .ZN(N43606));
    NOR2X1 U30735 (.A1(N2433), .A2(n42829), .ZN(N43607));
    NOR2X1 U30736 (.A1(n40079), .A2(n18165), .ZN(N43608));
    NOR2X1 U30737 (.A1(N12115), .A2(n38272), .ZN(N43609));
    INVX1 U30738 (.I(N2313), .ZN(N43610));
    NANDX1 U30739 (.A1(n26626), .A2(n17092), .ZN(N43611));
    NOR2X1 U30740 (.A1(n36745), .A2(n15135), .ZN(N43612));
    NOR2X1 U30741 (.A1(n19146), .A2(n30090), .ZN(N43613));
    INVX1 U30742 (.I(n16615), .ZN(N43614));
    NOR2X1 U30743 (.A1(n36104), .A2(n23692), .ZN(N43615));
    INVX1 U30744 (.I(n15256), .ZN(N43616));
    NOR2X1 U30745 (.A1(n28920), .A2(n20355), .ZN(N43617));
    NANDX1 U30746 (.A1(n41011), .A2(N12468), .ZN(N43618));
    NANDX1 U30747 (.A1(n38612), .A2(n42226), .ZN(N43619));
    NOR2X1 U30748 (.A1(n38908), .A2(N548), .ZN(n43620));
    NANDX1 U30749 (.A1(n31804), .A2(n36012), .ZN(N43621));
    INVX1 U30750 (.I(n14957), .ZN(N43622));
    NANDX1 U30751 (.A1(n20083), .A2(N8229), .ZN(N43623));
    NOR2X1 U30752 (.A1(N9576), .A2(n17054), .ZN(N43624));
    NANDX1 U30753 (.A1(n13476), .A2(n23348), .ZN(N43625));
    INVX1 U30754 (.I(n39259), .ZN(N43626));
    INVX1 U30755 (.I(n15728), .ZN(n43627));
    NOR2X1 U30756 (.A1(N3490), .A2(n34327), .ZN(N43628));
    NOR2X1 U30757 (.A1(n36670), .A2(n21545), .ZN(N43629));
    INVX1 U30758 (.I(n15415), .ZN(N43630));
    INVX1 U30759 (.I(n21977), .ZN(n43631));
    NOR2X1 U30760 (.A1(N1800), .A2(n22524), .ZN(N43632));
    NANDX1 U30761 (.A1(n33603), .A2(N4743), .ZN(n43633));
    NOR2X1 U30762 (.A1(n38239), .A2(n14373), .ZN(N43634));
    INVX1 U30763 (.I(n36147), .ZN(N43635));
    NOR2X1 U30764 (.A1(N12743), .A2(N9729), .ZN(N43636));
    NOR2X1 U30765 (.A1(n15898), .A2(n33076), .ZN(N43637));
    INVX1 U30766 (.I(N11684), .ZN(N43638));
    NOR2X1 U30767 (.A1(N6563), .A2(N12406), .ZN(N43639));
    NOR2X1 U30768 (.A1(n40889), .A2(n33483), .ZN(N43640));
    NANDX1 U30769 (.A1(n18962), .A2(N2914), .ZN(N43641));
    INVX1 U30770 (.I(n25326), .ZN(N43642));
    NANDX1 U30771 (.A1(N9468), .A2(n27125), .ZN(n43643));
    NOR2X1 U30772 (.A1(n26012), .A2(N6935), .ZN(N43644));
    NOR2X1 U30773 (.A1(n19416), .A2(N1701), .ZN(N43645));
    INVX1 U30774 (.I(n22582), .ZN(N43646));
    NANDX1 U30775 (.A1(N10594), .A2(n25004), .ZN(N43647));
    INVX1 U30776 (.I(n30152), .ZN(N43648));
    NANDX1 U30777 (.A1(n16539), .A2(n31307), .ZN(N43649));
    NOR2X1 U30778 (.A1(n32541), .A2(n37870), .ZN(N43650));
    NANDX1 U30779 (.A1(n41713), .A2(n24966), .ZN(N43651));
    NANDX1 U30780 (.A1(N610), .A2(n33607), .ZN(N43652));
    NOR2X1 U30781 (.A1(N8073), .A2(n15460), .ZN(N43653));
    INVX1 U30782 (.I(n17540), .ZN(N43654));
    NANDX1 U30783 (.A1(n24825), .A2(N79), .ZN(N43655));
    NOR2X1 U30784 (.A1(N12869), .A2(N9174), .ZN(N43656));
    INVX1 U30785 (.I(N4966), .ZN(N43657));
    NOR2X1 U30786 (.A1(N4313), .A2(N5239), .ZN(N43658));
    NOR2X1 U30787 (.A1(n31247), .A2(n35390), .ZN(N43659));
    NOR2X1 U30788 (.A1(n37465), .A2(n12904), .ZN(N43660));
    NANDX1 U30789 (.A1(n16214), .A2(n40453), .ZN(N43661));
    INVX1 U30790 (.I(n14454), .ZN(N43662));
    NOR2X1 U30791 (.A1(n24105), .A2(n15063), .ZN(N43663));
    NANDX1 U30792 (.A1(n17906), .A2(N12815), .ZN(N43664));
    NANDX1 U30793 (.A1(n15957), .A2(n30355), .ZN(N43665));
    INVX1 U30794 (.I(n40781), .ZN(N43666));
    NOR2X1 U30795 (.A1(n34890), .A2(n43330), .ZN(N43667));
    NANDX1 U30796 (.A1(N11675), .A2(n37975), .ZN(N43668));
    NANDX1 U30797 (.A1(n15987), .A2(n43213), .ZN(N43669));
    NANDX1 U30798 (.A1(n36914), .A2(n35130), .ZN(N43670));
    INVX1 U30799 (.I(n30906), .ZN(N43671));
    INVX1 U30800 (.I(N1670), .ZN(N43672));
    NANDX1 U30801 (.A1(n34694), .A2(n34887), .ZN(N43673));
    NOR2X1 U30802 (.A1(N2848), .A2(N5199), .ZN(N43674));
    INVX1 U30803 (.I(n37760), .ZN(n43675));
    NANDX1 U30804 (.A1(n35657), .A2(N11508), .ZN(N43676));
    NANDX1 U30805 (.A1(N12219), .A2(N7200), .ZN(N43677));
    NANDX1 U30806 (.A1(n32331), .A2(n31769), .ZN(N43678));
    NANDX1 U30807 (.A1(n18145), .A2(n33123), .ZN(N43679));
    NOR2X1 U30808 (.A1(N4754), .A2(n38790), .ZN(N43680));
    INVX1 U30809 (.I(n37802), .ZN(N43681));
    NOR2X1 U30810 (.A1(n24316), .A2(N7132), .ZN(N43682));
    NANDX1 U30811 (.A1(n18557), .A2(n41954), .ZN(N43683));
    INVX1 U30812 (.I(n42930), .ZN(N43684));
    INVX1 U30813 (.I(n20770), .ZN(N43685));
    INVX1 U30814 (.I(n28246), .ZN(N43686));
    NANDX1 U30815 (.A1(n29744), .A2(N7877), .ZN(N43687));
    NANDX1 U30816 (.A1(n30932), .A2(n26296), .ZN(N43688));
    NANDX1 U30817 (.A1(n38131), .A2(n42023), .ZN(N43689));
    INVX1 U30818 (.I(n16107), .ZN(n43690));
    NOR2X1 U30819 (.A1(n34377), .A2(N5757), .ZN(N43691));
    NOR2X1 U30820 (.A1(n39130), .A2(n34226), .ZN(N43692));
    INVX1 U30821 (.I(n33459), .ZN(N43693));
    NANDX1 U30822 (.A1(n27404), .A2(n30271), .ZN(N43694));
    INVX1 U30823 (.I(n35640), .ZN(N43695));
    INVX1 U30824 (.I(n34998), .ZN(N43696));
    INVX1 U30825 (.I(N8327), .ZN(N43697));
    NANDX1 U30826 (.A1(n16761), .A2(n36572), .ZN(N43698));
    INVX1 U30827 (.I(N3033), .ZN(N43699));
    NOR2X1 U30828 (.A1(n27589), .A2(n33964), .ZN(N43700));
    INVX1 U30829 (.I(n21810), .ZN(N43701));
    NOR2X1 U30830 (.A1(N5181), .A2(n38042), .ZN(N43702));
    NOR2X1 U30831 (.A1(n42148), .A2(n28946), .ZN(n43703));
    NOR2X1 U30832 (.A1(n35410), .A2(n14283), .ZN(N43704));
    NOR2X1 U30833 (.A1(n28178), .A2(n37422), .ZN(N43705));
    NANDX1 U30834 (.A1(N1789), .A2(n24220), .ZN(N43706));
    NOR2X1 U30835 (.A1(n37429), .A2(N9499), .ZN(N43707));
    INVX1 U30836 (.I(n18733), .ZN(N43708));
    NOR2X1 U30837 (.A1(N5296), .A2(n35494), .ZN(N43709));
    NANDX1 U30838 (.A1(N7409), .A2(n38526), .ZN(N43710));
    INVX1 U30839 (.I(n34998), .ZN(N43711));
    NOR2X1 U30840 (.A1(n41361), .A2(N3015), .ZN(N43712));
    NANDX1 U30841 (.A1(n36221), .A2(n41056), .ZN(N43713));
    INVX1 U30842 (.I(n24577), .ZN(N43714));
    INVX1 U30843 (.I(n14304), .ZN(N43715));
    NOR2X1 U30844 (.A1(n40812), .A2(n24581), .ZN(N43716));
    NANDX1 U30845 (.A1(n24441), .A2(n14370), .ZN(N43717));
    NANDX1 U30846 (.A1(N5188), .A2(n26165), .ZN(N43718));
    NOR2X1 U30847 (.A1(N4366), .A2(n19166), .ZN(N43719));
    NANDX1 U30848 (.A1(N11870), .A2(n24461), .ZN(N43720));
    NANDX1 U30849 (.A1(N12473), .A2(n31869), .ZN(N43721));
    NANDX1 U30850 (.A1(n36883), .A2(n13074), .ZN(N43722));
    INVX1 U30851 (.I(n24451), .ZN(N43723));
    NOR2X1 U30852 (.A1(n37823), .A2(n17199), .ZN(N43724));
    NOR2X1 U30853 (.A1(N11963), .A2(n31455), .ZN(N43725));
    NANDX1 U30854 (.A1(n26266), .A2(N4496), .ZN(N43726));
    NOR2X1 U30855 (.A1(N7375), .A2(n38866), .ZN(N43727));
    INVX1 U30856 (.I(N11424), .ZN(N43728));
    NANDX1 U30857 (.A1(n36207), .A2(n27268), .ZN(n43729));
    NANDX1 U30858 (.A1(n40572), .A2(N2961), .ZN(N43730));
    NOR2X1 U30859 (.A1(N8969), .A2(n27421), .ZN(N43731));
    NANDX1 U30860 (.A1(N11121), .A2(N5498), .ZN(N43732));
    NOR2X1 U30861 (.A1(n37683), .A2(n18571), .ZN(N43733));
    INVX1 U30862 (.I(n18661), .ZN(N43734));
    NOR2X1 U30863 (.A1(N10782), .A2(n25539), .ZN(N43735));
    NOR2X1 U30864 (.A1(n22744), .A2(n13522), .ZN(N43736));
    NANDX1 U30865 (.A1(n38690), .A2(N7697), .ZN(N43737));
    INVX1 U30866 (.I(n35744), .ZN(N43738));
    NOR2X1 U30867 (.A1(n18545), .A2(n36847), .ZN(N43739));
    INVX1 U30868 (.I(N11279), .ZN(N43740));
    NANDX1 U30869 (.A1(n32197), .A2(N8378), .ZN(N43741));
    NOR2X1 U30870 (.A1(n35127), .A2(N7026), .ZN(N43742));
    NOR2X1 U30871 (.A1(n35452), .A2(N7826), .ZN(N43743));
    INVX1 U30872 (.I(N7587), .ZN(N43744));
    NANDX1 U30873 (.A1(N659), .A2(n24018), .ZN(N43745));
    NANDX1 U30874 (.A1(n24997), .A2(n24480), .ZN(N43746));
    NOR2X1 U30875 (.A1(N9215), .A2(n36903), .ZN(n43747));
    NOR2X1 U30876 (.A1(n23313), .A2(n21800), .ZN(N43748));
    NOR2X1 U30877 (.A1(N518), .A2(N3751), .ZN(N43749));
    NANDX1 U30878 (.A1(n19062), .A2(n40597), .ZN(N43750));
    NOR2X1 U30879 (.A1(n30340), .A2(n17767), .ZN(N43751));
    NANDX1 U30880 (.A1(n28397), .A2(n31049), .ZN(N43752));
    INVX1 U30881 (.I(n25102), .ZN(N43753));
    NOR2X1 U30882 (.A1(N5302), .A2(n32927), .ZN(N43754));
    INVX1 U30883 (.I(n12888), .ZN(N43755));
    NANDX1 U30884 (.A1(N11025), .A2(n26585), .ZN(N43756));
    NOR2X1 U30885 (.A1(n25701), .A2(N7592), .ZN(N43757));
    NOR2X1 U30886 (.A1(n34916), .A2(N1023), .ZN(N43758));
    NANDX1 U30887 (.A1(N4436), .A2(N12502), .ZN(N43759));
    NANDX1 U30888 (.A1(N4954), .A2(n16253), .ZN(n43760));
    INVX1 U30889 (.I(n13695), .ZN(N43761));
    NOR2X1 U30890 (.A1(N12020), .A2(n33715), .ZN(n43762));
    NOR2X1 U30891 (.A1(N536), .A2(N8319), .ZN(N43763));
    NANDX1 U30892 (.A1(n13857), .A2(n33421), .ZN(n43764));
    NOR2X1 U30893 (.A1(n19158), .A2(N12555), .ZN(N43765));
    NOR2X1 U30894 (.A1(n21725), .A2(n26877), .ZN(N43766));
    NANDX1 U30895 (.A1(N4838), .A2(n18421), .ZN(N43767));
    NANDX1 U30896 (.A1(N2109), .A2(n35559), .ZN(N43768));
    NANDX1 U30897 (.A1(n36283), .A2(N4868), .ZN(N43769));
    NOR2X1 U30898 (.A1(N5313), .A2(n20987), .ZN(n43770));
    NOR2X1 U30899 (.A1(n21565), .A2(N12576), .ZN(n43771));
    INVX1 U30900 (.I(n34941), .ZN(N43772));
    NOR2X1 U30901 (.A1(n16296), .A2(N12292), .ZN(N43773));
    NANDX1 U30902 (.A1(n14295), .A2(N10370), .ZN(N43774));
    NOR2X1 U30903 (.A1(n37395), .A2(n26407), .ZN(N43775));
    NANDX1 U30904 (.A1(N6477), .A2(n42490), .ZN(n43776));
    NANDX1 U30905 (.A1(n23033), .A2(n26125), .ZN(N43777));
    NANDX1 U30906 (.A1(n41454), .A2(n25141), .ZN(N43778));
    NANDX1 U30907 (.A1(n23220), .A2(N5279), .ZN(N43779));
    NANDX1 U30908 (.A1(n28087), .A2(n23005), .ZN(N43780));
    NANDX1 U30909 (.A1(n38754), .A2(N2212), .ZN(N43781));
    INVX1 U30910 (.I(N7857), .ZN(N43782));
    NOR2X1 U30911 (.A1(n36049), .A2(n22131), .ZN(N43783));
    NANDX1 U30912 (.A1(n38020), .A2(n36941), .ZN(N43784));
    NOR2X1 U30913 (.A1(N4918), .A2(N11815), .ZN(N43785));
    NANDX1 U30914 (.A1(n21004), .A2(n38998), .ZN(N43786));
    INVX1 U30915 (.I(n20022), .ZN(N43787));
    NOR2X1 U30916 (.A1(N7854), .A2(n35826), .ZN(N43788));
    NANDX1 U30917 (.A1(N5835), .A2(N7174), .ZN(N43789));
    INVX1 U30918 (.I(n29055), .ZN(N43790));
    INVX1 U30919 (.I(N41), .ZN(N43791));
    INVX1 U30920 (.I(n25137), .ZN(N43792));
    INVX1 U30921 (.I(n31782), .ZN(N43793));
    INVX1 U30922 (.I(n34485), .ZN(N43794));
    INVX1 U30923 (.I(n34974), .ZN(N43795));
    INVX1 U30924 (.I(n18297), .ZN(n43796));
    NANDX1 U30925 (.A1(N11289), .A2(N1445), .ZN(N43797));
    NANDX1 U30926 (.A1(N5886), .A2(N2939), .ZN(N43798));
    NOR2X1 U30927 (.A1(n26889), .A2(n31616), .ZN(N43799));
    INVX1 U30928 (.I(n36590), .ZN(N43800));
    NOR2X1 U30929 (.A1(n24656), .A2(n18624), .ZN(N43801));
    INVX1 U30930 (.I(n30490), .ZN(N43802));
    NANDX1 U30931 (.A1(N7700), .A2(N5752), .ZN(n43803));
    NOR2X1 U30932 (.A1(N7740), .A2(n42253), .ZN(N43804));
    NOR2X1 U30933 (.A1(n41116), .A2(n30562), .ZN(N43805));
    INVX1 U30934 (.I(n32128), .ZN(N43806));
    NANDX1 U30935 (.A1(n20315), .A2(N5397), .ZN(N43807));
    NANDX1 U30936 (.A1(n25416), .A2(n16685), .ZN(N43808));
    NANDX1 U30937 (.A1(n35580), .A2(n22570), .ZN(N43809));
    NOR2X1 U30938 (.A1(n24089), .A2(n39138), .ZN(N43810));
    NANDX1 U30939 (.A1(n30570), .A2(n32256), .ZN(N43811));
    INVX1 U30940 (.I(N11753), .ZN(N43812));
    NANDX1 U30941 (.A1(N418), .A2(n31923), .ZN(N43813));
    INVX1 U30942 (.I(n41269), .ZN(N43814));
    NOR2X1 U30943 (.A1(n30172), .A2(N5537), .ZN(N43815));
    NOR2X1 U30944 (.A1(n19125), .A2(n36332), .ZN(N43816));
    INVX1 U30945 (.I(N4466), .ZN(N43817));
    NOR2X1 U30946 (.A1(n19311), .A2(n24780), .ZN(N43818));
    NOR2X1 U30947 (.A1(N222), .A2(N6723), .ZN(N43819));
    INVX1 U30948 (.I(n15729), .ZN(N43820));
    NOR2X1 U30949 (.A1(n38677), .A2(n23854), .ZN(N43821));
    NANDX1 U30950 (.A1(n34342), .A2(n20122), .ZN(N43822));
    INVX1 U30951 (.I(N12805), .ZN(N43823));
    INVX1 U30952 (.I(N1129), .ZN(N43824));
    NANDX1 U30953 (.A1(n18425), .A2(n33051), .ZN(N43825));
    NOR2X1 U30954 (.A1(n16221), .A2(n16932), .ZN(N43826));
    NANDX1 U30955 (.A1(n21757), .A2(n32746), .ZN(N43827));
    NANDX1 U30956 (.A1(n14617), .A2(n25329), .ZN(N43828));
    INVX1 U30957 (.I(n29284), .ZN(N43829));
    NOR2X1 U30958 (.A1(N3729), .A2(n39027), .ZN(N43830));
    NOR2X1 U30959 (.A1(N10451), .A2(N11662), .ZN(N43831));
    NANDX1 U30960 (.A1(n32113), .A2(N6866), .ZN(N43832));
    NOR2X1 U30961 (.A1(n34391), .A2(n41207), .ZN(N43833));
    NANDX1 U30962 (.A1(n13447), .A2(N10540), .ZN(N43834));
    NOR2X1 U30963 (.A1(N4255), .A2(n20430), .ZN(N43835));
    NANDX1 U30964 (.A1(n26985), .A2(n42883), .ZN(N43836));
    NANDX1 U30965 (.A1(n33596), .A2(N8563), .ZN(N43837));
    NOR2X1 U30966 (.A1(n22869), .A2(n26519), .ZN(N43838));
    INVX1 U30967 (.I(N4725), .ZN(N43839));
    INVX1 U30968 (.I(n40853), .ZN(N43840));
    NANDX1 U30969 (.A1(n42348), .A2(n36407), .ZN(N43841));
    INVX1 U30970 (.I(n42479), .ZN(N43842));
    NOR2X1 U30971 (.A1(n16265), .A2(n31119), .ZN(N43843));
    NANDX1 U30972 (.A1(n36593), .A2(N11718), .ZN(n43844));
    NANDX1 U30973 (.A1(n33571), .A2(n25164), .ZN(N43845));
    NANDX1 U30974 (.A1(N5083), .A2(n19098), .ZN(N43846));
    NANDX1 U30975 (.A1(n28172), .A2(N2610), .ZN(N43847));
    INVX1 U30976 (.I(n34329), .ZN(N43848));
    NOR2X1 U30977 (.A1(n17177), .A2(n41602), .ZN(N43849));
    INVX1 U30978 (.I(n33376), .ZN(N43850));
    NANDX1 U30979 (.A1(N10006), .A2(n28523), .ZN(N43851));
    NANDX1 U30980 (.A1(n38729), .A2(n27399), .ZN(N43852));
    NOR2X1 U30981 (.A1(n25366), .A2(n26405), .ZN(N43853));
    NOR2X1 U30982 (.A1(n41631), .A2(n14051), .ZN(N43854));
    NANDX1 U30983 (.A1(n24431), .A2(n15448), .ZN(N43855));
    NOR2X1 U30984 (.A1(N4209), .A2(n30291), .ZN(N43856));
    NANDX1 U30985 (.A1(n42444), .A2(N5916), .ZN(N43857));
    NOR2X1 U30986 (.A1(n27143), .A2(N8525), .ZN(n43858));
    INVX1 U30987 (.I(N7679), .ZN(N43859));
    INVX1 U30988 (.I(N7754), .ZN(N43860));
    INVX1 U30989 (.I(N6539), .ZN(N43861));
    INVX1 U30990 (.I(n25827), .ZN(N43862));
    NANDX1 U30991 (.A1(n15859), .A2(n43227), .ZN(N43863));
    INVX1 U30992 (.I(n43257), .ZN(N43864));
    INVX1 U30993 (.I(n16526), .ZN(N43865));
    INVX1 U30994 (.I(n27210), .ZN(N43866));
    NANDX1 U30995 (.A1(n29920), .A2(n22640), .ZN(N43867));
    NOR2X1 U30996 (.A1(n35047), .A2(N6625), .ZN(N43868));
    NOR2X1 U30997 (.A1(n21866), .A2(n33176), .ZN(N43869));
    NOR2X1 U30998 (.A1(n17461), .A2(n25459), .ZN(N43870));
    NOR2X1 U30999 (.A1(n25986), .A2(n26355), .ZN(N43871));
    NOR2X1 U31000 (.A1(n16923), .A2(n23788), .ZN(N43872));
    NOR2X1 U31001 (.A1(n13141), .A2(n21444), .ZN(N43873));
    NOR2X1 U31002 (.A1(N9044), .A2(n37303), .ZN(N43874));
    INVX1 U31003 (.I(N10524), .ZN(N43875));
    NANDX1 U31004 (.A1(n13198), .A2(n27049), .ZN(N43876));
    INVX1 U31005 (.I(n40407), .ZN(N43877));
    NOR2X1 U31006 (.A1(n29083), .A2(N9255), .ZN(n43878));
    NANDX1 U31007 (.A1(n20657), .A2(n15879), .ZN(N43879));
    NANDX1 U31008 (.A1(n32202), .A2(n38735), .ZN(N43880));
    NANDX1 U31009 (.A1(N6191), .A2(N10401), .ZN(N43881));
    INVX1 U31010 (.I(n21856), .ZN(N43882));
    NANDX1 U31011 (.A1(n15280), .A2(n28458), .ZN(N43883));
    NOR2X1 U31012 (.A1(n34089), .A2(n31278), .ZN(N43884));
    INVX1 U31013 (.I(n14612), .ZN(N43885));
    NOR2X1 U31014 (.A1(N11704), .A2(n38361), .ZN(N43886));
    NANDX1 U31015 (.A1(n28151), .A2(N8086), .ZN(N43887));
    NOR2X1 U31016 (.A1(n27314), .A2(n38172), .ZN(N43888));
    NANDX1 U31017 (.A1(N2604), .A2(N3954), .ZN(N43889));
    NANDX1 U31018 (.A1(n12940), .A2(N9513), .ZN(n43890));
    INVX1 U31019 (.I(N1670), .ZN(N43891));
    INVX1 U31020 (.I(n23862), .ZN(N43892));
    NOR2X1 U31021 (.A1(N4855), .A2(n26140), .ZN(N43893));
    NOR2X1 U31022 (.A1(n31289), .A2(n41420), .ZN(N43894));
    NANDX1 U31023 (.A1(n38039), .A2(n21716), .ZN(N43895));
    NOR2X1 U31024 (.A1(N12441), .A2(n36327), .ZN(N43896));
    NANDX1 U31025 (.A1(n13824), .A2(n20895), .ZN(N43897));
    NANDX1 U31026 (.A1(n41974), .A2(n28980), .ZN(N43898));
    INVX1 U31027 (.I(n15495), .ZN(n43899));
    NANDX1 U31028 (.A1(N1583), .A2(n18098), .ZN(N43900));
    INVX1 U31029 (.I(n32546), .ZN(N43901));
    NANDX1 U31030 (.A1(n16505), .A2(N5659), .ZN(N43902));
    NOR2X1 U31031 (.A1(N10959), .A2(n19200), .ZN(N43903));
    NANDX1 U31032 (.A1(n15813), .A2(N1868), .ZN(N43904));
    NANDX1 U31033 (.A1(N3629), .A2(n32967), .ZN(N43905));
    INVX1 U31034 (.I(n31348), .ZN(N43906));
    NANDX1 U31035 (.A1(N4923), .A2(N316), .ZN(N43907));
    NANDX1 U31036 (.A1(n16787), .A2(N3819), .ZN(N43908));
    NANDX1 U31037 (.A1(n36023), .A2(n35473), .ZN(N43909));
    NOR2X1 U31038 (.A1(n35887), .A2(N7495), .ZN(N43910));
    INVX1 U31039 (.I(n27149), .ZN(N43911));
    NANDX1 U31040 (.A1(N10175), .A2(n16222), .ZN(N43912));
    NOR2X1 U31041 (.A1(n16359), .A2(N11560), .ZN(N43913));
    NOR2X1 U31042 (.A1(n27317), .A2(n30760), .ZN(N43914));
    NANDX1 U31043 (.A1(n43129), .A2(n32627), .ZN(N43915));
    INVX1 U31044 (.I(n36438), .ZN(N43916));
    INVX1 U31045 (.I(n20582), .ZN(N43917));
    NOR2X1 U31046 (.A1(N12690), .A2(n15184), .ZN(N43918));
    NANDX1 U31047 (.A1(n29265), .A2(n31970), .ZN(N43919));
    INVX1 U31048 (.I(n33582), .ZN(n43920));
    NANDX1 U31049 (.A1(n43278), .A2(n13086), .ZN(N43921));
    NOR2X1 U31050 (.A1(N7301), .A2(n39100), .ZN(N43922));
    NOR2X1 U31051 (.A1(n22573), .A2(n38955), .ZN(N43923));
    NANDX1 U31052 (.A1(n35730), .A2(N11841), .ZN(N43924));
    NOR2X1 U31053 (.A1(n27801), .A2(n39158), .ZN(N43925));
    NANDX1 U31054 (.A1(n29477), .A2(n38814), .ZN(N43926));
    INVX1 U31055 (.I(n27000), .ZN(N43927));
    NOR2X1 U31056 (.A1(N8504), .A2(N4109), .ZN(N43928));
    NOR2X1 U31057 (.A1(n21193), .A2(n19292), .ZN(N43929));
    INVX1 U31058 (.I(N6985), .ZN(N43930));
    NOR2X1 U31059 (.A1(n24412), .A2(n30246), .ZN(N43931));
    NANDX1 U31060 (.A1(n24217), .A2(n43331), .ZN(N43932));
    INVX1 U31061 (.I(n21197), .ZN(n43933));
    NANDX1 U31062 (.A1(N8573), .A2(N297), .ZN(N43934));
    NANDX1 U31063 (.A1(n37916), .A2(n25706), .ZN(N43935));
    NANDX1 U31064 (.A1(n35347), .A2(n43186), .ZN(N43936));
    NANDX1 U31065 (.A1(N9744), .A2(n29190), .ZN(N43937));
    NANDX1 U31066 (.A1(n16768), .A2(N12717), .ZN(N43938));
    NANDX1 U31067 (.A1(n25271), .A2(n16825), .ZN(N43939));
    NANDX1 U31068 (.A1(n36144), .A2(n25796), .ZN(n43940));
    NOR2X1 U31069 (.A1(n32808), .A2(n23265), .ZN(n43941));
    NOR2X1 U31070 (.A1(n19582), .A2(N1781), .ZN(N43942));
    NOR2X1 U31071 (.A1(N9120), .A2(n30384), .ZN(N43943));
    INVX1 U31072 (.I(n37758), .ZN(N43944));
    INVX1 U31073 (.I(N9247), .ZN(N43945));
    NANDX1 U31074 (.A1(n23080), .A2(n34952), .ZN(N43946));
    INVX1 U31075 (.I(N4634), .ZN(N43947));
    NOR2X1 U31076 (.A1(n42540), .A2(n14377), .ZN(N43948));
    INVX1 U31077 (.I(n15735), .ZN(N43949));
    NANDX1 U31078 (.A1(n33100), .A2(N10389), .ZN(N43950));
    NOR2X1 U31079 (.A1(n39604), .A2(n17661), .ZN(N43951));
    NANDX1 U31080 (.A1(N11608), .A2(n20898), .ZN(N43952));
    NOR2X1 U31081 (.A1(n34872), .A2(N5075), .ZN(N43953));
    INVX1 U31082 (.I(n36652), .ZN(n43954));
    INVX1 U31083 (.I(n36162), .ZN(N43955));
    INVX1 U31084 (.I(n22417), .ZN(N43956));
    NANDX1 U31085 (.A1(n41879), .A2(n21343), .ZN(N43957));
    NANDX1 U31086 (.A1(N11166), .A2(N12823), .ZN(N43958));
    NOR2X1 U31087 (.A1(N5479), .A2(n37168), .ZN(N43959));
    NANDX1 U31088 (.A1(n19855), .A2(n14078), .ZN(N43960));
    NOR2X1 U31089 (.A1(n40679), .A2(n36857), .ZN(N43961));
    INVX1 U31090 (.I(n32981), .ZN(N43962));
    NOR2X1 U31091 (.A1(N7525), .A2(n17954), .ZN(n43963));
    NANDX1 U31092 (.A1(n18102), .A2(n25414), .ZN(N43964));
    INVX1 U31093 (.I(n23176), .ZN(N43965));
    NOR2X1 U31094 (.A1(n18854), .A2(n26323), .ZN(N43966));
    INVX1 U31095 (.I(n21777), .ZN(N43967));
    INVX1 U31096 (.I(N1159), .ZN(N43968));
    NANDX1 U31097 (.A1(N5970), .A2(n29371), .ZN(N43969));
    INVX1 U31098 (.I(n18792), .ZN(N43970));
    NOR2X1 U31099 (.A1(n26506), .A2(N12487), .ZN(N43971));
    NANDX1 U31100 (.A1(n36040), .A2(n16245), .ZN(N43972));
    NANDX1 U31101 (.A1(n22926), .A2(N9629), .ZN(N43973));
    NANDX1 U31102 (.A1(N12434), .A2(n21977), .ZN(N43974));
    INVX1 U31103 (.I(n20067), .ZN(N43975));
    NOR2X1 U31104 (.A1(n16864), .A2(N2009), .ZN(N43976));
    NOR2X1 U31105 (.A1(n40040), .A2(N672), .ZN(N43977));
    NANDX1 U31106 (.A1(N12570), .A2(n25176), .ZN(N43978));
    INVX1 U31107 (.I(n40669), .ZN(N43979));
    NANDX1 U31108 (.A1(n24834), .A2(N3167), .ZN(N43980));
    NOR2X1 U31109 (.A1(N2389), .A2(N11638), .ZN(N43981));
    NANDX1 U31110 (.A1(n18574), .A2(n24125), .ZN(N43982));
    INVX1 U31111 (.I(N821), .ZN(N43983));
    NOR2X1 U31112 (.A1(n17037), .A2(n23747), .ZN(N43984));
    NANDX1 U31113 (.A1(N8275), .A2(n25860), .ZN(N43985));
    INVX1 U31114 (.I(N7037), .ZN(N43986));
    NOR2X1 U31115 (.A1(n20641), .A2(n23901), .ZN(N43987));
    NANDX1 U31116 (.A1(N5303), .A2(N10148), .ZN(N43988));
    NOR2X1 U31117 (.A1(N8818), .A2(N12397), .ZN(N43989));
    NANDX1 U31118 (.A1(n23789), .A2(N9594), .ZN(N43990));
    NOR2X1 U31119 (.A1(N5150), .A2(N2440), .ZN(N43991));
    NOR2X1 U31120 (.A1(n40690), .A2(n14077), .ZN(N43992));
    NOR2X1 U31121 (.A1(N5471), .A2(n27881), .ZN(n43993));
    NOR2X1 U31122 (.A1(N6291), .A2(n14457), .ZN(N43994));
    NOR2X1 U31123 (.A1(n19717), .A2(N342), .ZN(N43995));
    NOR2X1 U31124 (.A1(N2105), .A2(N8203), .ZN(N43996));
    INVX1 U31125 (.I(N4559), .ZN(N43997));
    NANDX1 U31126 (.A1(n18837), .A2(n42173), .ZN(n43998));
    NANDX1 U31127 (.A1(n18664), .A2(n26666), .ZN(N43999));
    INVX1 U31128 (.I(n31060), .ZN(N44000));
    NOR2X1 U31129 (.A1(n35790), .A2(n40653), .ZN(N44001));
    NOR2X1 U31130 (.A1(n30619), .A2(n43092), .ZN(N44002));
    NOR2X1 U31131 (.A1(n17516), .A2(N3377), .ZN(N44003));
    NANDX1 U31132 (.A1(n22986), .A2(n31257), .ZN(N44004));
    NANDX1 U31133 (.A1(n18957), .A2(N2242), .ZN(N44005));
    INVX1 U31134 (.I(n28353), .ZN(n44006));
    INVX1 U31135 (.I(n16056), .ZN(N44007));
    NANDX1 U31136 (.A1(n33617), .A2(N10992), .ZN(N44008));
    NOR2X1 U31137 (.A1(N8667), .A2(n29828), .ZN(N44009));
    NANDX1 U31138 (.A1(n22172), .A2(N5019), .ZN(N44010));
    NOR2X1 U31139 (.A1(n34173), .A2(n25758), .ZN(N44011));
    NOR2X1 U31140 (.A1(n16171), .A2(N12619), .ZN(N44012));
    NOR2X1 U31141 (.A1(N3317), .A2(N1918), .ZN(N44013));
    NOR2X1 U31142 (.A1(n20833), .A2(N5294), .ZN(N44014));
    NANDX1 U31143 (.A1(n33498), .A2(n36551), .ZN(N44015));
    NOR2X1 U31144 (.A1(n42134), .A2(n28472), .ZN(N44016));
    NANDX1 U31145 (.A1(n27015), .A2(n20734), .ZN(N44017));
    NOR2X1 U31146 (.A1(N3679), .A2(N10878), .ZN(N44018));
    NOR2X1 U31147 (.A1(n28374), .A2(N9224), .ZN(N44019));
    INVX1 U31148 (.I(n41448), .ZN(N44020));
    INVX1 U31149 (.I(n40327), .ZN(N44021));
    INVX1 U31150 (.I(N11776), .ZN(N44022));
    NANDX1 U31151 (.A1(n16524), .A2(n27946), .ZN(N44023));
    NOR2X1 U31152 (.A1(n34515), .A2(n20942), .ZN(N44024));
    NANDX1 U31153 (.A1(n42658), .A2(n41774), .ZN(N44025));
    NANDX1 U31154 (.A1(n29159), .A2(n21480), .ZN(N44026));
    NOR2X1 U31155 (.A1(N79), .A2(N9821), .ZN(N44027));
    INVX1 U31156 (.I(n42626), .ZN(N44028));
    NANDX1 U31157 (.A1(n20611), .A2(N3964), .ZN(N44029));
    INVX1 U31158 (.I(n21168), .ZN(N44030));
    NANDX1 U31159 (.A1(n15095), .A2(n30392), .ZN(N44031));
    NOR2X1 U31160 (.A1(N2750), .A2(N7994), .ZN(N44032));
    INVX1 U31161 (.I(n30145), .ZN(N44033));
    NOR2X1 U31162 (.A1(N10426), .A2(n36349), .ZN(N44034));
    INVX1 U31163 (.I(n35336), .ZN(N44035));
    NANDX1 U31164 (.A1(n14864), .A2(n18691), .ZN(N44036));
    NOR2X1 U31165 (.A1(N2845), .A2(N7339), .ZN(N44037));
    NOR2X1 U31166 (.A1(n24324), .A2(n32538), .ZN(N44038));
    INVX1 U31167 (.I(n23825), .ZN(N44039));
    NANDX1 U31168 (.A1(n34326), .A2(N6867), .ZN(N44040));
    NOR2X1 U31169 (.A1(n27969), .A2(n37060), .ZN(N44041));
    NOR2X1 U31170 (.A1(n37413), .A2(n41834), .ZN(N44042));
    NANDX1 U31171 (.A1(n38693), .A2(n34264), .ZN(N44043));
    NANDX1 U31172 (.A1(n36827), .A2(n20936), .ZN(N44044));
    NANDX1 U31173 (.A1(N3781), .A2(N3492), .ZN(N44045));
    NOR2X1 U31174 (.A1(n28796), .A2(n20563), .ZN(N44046));
    INVX1 U31175 (.I(N4014), .ZN(N44047));
    NOR2X1 U31176 (.A1(n26071), .A2(N11352), .ZN(N44048));
    NANDX1 U31177 (.A1(n40075), .A2(n33569), .ZN(N44049));
    INVX1 U31178 (.I(n20427), .ZN(N44050));
    NOR2X1 U31179 (.A1(N10995), .A2(n27293), .ZN(N44051));
    NOR2X1 U31180 (.A1(n28644), .A2(n20881), .ZN(N44052));
    NANDX1 U31181 (.A1(n22584), .A2(N8922), .ZN(N44053));
    NANDX1 U31182 (.A1(N7485), .A2(n43185), .ZN(n44054));
    NOR2X1 U31183 (.A1(N839), .A2(N10329), .ZN(N44055));
    INVX1 U31184 (.I(n37771), .ZN(N44056));
    NOR2X1 U31185 (.A1(n25662), .A2(n23094), .ZN(N44057));
    NOR2X1 U31186 (.A1(N5416), .A2(n27107), .ZN(N44058));
    NOR2X1 U31187 (.A1(n31487), .A2(n28139), .ZN(N44059));
    NOR2X1 U31188 (.A1(n17769), .A2(n18235), .ZN(N44060));
    NOR2X1 U31189 (.A1(n38195), .A2(n20106), .ZN(N44061));
    NANDX1 U31190 (.A1(N11695), .A2(n21210), .ZN(N44062));
    NOR2X1 U31191 (.A1(n22255), .A2(n42715), .ZN(N44063));
    INVX1 U31192 (.I(n31177), .ZN(N44064));
    NANDX1 U31193 (.A1(n28111), .A2(n30889), .ZN(N44065));
    NANDX1 U31194 (.A1(n28949), .A2(n41217), .ZN(N44066));
    NOR2X1 U31195 (.A1(n12928), .A2(N1245), .ZN(N44067));
    INVX1 U31196 (.I(n36021), .ZN(n44068));
    NOR2X1 U31197 (.A1(N4867), .A2(N9336), .ZN(N44069));
    NOR2X1 U31198 (.A1(n26033), .A2(n37474), .ZN(N44070));
    NANDX1 U31199 (.A1(N329), .A2(N1916), .ZN(N44071));
    NANDX1 U31200 (.A1(n38523), .A2(n22022), .ZN(N44072));
    INVX1 U31201 (.I(n39898), .ZN(N44073));
    NOR2X1 U31202 (.A1(N12217), .A2(n18680), .ZN(N44074));
    INVX1 U31203 (.I(n32843), .ZN(N44075));
    NOR2X1 U31204 (.A1(n29259), .A2(n17481), .ZN(N44076));
    INVX1 U31205 (.I(n39542), .ZN(N44077));
    INVX1 U31206 (.I(n14377), .ZN(N44078));
    NANDX1 U31207 (.A1(N5564), .A2(n15621), .ZN(N44079));
    NANDX1 U31208 (.A1(n31265), .A2(n30607), .ZN(N44080));
    INVX1 U31209 (.I(n40600), .ZN(N44081));
    NANDX1 U31210 (.A1(N210), .A2(n24281), .ZN(N44082));
    NOR2X1 U31211 (.A1(N538), .A2(n15876), .ZN(N44083));
    NANDX1 U31212 (.A1(n28741), .A2(n37897), .ZN(N44084));
    NANDX1 U31213 (.A1(n25166), .A2(n27336), .ZN(N44085));
    NANDX1 U31214 (.A1(N373), .A2(n16016), .ZN(N44086));
    NANDX1 U31215 (.A1(N6757), .A2(N1803), .ZN(N44087));
    NOR2X1 U31216 (.A1(n23389), .A2(n31024), .ZN(N44088));
    INVX1 U31217 (.I(n37765), .ZN(N44089));
    INVX1 U31218 (.I(N2286), .ZN(N44090));
    INVX1 U31219 (.I(N3345), .ZN(N44091));
    NOR2X1 U31220 (.A1(n30200), .A2(n20994), .ZN(N44092));
    INVX1 U31221 (.I(n16575), .ZN(N44093));
    NANDX1 U31222 (.A1(n34317), .A2(n37719), .ZN(N44094));
    NOR2X1 U31223 (.A1(N6721), .A2(n39525), .ZN(N44095));
    INVX1 U31224 (.I(n34297), .ZN(n44096));
    NOR2X1 U31225 (.A1(n21853), .A2(n18160), .ZN(N44097));
    NOR2X1 U31226 (.A1(N11906), .A2(n34176), .ZN(N44098));
    NANDX1 U31227 (.A1(N8342), .A2(n25658), .ZN(N44099));
    NANDX1 U31228 (.A1(n31730), .A2(N2889), .ZN(N44100));
    NOR2X1 U31229 (.A1(n26022), .A2(n36924), .ZN(N44101));
    INVX1 U31230 (.I(n25615), .ZN(N44102));
    INVX1 U31231 (.I(n42836), .ZN(N44103));
    INVX1 U31232 (.I(n17789), .ZN(n44104));
    NANDX1 U31233 (.A1(n18596), .A2(n38991), .ZN(N44105));
    NOR2X1 U31234 (.A1(N12842), .A2(N6939), .ZN(N44106));
    NOR2X1 U31235 (.A1(N8894), .A2(N3626), .ZN(N44107));
    NANDX1 U31236 (.A1(N286), .A2(n15159), .ZN(N44108));
    NANDX1 U31237 (.A1(n42705), .A2(n27064), .ZN(N44109));
    NOR2X1 U31238 (.A1(N5425), .A2(n35405), .ZN(N44110));
    NANDX1 U31239 (.A1(n15703), .A2(n23662), .ZN(N44111));
    NANDX1 U31240 (.A1(n33023), .A2(n39363), .ZN(N44112));
    INVX1 U31241 (.I(n42309), .ZN(N44113));
    NOR2X1 U31242 (.A1(n37956), .A2(n41672), .ZN(N44114));
    INVX1 U31243 (.I(N1952), .ZN(N44115));
    NANDX1 U31244 (.A1(n42123), .A2(n40943), .ZN(N44116));
    NANDX1 U31245 (.A1(N1172), .A2(n37561), .ZN(N44117));
    INVX1 U31246 (.I(n43218), .ZN(N44118));
    NANDX1 U31247 (.A1(N2276), .A2(N31), .ZN(N44119));
    NOR2X1 U31248 (.A1(n18224), .A2(n42735), .ZN(n44120));
    INVX1 U31249 (.I(N4235), .ZN(N44121));
    NANDX1 U31250 (.A1(N11227), .A2(n15903), .ZN(N44122));
    NOR2X1 U31251 (.A1(n24568), .A2(n20139), .ZN(N44123));
    NOR2X1 U31252 (.A1(n20459), .A2(n17827), .ZN(N44124));
    INVX1 U31253 (.I(n31644), .ZN(N44125));
    INVX1 U31254 (.I(n29807), .ZN(N44126));
    INVX1 U31255 (.I(n14261), .ZN(N44127));
    NOR2X1 U31256 (.A1(N28), .A2(N1411), .ZN(N44128));
    INVX1 U31257 (.I(N1200), .ZN(N44129));
    INVX1 U31258 (.I(n39415), .ZN(N44130));
    NANDX1 U31259 (.A1(n16045), .A2(n41690), .ZN(N44131));
    NANDX1 U31260 (.A1(N8276), .A2(N6121), .ZN(N44132));
    NANDX1 U31261 (.A1(n27571), .A2(N10355), .ZN(N44133));
    NOR2X1 U31262 (.A1(n28477), .A2(n15937), .ZN(n44134));
    NANDX1 U31263 (.A1(N9573), .A2(n36075), .ZN(N44135));
    NANDX1 U31264 (.A1(n19711), .A2(N10429), .ZN(N44136));
    NOR2X1 U31265 (.A1(N7882), .A2(n22738), .ZN(N44137));
    INVX1 U31266 (.I(N9259), .ZN(n44138));
    INVX1 U31267 (.I(n41191), .ZN(N44139));
    NANDX1 U31268 (.A1(n17769), .A2(n32646), .ZN(n44140));
    NANDX1 U31269 (.A1(N2948), .A2(n28588), .ZN(N44141));
    INVX1 U31270 (.I(n18992), .ZN(N44142));
    NANDX1 U31271 (.A1(n24916), .A2(n27267), .ZN(N44143));
    NOR2X1 U31272 (.A1(N4512), .A2(N1045), .ZN(N44144));
    NANDX1 U31273 (.A1(N11626), .A2(n29522), .ZN(N44145));
    NANDX1 U31274 (.A1(n28810), .A2(n39094), .ZN(N44146));
    NOR2X1 U31275 (.A1(n35293), .A2(n15332), .ZN(N44147));
    NANDX1 U31276 (.A1(n29911), .A2(n12893), .ZN(N44148));
    NOR2X1 U31277 (.A1(N544), .A2(n22151), .ZN(N44149));
    INVX1 U31278 (.I(n41734), .ZN(N44150));
    INVX1 U31279 (.I(N1206), .ZN(N44151));
    INVX1 U31280 (.I(N10962), .ZN(N44152));
    NOR2X1 U31281 (.A1(n38855), .A2(N1751), .ZN(N44153));
    NOR2X1 U31282 (.A1(N11868), .A2(n16346), .ZN(N44154));
    NOR2X1 U31283 (.A1(n34472), .A2(n20857), .ZN(N44155));
    NOR2X1 U31284 (.A1(n13639), .A2(n22163), .ZN(N44156));
    INVX1 U31285 (.I(N8741), .ZN(n44157));
    INVX1 U31286 (.I(n35317), .ZN(N44158));
    NANDX1 U31287 (.A1(n42792), .A2(n40328), .ZN(N44159));
    INVX1 U31288 (.I(n29230), .ZN(N44160));
    INVX1 U31289 (.I(n27963), .ZN(N44161));
    INVX1 U31290 (.I(n21579), .ZN(N44162));
    INVX1 U31291 (.I(N7395), .ZN(N44163));
    NANDX1 U31292 (.A1(N2285), .A2(n27982), .ZN(N44164));
    NANDX1 U31293 (.A1(n39590), .A2(n13045), .ZN(N44165));
    INVX1 U31294 (.I(n42093), .ZN(N44166));
    INVX1 U31295 (.I(n17961), .ZN(N44167));
    NANDX1 U31296 (.A1(n38743), .A2(n28497), .ZN(N44168));
    NANDX1 U31297 (.A1(N8909), .A2(N7187), .ZN(N44169));
    NANDX1 U31298 (.A1(N7330), .A2(N4366), .ZN(n44170));
    NOR2X1 U31299 (.A1(n26607), .A2(N3685), .ZN(N44171));
    NOR2X1 U31300 (.A1(N546), .A2(n32915), .ZN(N44172));
    INVX1 U31301 (.I(n28508), .ZN(n44173));
    INVX1 U31302 (.I(N1023), .ZN(N44174));
    NOR2X1 U31303 (.A1(N5970), .A2(n33397), .ZN(N44175));
    NANDX1 U31304 (.A1(n23632), .A2(n33261), .ZN(n44176));
    NOR2X1 U31305 (.A1(n36676), .A2(n24556), .ZN(N44177));
    INVX1 U31306 (.I(N7795), .ZN(N44178));
    NANDX1 U31307 (.A1(n34360), .A2(n36217), .ZN(n44179));
    NOR2X1 U31308 (.A1(n29453), .A2(N1654), .ZN(n44180));
    NOR2X1 U31309 (.A1(n20769), .A2(n42135), .ZN(N44181));
    NANDX1 U31310 (.A1(N3930), .A2(n14949), .ZN(N44182));
    NOR2X1 U31311 (.A1(n27419), .A2(n15495), .ZN(N44183));
    NOR2X1 U31312 (.A1(N6863), .A2(n33682), .ZN(N44184));
    NOR2X1 U31313 (.A1(N7885), .A2(n19797), .ZN(N44185));
    INVX1 U31314 (.I(n41281), .ZN(N44186));
    INVX1 U31315 (.I(n19114), .ZN(N44187));
    NOR2X1 U31316 (.A1(N5224), .A2(N1997), .ZN(N44188));
    NANDX1 U31317 (.A1(N11192), .A2(n42943), .ZN(N44189));
    INVX1 U31318 (.I(n35231), .ZN(N44190));
    NANDX1 U31319 (.A1(N7775), .A2(N10891), .ZN(N44191));
    INVX1 U31320 (.I(n21861), .ZN(N44192));
    NOR2X1 U31321 (.A1(n15363), .A2(n29993), .ZN(N44193));
    NOR2X1 U31322 (.A1(n30311), .A2(N8657), .ZN(N44194));
    NANDX1 U31323 (.A1(N2333), .A2(n43067), .ZN(N44195));
    NOR2X1 U31324 (.A1(n36015), .A2(n32580), .ZN(N44196));
    INVX1 U31325 (.I(N2019), .ZN(N44197));
    INVX1 U31326 (.I(N1130), .ZN(N44198));
    INVX1 U31327 (.I(N3704), .ZN(N44199));
    NANDX1 U31328 (.A1(n38269), .A2(n38852), .ZN(N44200));
    NOR2X1 U31329 (.A1(n39140), .A2(n38323), .ZN(N44201));
    NOR2X1 U31330 (.A1(n30899), .A2(n30538), .ZN(N44202));
    NOR2X1 U31331 (.A1(n41789), .A2(N3766), .ZN(N44203));
    NOR2X1 U31332 (.A1(n19656), .A2(n19128), .ZN(N44204));
    INVX1 U31333 (.I(N1453), .ZN(N44205));
    NOR2X1 U31334 (.A1(n18437), .A2(N347), .ZN(N44206));
    NOR2X1 U31335 (.A1(N7711), .A2(n39256), .ZN(N44207));
    NOR2X1 U31336 (.A1(n40290), .A2(N9424), .ZN(N44208));
    NANDX1 U31337 (.A1(n24879), .A2(N233), .ZN(N44209));
    NOR2X1 U31338 (.A1(n18262), .A2(n22111), .ZN(N44210));
    NOR2X1 U31339 (.A1(n13642), .A2(N2349), .ZN(n44211));
    NOR2X1 U31340 (.A1(N8492), .A2(N6294), .ZN(N44212));
    INVX1 U31341 (.I(n28709), .ZN(N44213));
    INVX1 U31342 (.I(n14302), .ZN(n44214));
    NOR2X1 U31343 (.A1(n30954), .A2(n23637), .ZN(N44215));
    INVX1 U31344 (.I(n40734), .ZN(N44216));
    INVX1 U31345 (.I(N3774), .ZN(N44217));
    NANDX1 U31346 (.A1(n15116), .A2(N1752), .ZN(N44218));
    NOR2X1 U31347 (.A1(N10899), .A2(n25424), .ZN(N44219));
    INVX1 U31348 (.I(N10002), .ZN(N44220));
    INVX1 U31349 (.I(n34783), .ZN(N44221));
    INVX1 U31350 (.I(n33225), .ZN(N44222));
    NANDX1 U31351 (.A1(n22025), .A2(n32964), .ZN(n44223));
    INVX1 U31352 (.I(n14054), .ZN(N44224));
    NOR2X1 U31353 (.A1(N11065), .A2(n20347), .ZN(N44225));
    INVX1 U31354 (.I(n29453), .ZN(N44226));
    NOR2X1 U31355 (.A1(N4864), .A2(N8134), .ZN(N44227));
    NOR2X1 U31356 (.A1(n28501), .A2(N5942), .ZN(n44228));
    NOR2X1 U31357 (.A1(n43269), .A2(N9715), .ZN(N44229));
    NANDX1 U31358 (.A1(N4592), .A2(N1147), .ZN(N44230));
    INVX1 U31359 (.I(n15490), .ZN(n44231));
    NOR2X1 U31360 (.A1(n30830), .A2(n15172), .ZN(N44232));
    NANDX1 U31361 (.A1(N11821), .A2(n15086), .ZN(N44233));
    NANDX1 U31362 (.A1(N11073), .A2(n37110), .ZN(N44234));
    NANDX1 U31363 (.A1(n23966), .A2(N7691), .ZN(N44235));
    NANDX1 U31364 (.A1(n24710), .A2(n17718), .ZN(N44236));
    NOR2X1 U31365 (.A1(N10690), .A2(n35437), .ZN(N44237));
    INVX1 U31366 (.I(n18823), .ZN(N44238));
    NOR2X1 U31367 (.A1(n34792), .A2(n24764), .ZN(N44239));
    NOR2X1 U31368 (.A1(n34588), .A2(n24158), .ZN(N44240));
    NANDX1 U31369 (.A1(n39180), .A2(n14984), .ZN(N44241));
    NANDX1 U31370 (.A1(N877), .A2(n31234), .ZN(N44242));
    INVX1 U31371 (.I(N5728), .ZN(N44243));
    NOR2X1 U31372 (.A1(n17249), .A2(n20813), .ZN(N44244));
    INVX1 U31373 (.I(n18001), .ZN(n44245));
    NANDX1 U31374 (.A1(n28431), .A2(n31646), .ZN(N44246));
    NOR2X1 U31375 (.A1(n39296), .A2(n12883), .ZN(n44247));
    NANDX1 U31376 (.A1(N7572), .A2(n13252), .ZN(N44248));
    NANDX1 U31377 (.A1(n13863), .A2(n32074), .ZN(N44249));
    INVX1 U31378 (.I(N5182), .ZN(N44250));
    NANDX1 U31379 (.A1(n41126), .A2(n39769), .ZN(N44251));
    NANDX1 U31380 (.A1(N5119), .A2(n25156), .ZN(N44252));
    INVX1 U31381 (.I(n23190), .ZN(n44253));
    NANDX1 U31382 (.A1(N9307), .A2(n28618), .ZN(N44254));
    NOR2X1 U31383 (.A1(n31279), .A2(n35546), .ZN(N44255));
    INVX1 U31384 (.I(n13102), .ZN(N44256));
    NOR2X1 U31385 (.A1(N2911), .A2(n41533), .ZN(N44257));
    NOR2X1 U31386 (.A1(N4411), .A2(n37356), .ZN(N44258));
    NOR2X1 U31387 (.A1(n23629), .A2(n34607), .ZN(N44259));
    NANDX1 U31388 (.A1(n24491), .A2(N4997), .ZN(n44260));
    INVX1 U31389 (.I(N12198), .ZN(N44261));
    NOR2X1 U31390 (.A1(n18217), .A2(N9851), .ZN(N44262));
    NOR2X1 U31391 (.A1(n24778), .A2(N4650), .ZN(N44263));
    INVX1 U31392 (.I(N2851), .ZN(N44264));
    INVX1 U31393 (.I(n37022), .ZN(N44265));
    NOR2X1 U31394 (.A1(N2664), .A2(n14990), .ZN(N44266));
    INVX1 U31395 (.I(n27889), .ZN(N44267));
    NOR2X1 U31396 (.A1(N2745), .A2(n27642), .ZN(N44268));
    INVX1 U31397 (.I(N805), .ZN(N44269));
    NOR2X1 U31398 (.A1(n21090), .A2(n27840), .ZN(n44270));
    NOR2X1 U31399 (.A1(n34398), .A2(n18975), .ZN(N44271));
    INVX1 U31400 (.I(N5096), .ZN(N44272));
    INVX1 U31401 (.I(N4327), .ZN(N44273));
    INVX1 U31402 (.I(n13509), .ZN(N44274));
    INVX1 U31403 (.I(n16824), .ZN(N44275));
    INVX1 U31404 (.I(N3848), .ZN(N44276));
    INVX1 U31405 (.I(N10332), .ZN(N44277));
    NANDX1 U31406 (.A1(n38991), .A2(n37034), .ZN(N44278));
    NANDX1 U31407 (.A1(n31334), .A2(N8551), .ZN(N44279));
    NOR2X1 U31408 (.A1(n15750), .A2(N12000), .ZN(n44280));
    NANDX1 U31409 (.A1(n33071), .A2(n28679), .ZN(N44281));
    NOR2X1 U31410 (.A1(n27998), .A2(n39448), .ZN(N44282));
    NOR2X1 U31411 (.A1(n13413), .A2(n20054), .ZN(N44283));
    NOR2X1 U31412 (.A1(n35719), .A2(n25149), .ZN(N44284));
    INVX1 U31413 (.I(n40045), .ZN(N44285));
    NOR2X1 U31414 (.A1(N1266), .A2(N8795), .ZN(N44286));
    NOR2X1 U31415 (.A1(n33760), .A2(N2322), .ZN(n44287));
    NOR2X1 U31416 (.A1(N619), .A2(n42172), .ZN(N44288));
    NANDX1 U31417 (.A1(n27332), .A2(n40387), .ZN(N44289));
    NANDX1 U31418 (.A1(n35882), .A2(n17924), .ZN(N44290));
    NOR2X1 U31419 (.A1(n37561), .A2(n41677), .ZN(N44291));
    INVX1 U31420 (.I(n22767), .ZN(N44292));
    NOR2X1 U31421 (.A1(N12708), .A2(N8423), .ZN(N44293));
    NOR2X1 U31422 (.A1(n15800), .A2(n28476), .ZN(N44294));
    NOR2X1 U31423 (.A1(N8046), .A2(N10152), .ZN(N44295));
    INVX1 U31424 (.I(N4618), .ZN(N44296));
    NANDX1 U31425 (.A1(N7327), .A2(N3092), .ZN(N44297));
    NANDX1 U31426 (.A1(n41086), .A2(N5413), .ZN(N44298));
    INVX1 U31427 (.I(n31384), .ZN(N44299));
    INVX1 U31428 (.I(n22719), .ZN(N44300));
    NANDX1 U31429 (.A1(n23859), .A2(N12402), .ZN(N44301));
    INVX1 U31430 (.I(n41782), .ZN(N44302));
    INVX1 U31431 (.I(n34894), .ZN(N44303));
    INVX1 U31432 (.I(N2544), .ZN(N44304));
    INVX1 U31433 (.I(N8955), .ZN(N44305));
    NANDX1 U31434 (.A1(N12290), .A2(n30320), .ZN(N44306));
    NANDX1 U31435 (.A1(n40765), .A2(n15472), .ZN(N44307));
    NOR2X1 U31436 (.A1(n40597), .A2(n31853), .ZN(N44308));
    NANDX1 U31437 (.A1(n39397), .A2(n28859), .ZN(N44309));
    NOR2X1 U31438 (.A1(n33350), .A2(n26472), .ZN(N44310));
    INVX1 U31439 (.I(N454), .ZN(N44311));
    INVX1 U31440 (.I(N4728), .ZN(N44312));
    NOR2X1 U31441 (.A1(n19307), .A2(n28586), .ZN(N44313));
    INVX1 U31442 (.I(N6319), .ZN(N44314));
    INVX1 U31443 (.I(n32768), .ZN(n44315));
    NOR2X1 U31444 (.A1(n13088), .A2(n24991), .ZN(N44316));
    INVX1 U31445 (.I(N11722), .ZN(N44317));
    NOR2X1 U31446 (.A1(N3577), .A2(n31721), .ZN(N44318));
    NANDX1 U31447 (.A1(n34022), .A2(N3721), .ZN(N44319));
    NOR2X1 U31448 (.A1(n31146), .A2(n25253), .ZN(N44320));
    INVX1 U31449 (.I(n16750), .ZN(N44321));
    INVX1 U31450 (.I(n23268), .ZN(N44322));
    NANDX1 U31451 (.A1(n26791), .A2(n34203), .ZN(N44323));
    NANDX1 U31452 (.A1(n30854), .A2(n38930), .ZN(N44324));
    INVX1 U31453 (.I(n39840), .ZN(N44325));
    NANDX1 U31454 (.A1(n14226), .A2(n35839), .ZN(N44326));
    NANDX1 U31455 (.A1(N3521), .A2(n23258), .ZN(N44327));
    NANDX1 U31456 (.A1(n28512), .A2(n14545), .ZN(N44328));
    INVX1 U31457 (.I(N4641), .ZN(N44329));
    NOR2X1 U31458 (.A1(n33033), .A2(N1499), .ZN(N44330));
    INVX1 U31459 (.I(n26433), .ZN(N44331));
    NANDX1 U31460 (.A1(n19176), .A2(n41366), .ZN(N44332));
    INVX1 U31461 (.I(n35925), .ZN(N44333));
    NANDX1 U31462 (.A1(n37184), .A2(n21912), .ZN(N44334));
    NOR2X1 U31463 (.A1(n17594), .A2(N8352), .ZN(N44335));
    NOR2X1 U31464 (.A1(n13051), .A2(n40796), .ZN(n44336));
    INVX1 U31465 (.I(n26773), .ZN(n44337));
    NOR2X1 U31466 (.A1(n23950), .A2(N3277), .ZN(N44338));
    NANDX1 U31467 (.A1(N3736), .A2(n36340), .ZN(N44339));
    NOR2X1 U31468 (.A1(n18280), .A2(n37652), .ZN(n44340));
    INVX1 U31469 (.I(n26081), .ZN(N44341));
    NANDX1 U31470 (.A1(n29079), .A2(n14111), .ZN(N44342));
    NOR2X1 U31471 (.A1(n25251), .A2(n33286), .ZN(N44343));
    NOR2X1 U31472 (.A1(n39167), .A2(n15419), .ZN(n44344));
    NANDX1 U31473 (.A1(n22558), .A2(n37330), .ZN(N44345));
    INVX1 U31474 (.I(n40151), .ZN(N44346));
    NOR2X1 U31475 (.A1(N12704), .A2(n42881), .ZN(N44347));
    INVX1 U31476 (.I(N816), .ZN(N44348));
    NANDX1 U31477 (.A1(n33912), .A2(n24765), .ZN(N44349));
    NOR2X1 U31478 (.A1(n38661), .A2(n28500), .ZN(N44350));
    NOR2X1 U31479 (.A1(n18129), .A2(n36460), .ZN(n44351));
    INVX1 U31480 (.I(N12557), .ZN(N44352));
    NANDX1 U31481 (.A1(n23074), .A2(n31316), .ZN(N44353));
    NANDX1 U31482 (.A1(n22926), .A2(n13094), .ZN(N44354));
    NOR2X1 U31483 (.A1(n20671), .A2(n41940), .ZN(N44355));
    NANDX1 U31484 (.A1(n16628), .A2(N10705), .ZN(N44356));
    INVX1 U31485 (.I(n27268), .ZN(N44357));
    INVX1 U31486 (.I(N3515), .ZN(n44358));
    NANDX1 U31487 (.A1(n39943), .A2(n25878), .ZN(N44359));
    INVX1 U31488 (.I(N2011), .ZN(N44360));
    NOR2X1 U31489 (.A1(N11759), .A2(n21147), .ZN(n44361));
    NANDX1 U31490 (.A1(n29938), .A2(n22830), .ZN(n44362));
    INVX1 U31491 (.I(N12605), .ZN(N44363));
    INVX1 U31492 (.I(N11231), .ZN(N44364));
    NANDX1 U31493 (.A1(n31445), .A2(n42546), .ZN(N44365));
    NOR2X1 U31494 (.A1(N579), .A2(N1847), .ZN(N44366));
    NOR2X1 U31495 (.A1(N10929), .A2(N314), .ZN(N44367));
    NOR2X1 U31496 (.A1(n17237), .A2(N11018), .ZN(N44368));
    INVX1 U31497 (.I(N1032), .ZN(N44369));
    INVX1 U31498 (.I(n25681), .ZN(N44370));
    NOR2X1 U31499 (.A1(n37702), .A2(n41238), .ZN(N44371));
    INVX1 U31500 (.I(n39712), .ZN(N44372));
    INVX1 U31501 (.I(n29434), .ZN(N44373));
    NANDX1 U31502 (.A1(n38101), .A2(N5579), .ZN(n44374));
    NOR2X1 U31503 (.A1(n36775), .A2(n18184), .ZN(N44375));
    INVX1 U31504 (.I(N4533), .ZN(N44376));
    NANDX1 U31505 (.A1(n26239), .A2(n36759), .ZN(N44377));
    NANDX1 U31506 (.A1(n26817), .A2(n38605), .ZN(N44378));
    NANDX1 U31507 (.A1(n27425), .A2(n28599), .ZN(N44379));
    NANDX1 U31508 (.A1(N1189), .A2(n29296), .ZN(N44380));
    NOR2X1 U31509 (.A1(N2220), .A2(n27056), .ZN(N44381));
    INVX1 U31510 (.I(n32902), .ZN(n44382));
    NOR2X1 U31511 (.A1(n25081), .A2(n40257), .ZN(n44383));
    NANDX1 U31512 (.A1(n28844), .A2(n15898), .ZN(N44384));
    INVX1 U31513 (.I(n13152), .ZN(N44385));
    NOR2X1 U31514 (.A1(N11013), .A2(N6454), .ZN(N44386));
    INVX1 U31515 (.I(N5806), .ZN(N44387));
    NOR2X1 U31516 (.A1(n15082), .A2(n21724), .ZN(N44388));
    INVX1 U31517 (.I(n34715), .ZN(N44389));
    NANDX1 U31518 (.A1(N11917), .A2(N3646), .ZN(N44390));
    INVX1 U31519 (.I(n40515), .ZN(N44391));
    NOR2X1 U31520 (.A1(n23361), .A2(n16018), .ZN(N44392));
    NOR2X1 U31521 (.A1(n15261), .A2(n43073), .ZN(N44393));
    INVX1 U31522 (.I(n37842), .ZN(N44394));
    INVX1 U31523 (.I(n37146), .ZN(N44395));
    NANDX1 U31524 (.A1(n28090), .A2(N12197), .ZN(N44396));
    INVX1 U31525 (.I(n42359), .ZN(N44397));
    NOR2X1 U31526 (.A1(n18206), .A2(N9899), .ZN(n44398));
    NANDX1 U31527 (.A1(n37225), .A2(N5385), .ZN(N44399));
    NANDX1 U31528 (.A1(N8834), .A2(n16788), .ZN(N44400));
    NOR2X1 U31529 (.A1(N77), .A2(N11536), .ZN(N44401));
    NANDX1 U31530 (.A1(N3722), .A2(n23388), .ZN(N44402));
    NANDX1 U31531 (.A1(n30308), .A2(N3276), .ZN(N44403));
    NANDX1 U31532 (.A1(n15058), .A2(N8216), .ZN(N44404));
    NOR2X1 U31533 (.A1(n27122), .A2(N2585), .ZN(N44405));
    NOR2X1 U31534 (.A1(n20795), .A2(n26890), .ZN(N44406));
    NANDX1 U31535 (.A1(n22671), .A2(n23620), .ZN(N44407));
    INVX1 U31536 (.I(n37698), .ZN(N44408));
    NOR2X1 U31537 (.A1(n26193), .A2(N5386), .ZN(N44409));
    NANDX1 U31538 (.A1(n31577), .A2(n17212), .ZN(N44410));
    NOR2X1 U31539 (.A1(N4892), .A2(N2349), .ZN(N44411));
    INVX1 U31540 (.I(N6107), .ZN(N44412));
    INVX1 U31541 (.I(n17248), .ZN(N44413));
    NOR2X1 U31542 (.A1(n36969), .A2(n37236), .ZN(N44414));
    NANDX1 U31543 (.A1(n36761), .A2(N8821), .ZN(N44415));
    NANDX1 U31544 (.A1(n25834), .A2(n35942), .ZN(N44416));
    INVX1 U31545 (.I(n35792), .ZN(N44417));
    INVX1 U31546 (.I(N6347), .ZN(N44418));
    NANDX1 U31547 (.A1(n15295), .A2(n29967), .ZN(N44419));
    NOR2X1 U31548 (.A1(N9521), .A2(n18000), .ZN(N44420));
    INVX1 U31549 (.I(N4586), .ZN(N44421));
    INVX1 U31550 (.I(n40317), .ZN(N44422));
    NOR2X1 U31551 (.A1(n23555), .A2(n34888), .ZN(N44423));
    INVX1 U31552 (.I(n37082), .ZN(N44424));
    INVX1 U31553 (.I(N2906), .ZN(N44425));
    NOR2X1 U31554 (.A1(n16696), .A2(n39874), .ZN(N44426));
    NANDX1 U31555 (.A1(n39145), .A2(n22843), .ZN(N44427));
    INVX1 U31556 (.I(n26338), .ZN(N44428));
    NANDX1 U31557 (.A1(n18422), .A2(N5795), .ZN(N44429));
    NOR2X1 U31558 (.A1(n21366), .A2(N1821), .ZN(N44430));
    INVX1 U31559 (.I(n36660), .ZN(N44431));
    INVX1 U31560 (.I(n33270), .ZN(N44432));
    NOR2X1 U31561 (.A1(n39466), .A2(n42010), .ZN(N44433));
    NANDX1 U31562 (.A1(n28930), .A2(n38854), .ZN(N44434));
    INVX1 U31563 (.I(n42165), .ZN(N44435));
    NOR2X1 U31564 (.A1(N1635), .A2(n35774), .ZN(N44436));
    NOR2X1 U31565 (.A1(N4540), .A2(n25990), .ZN(N44437));
    INVX1 U31566 (.I(n34094), .ZN(N44438));
    NANDX1 U31567 (.A1(n19520), .A2(n13464), .ZN(n44439));
    NOR2X1 U31568 (.A1(n35537), .A2(N8347), .ZN(N44440));
    NANDX1 U31569 (.A1(n31011), .A2(n39022), .ZN(N44441));
    NANDX1 U31570 (.A1(n32831), .A2(n25632), .ZN(N44442));
    NANDX1 U31571 (.A1(N10826), .A2(N5109), .ZN(N44443));
    INVX1 U31572 (.I(n39971), .ZN(N44444));
    INVX1 U31573 (.I(n37615), .ZN(N44445));
    INVX1 U31574 (.I(n32180), .ZN(N44446));
    INVX1 U31575 (.I(n24121), .ZN(N44447));
    INVX1 U31576 (.I(n27059), .ZN(N44448));
    INVX1 U31577 (.I(n15808), .ZN(n44449));
    NOR2X1 U31578 (.A1(n32091), .A2(n39655), .ZN(N44450));
    NANDX1 U31579 (.A1(n42060), .A2(N5382), .ZN(N44451));
    INVX1 U31580 (.I(N1357), .ZN(N44452));
    NANDX1 U31581 (.A1(n23389), .A2(n22546), .ZN(N44453));
    INVX1 U31582 (.I(n18938), .ZN(n44454));
    NOR2X1 U31583 (.A1(N7494), .A2(n34249), .ZN(n44455));
    INVX1 U31584 (.I(N7999), .ZN(N44456));
    INVX1 U31585 (.I(n13260), .ZN(N44457));
    NANDX1 U31586 (.A1(n32684), .A2(N7403), .ZN(N44458));
    NOR2X1 U31587 (.A1(n21391), .A2(n22507), .ZN(N44459));
    NOR2X1 U31588 (.A1(n30048), .A2(N6093), .ZN(n44460));
    INVX1 U31589 (.I(n35535), .ZN(N44461));
    INVX1 U31590 (.I(n28125), .ZN(N44462));
    NOR2X1 U31591 (.A1(n39269), .A2(n16393), .ZN(N44463));
    INVX1 U31592 (.I(N10838), .ZN(N44464));
    NANDX1 U31593 (.A1(n24223), .A2(n34226), .ZN(N44465));
    NANDX1 U31594 (.A1(n42358), .A2(n42844), .ZN(N44466));
    INVX1 U31595 (.I(n39532), .ZN(N44467));
    NOR2X1 U31596 (.A1(n36732), .A2(n37210), .ZN(n44468));
    INVX1 U31597 (.I(N6520), .ZN(N44469));
    INVX1 U31598 (.I(N8396), .ZN(N44470));
    INVX1 U31599 (.I(n17840), .ZN(N44471));
    NANDX1 U31600 (.A1(n26108), .A2(N7773), .ZN(N44472));
    NOR2X1 U31601 (.A1(n21880), .A2(N3807), .ZN(N44473));
    INVX1 U31602 (.I(N5777), .ZN(N44474));
    INVX1 U31603 (.I(n29821), .ZN(N44475));
    NOR2X1 U31604 (.A1(n27684), .A2(n13126), .ZN(N44476));
    INVX1 U31605 (.I(n35112), .ZN(n44477));
    NOR2X1 U31606 (.A1(n36316), .A2(N11293), .ZN(N44478));
    NANDX1 U31607 (.A1(n25367), .A2(n31935), .ZN(N44479));
    NANDX1 U31608 (.A1(n15515), .A2(n14874), .ZN(N44480));
    NANDX1 U31609 (.A1(n24379), .A2(n21393), .ZN(N44481));
    NOR2X1 U31610 (.A1(n32775), .A2(n14674), .ZN(N44482));
    INVX1 U31611 (.I(n19089), .ZN(N44483));
    NOR2X1 U31612 (.A1(N8597), .A2(n14810), .ZN(N44484));
    NANDX1 U31613 (.A1(N2084), .A2(n12913), .ZN(n44485));
    NOR2X1 U31614 (.A1(n13375), .A2(n32413), .ZN(N44486));
    NANDX1 U31615 (.A1(n41058), .A2(n35219), .ZN(n44487));
    NOR2X1 U31616 (.A1(n32697), .A2(n18775), .ZN(N44488));
    INVX1 U31617 (.I(n33669), .ZN(N44489));
    INVX1 U31618 (.I(N5557), .ZN(n44490));
    NOR2X1 U31619 (.A1(N2549), .A2(n21071), .ZN(N44491));
    NANDX1 U31620 (.A1(n41091), .A2(n35130), .ZN(N44492));
    NOR2X1 U31621 (.A1(n34395), .A2(n24432), .ZN(N44493));
    NANDX1 U31622 (.A1(n24899), .A2(n33200), .ZN(N44494));
    NANDX1 U31623 (.A1(n23176), .A2(N4537), .ZN(N44495));
    NANDX1 U31624 (.A1(n25259), .A2(N7129), .ZN(N44496));
    INVX1 U31625 (.I(n28313), .ZN(N44497));
    NANDX1 U31626 (.A1(n25355), .A2(n15578), .ZN(N44498));
    INVX1 U31627 (.I(n23022), .ZN(N44499));
    NOR2X1 U31628 (.A1(n39742), .A2(N3212), .ZN(N44500));
    NOR2X1 U31629 (.A1(n30637), .A2(N8768), .ZN(n44501));
    NOR2X1 U31630 (.A1(n22865), .A2(n19519), .ZN(N44502));
    NANDX1 U31631 (.A1(N10163), .A2(N11176), .ZN(N44503));
    INVX1 U31632 (.I(n34238), .ZN(N44504));
    INVX1 U31633 (.I(N3583), .ZN(N44505));
    INVX1 U31634 (.I(n15014), .ZN(N44506));
    NANDX1 U31635 (.A1(n38839), .A2(N9230), .ZN(N44507));
    NOR2X1 U31636 (.A1(N10305), .A2(n16358), .ZN(N44508));
    INVX1 U31637 (.I(n38617), .ZN(N44509));
    NANDX1 U31638 (.A1(n26324), .A2(N10722), .ZN(N44510));
    NOR2X1 U31639 (.A1(N5873), .A2(N5203), .ZN(N44511));
    INVX1 U31640 (.I(n42236), .ZN(N44512));
    INVX1 U31641 (.I(n29340), .ZN(N44513));
    NANDX1 U31642 (.A1(n29841), .A2(n41884), .ZN(N44514));
    NOR2X1 U31643 (.A1(N9541), .A2(N8575), .ZN(N44515));
    NANDX1 U31644 (.A1(n37317), .A2(n42812), .ZN(N44516));
    NOR2X1 U31645 (.A1(n40900), .A2(N4683), .ZN(N44517));
    NANDX1 U31646 (.A1(n40429), .A2(N50), .ZN(N44518));
    NANDX1 U31647 (.A1(N11620), .A2(N10354), .ZN(N44519));
    NANDX1 U31648 (.A1(N12589), .A2(n38651), .ZN(N44520));
    NANDX1 U31649 (.A1(n38912), .A2(n39052), .ZN(N44521));
    INVX1 U31650 (.I(n34465), .ZN(N44522));
    NANDX1 U31651 (.A1(N10089), .A2(n33228), .ZN(N44523));
    NOR2X1 U31652 (.A1(n29108), .A2(n30439), .ZN(n44524));
    INVX1 U31653 (.I(n17199), .ZN(N44525));
    NANDX1 U31654 (.A1(n42555), .A2(n25773), .ZN(N44526));
    INVX1 U31655 (.I(n36399), .ZN(N44527));
    INVX1 U31656 (.I(N8166), .ZN(N44528));
    INVX1 U31657 (.I(n19475), .ZN(N44529));
    NANDX1 U31658 (.A1(N10142), .A2(N9204), .ZN(N44530));
    NOR2X1 U31659 (.A1(n21761), .A2(N9237), .ZN(N44531));
    NOR2X1 U31660 (.A1(n34349), .A2(N4415), .ZN(N44532));
    NANDX1 U31661 (.A1(n19469), .A2(n33147), .ZN(N44533));
    NOR2X1 U31662 (.A1(N141), .A2(n23609), .ZN(N44534));
    NANDX1 U31663 (.A1(n23048), .A2(n26783), .ZN(n44535));
    NOR2X1 U31664 (.A1(N10015), .A2(n16325), .ZN(N44536));
    NANDX1 U31665 (.A1(n24030), .A2(n15407), .ZN(N44537));
    NANDX1 U31666 (.A1(N12158), .A2(n41485), .ZN(N44538));
    INVX1 U31667 (.I(n20323), .ZN(N44539));
    INVX1 U31668 (.I(n40968), .ZN(N44540));
    INVX1 U31669 (.I(n21340), .ZN(N44541));
    NANDX1 U31670 (.A1(n22812), .A2(n43101), .ZN(n44542));
    INVX1 U31671 (.I(n42722), .ZN(N44543));
    NOR2X1 U31672 (.A1(N10030), .A2(N7472), .ZN(N44544));
    INVX1 U31673 (.I(n32856), .ZN(N44545));
    INVX1 U31674 (.I(n43265), .ZN(n44546));
    NANDX1 U31675 (.A1(n25815), .A2(n22841), .ZN(N44547));
    INVX1 U31676 (.I(N10186), .ZN(N44548));
    INVX1 U31677 (.I(N2306), .ZN(N44549));
    NANDX1 U31678 (.A1(N3092), .A2(N7392), .ZN(N44550));
    INVX1 U31679 (.I(N4929), .ZN(N44551));
    INVX1 U31680 (.I(n17117), .ZN(N44552));
    NANDX1 U31681 (.A1(N6282), .A2(N4292), .ZN(N44553));
    NOR2X1 U31682 (.A1(n17302), .A2(N10990), .ZN(N44554));
    NOR2X1 U31683 (.A1(n16930), .A2(n16605), .ZN(N44555));
    NOR2X1 U31684 (.A1(n40586), .A2(n26634), .ZN(N44556));
    INVX1 U31685 (.I(n29919), .ZN(N44557));
    INVX1 U31686 (.I(N6858), .ZN(N44558));
    INVX1 U31687 (.I(N8368), .ZN(N44559));
    NANDX1 U31688 (.A1(n42231), .A2(n37821), .ZN(N44560));
    NOR2X1 U31689 (.A1(n21293), .A2(n29806), .ZN(N44561));
    INVX1 U31690 (.I(n14065), .ZN(N44562));
    INVX1 U31691 (.I(n29595), .ZN(N44563));
    NOR2X1 U31692 (.A1(n21960), .A2(n36392), .ZN(N44564));
    INVX1 U31693 (.I(n28242), .ZN(n44565));
    NOR2X1 U31694 (.A1(n15130), .A2(N2071), .ZN(N44566));
    NOR2X1 U31695 (.A1(n19148), .A2(N8680), .ZN(N44567));
    NOR2X1 U31696 (.A1(N12095), .A2(n38945), .ZN(N44568));
    NOR2X1 U31697 (.A1(N12513), .A2(n25391), .ZN(N44569));
    INVX1 U31698 (.I(n19371), .ZN(N44570));
    NOR2X1 U31699 (.A1(N1389), .A2(n41723), .ZN(n44571));
    NOR2X1 U31700 (.A1(n28889), .A2(n30788), .ZN(N44572));
    NANDX1 U31701 (.A1(n15222), .A2(n31607), .ZN(N44573));
    NOR2X1 U31702 (.A1(n42098), .A2(N7409), .ZN(N44574));
    NANDX1 U31703 (.A1(n20585), .A2(n33480), .ZN(N44575));
    INVX1 U31704 (.I(N5354), .ZN(N44576));
    NOR2X1 U31705 (.A1(N6206), .A2(n40576), .ZN(N44577));
    NANDX1 U31706 (.A1(n25353), .A2(n38935), .ZN(N44578));
    NANDX1 U31707 (.A1(n37447), .A2(n34408), .ZN(N44579));
    NANDX1 U31708 (.A1(n39640), .A2(N6006), .ZN(N44580));
    NOR2X1 U31709 (.A1(n15538), .A2(N7315), .ZN(N44581));
    NANDX1 U31710 (.A1(n13788), .A2(N7383), .ZN(N44582));
    NANDX1 U31711 (.A1(n34255), .A2(n18423), .ZN(N44583));
    NOR2X1 U31712 (.A1(N12069), .A2(n33207), .ZN(n44584));
    NANDX1 U31713 (.A1(n19477), .A2(n33831), .ZN(N44585));
    NOR2X1 U31714 (.A1(n42637), .A2(n24907), .ZN(N44586));
    NOR2X1 U31715 (.A1(n19535), .A2(n20793), .ZN(N44587));
    NANDX1 U31716 (.A1(n27465), .A2(N2673), .ZN(N44588));
    NOR2X1 U31717 (.A1(n39559), .A2(n29800), .ZN(N44589));
    NANDX1 U31718 (.A1(n38978), .A2(n25967), .ZN(N44590));
    INVX1 U31719 (.I(n21098), .ZN(n44591));
    INVX1 U31720 (.I(n40874), .ZN(N44592));
    NANDX1 U31721 (.A1(n34651), .A2(n37936), .ZN(N44593));
    INVX1 U31722 (.I(n25433), .ZN(N44594));
    INVX1 U31723 (.I(N3339), .ZN(N44595));
    NANDX1 U31724 (.A1(n35772), .A2(N8941), .ZN(N44596));
    NANDX1 U31725 (.A1(n26130), .A2(n35127), .ZN(N44597));
    INVX1 U31726 (.I(n40717), .ZN(N44598));
    INVX1 U31727 (.I(N11563), .ZN(N44599));
    NANDX1 U31728 (.A1(n20879), .A2(n39027), .ZN(N44600));
    NOR2X1 U31729 (.A1(n24345), .A2(n24793), .ZN(N44601));
    NOR2X1 U31730 (.A1(n18746), .A2(N9978), .ZN(N44602));
    INVX1 U31731 (.I(N8832), .ZN(n44603));
    NOR2X1 U31732 (.A1(N73), .A2(N6233), .ZN(N44604));
    NANDX1 U31733 (.A1(n34723), .A2(N696), .ZN(N44605));
    NANDX1 U31734 (.A1(n16683), .A2(N3261), .ZN(N44606));
    NANDX1 U31735 (.A1(N391), .A2(n39032), .ZN(N44607));
    INVX1 U31736 (.I(n36728), .ZN(N44608));
    NANDX1 U31737 (.A1(n27846), .A2(n28756), .ZN(N44609));
    INVX1 U31738 (.I(n30400), .ZN(N44610));
    INVX1 U31739 (.I(N6010), .ZN(N44611));
    NOR2X1 U31740 (.A1(n25553), .A2(N6078), .ZN(N44612));
    NOR2X1 U31741 (.A1(N6874), .A2(n35946), .ZN(N44613));
    NANDX1 U31742 (.A1(n16851), .A2(N4835), .ZN(N44614));
    NOR2X1 U31743 (.A1(n37606), .A2(n38060), .ZN(N44615));
    NOR2X1 U31744 (.A1(n42325), .A2(n29310), .ZN(N44616));
    NANDX1 U31745 (.A1(n33086), .A2(n35673), .ZN(N44617));
    INVX1 U31746 (.I(n16864), .ZN(N44618));
    INVX1 U31747 (.I(n13875), .ZN(N44619));
    INVX1 U31748 (.I(n18998), .ZN(N44620));
    NOR2X1 U31749 (.A1(n27108), .A2(N4282), .ZN(N44621));
    NOR2X1 U31750 (.A1(n14035), .A2(n34280), .ZN(N44622));
    NOR2X1 U31751 (.A1(N11521), .A2(n16360), .ZN(n44623));
    NANDX1 U31752 (.A1(n33350), .A2(n12913), .ZN(n44624));
    INVX1 U31753 (.I(n20133), .ZN(N44625));
    NANDX1 U31754 (.A1(N12291), .A2(n15747), .ZN(N44626));
    INVX1 U31755 (.I(n40030), .ZN(N44627));
    INVX1 U31756 (.I(N2109), .ZN(N44628));
    NANDX1 U31757 (.A1(n32647), .A2(n24874), .ZN(N44629));
    NANDX1 U31758 (.A1(n17810), .A2(n41738), .ZN(N44630));
    INVX1 U31759 (.I(n21364), .ZN(N44631));
    NOR2X1 U31760 (.A1(n42167), .A2(n36287), .ZN(N44632));
    NANDX1 U31761 (.A1(n36128), .A2(n39183), .ZN(N44633));
    INVX1 U31762 (.I(n16615), .ZN(N44634));
    NOR2X1 U31763 (.A1(n39869), .A2(n32975), .ZN(N44635));
    INVX1 U31764 (.I(n19427), .ZN(N44636));
    NANDX1 U31765 (.A1(n27054), .A2(n39559), .ZN(N44637));
    NOR2X1 U31766 (.A1(n29024), .A2(N1513), .ZN(N44638));
    INVX1 U31767 (.I(n15261), .ZN(N44639));
    NANDX1 U31768 (.A1(N6583), .A2(n30807), .ZN(n44640));
    NANDX1 U31769 (.A1(n21136), .A2(n28234), .ZN(N44641));
    NOR2X1 U31770 (.A1(n19401), .A2(N7931), .ZN(n44642));
    NANDX1 U31771 (.A1(n16928), .A2(n39777), .ZN(N44643));
    NOR2X1 U31772 (.A1(n31242), .A2(n22113), .ZN(N44644));
    NOR2X1 U31773 (.A1(n16119), .A2(n38727), .ZN(N44645));
    NOR2X1 U31774 (.A1(N2195), .A2(n17909), .ZN(N44646));
    NOR2X1 U31775 (.A1(n21621), .A2(N10004), .ZN(N44647));
    NANDX1 U31776 (.A1(N7387), .A2(N11221), .ZN(N44648));
    NANDX1 U31777 (.A1(N8899), .A2(n15695), .ZN(N44649));
    INVX1 U31778 (.I(N7364), .ZN(N44650));
    NOR2X1 U31779 (.A1(n36299), .A2(N5323), .ZN(N44651));
    NOR2X1 U31780 (.A1(n21060), .A2(N451), .ZN(N44652));
    NOR2X1 U31781 (.A1(n28990), .A2(N6622), .ZN(N44653));
    INVX1 U31782 (.I(n14974), .ZN(N44654));
    INVX1 U31783 (.I(n36550), .ZN(N44655));
    NOR2X1 U31784 (.A1(n33454), .A2(n42348), .ZN(N44656));
    NANDX1 U31785 (.A1(n22444), .A2(n34222), .ZN(N44657));
    NANDX1 U31786 (.A1(n20711), .A2(N2051), .ZN(N44658));
    INVX1 U31787 (.I(n35712), .ZN(N44659));
    NANDX1 U31788 (.A1(n17681), .A2(n25943), .ZN(N44660));
    NANDX1 U31789 (.A1(n33375), .A2(n31435), .ZN(N44661));
    NOR2X1 U31790 (.A1(n35011), .A2(n24261), .ZN(N44662));
    NOR2X1 U31791 (.A1(n24630), .A2(N1848), .ZN(n44663));
    NOR2X1 U31792 (.A1(n13010), .A2(n20517), .ZN(N44664));
    INVX1 U31793 (.I(n18318), .ZN(n44665));
    NANDX1 U31794 (.A1(N2418), .A2(N1075), .ZN(N44666));
    NANDX1 U31795 (.A1(n35871), .A2(n33102), .ZN(N44667));
    NOR2X1 U31796 (.A1(n14842), .A2(n23851), .ZN(N44668));
    NANDX1 U31797 (.A1(n25232), .A2(n25901), .ZN(N44669));
    INVX1 U31798 (.I(n17471), .ZN(N44670));
    NANDX1 U31799 (.A1(n38568), .A2(n33094), .ZN(N44671));
    NOR2X1 U31800 (.A1(n18150), .A2(n21056), .ZN(N44672));
    NANDX1 U31801 (.A1(N9688), .A2(N1844), .ZN(N44673));
    NANDX1 U31802 (.A1(n23997), .A2(n36843), .ZN(N44674));
    INVX1 U31803 (.I(n37007), .ZN(N44675));
    NANDX1 U31804 (.A1(N12640), .A2(N11852), .ZN(N44676));
    INVX1 U31805 (.I(n15057), .ZN(N44677));
    NANDX1 U31806 (.A1(n24687), .A2(N7455), .ZN(N44678));
    NOR2X1 U31807 (.A1(n32338), .A2(N11976), .ZN(N44679));
    NOR2X1 U31808 (.A1(n36446), .A2(n26887), .ZN(N44680));
    NOR2X1 U31809 (.A1(n13861), .A2(N886), .ZN(N44681));
    NANDX1 U31810 (.A1(N8956), .A2(n23659), .ZN(N44682));
    INVX1 U31811 (.I(n16785), .ZN(N44683));
    INVX1 U31812 (.I(n30541), .ZN(N44684));
    NANDX1 U31813 (.A1(n36237), .A2(n35539), .ZN(N44685));
    INVX1 U31814 (.I(n19287), .ZN(N44686));
    INVX1 U31815 (.I(n33682), .ZN(N44687));
    NANDX1 U31816 (.A1(n43366), .A2(n35213), .ZN(N44688));
    NOR2X1 U31817 (.A1(N4630), .A2(n37818), .ZN(N44689));
    NOR2X1 U31818 (.A1(N12084), .A2(n30052), .ZN(N44690));
    NANDX1 U31819 (.A1(n13739), .A2(n35817), .ZN(N44691));
    NOR2X1 U31820 (.A1(n40625), .A2(n13690), .ZN(N44692));
    INVX1 U31821 (.I(n31190), .ZN(N44693));
    NOR2X1 U31822 (.A1(n16816), .A2(N11376), .ZN(N44694));
    INVX1 U31823 (.I(n33600), .ZN(N44695));
    NOR2X1 U31824 (.A1(n29250), .A2(N6279), .ZN(N44696));
    NANDX1 U31825 (.A1(N10996), .A2(n13275), .ZN(n44697));
    NOR2X1 U31826 (.A1(n41722), .A2(N3484), .ZN(N44698));
    INVX1 U31827 (.I(n41615), .ZN(N44699));
    INVX1 U31828 (.I(N1843), .ZN(N44700));
    NOR2X1 U31829 (.A1(n22722), .A2(n34645), .ZN(N44701));
    NOR2X1 U31830 (.A1(n42454), .A2(N2520), .ZN(N44702));
    INVX1 U31831 (.I(n24478), .ZN(n44703));
    NANDX1 U31832 (.A1(n38257), .A2(n38167), .ZN(N44704));
    NOR2X1 U31833 (.A1(n15655), .A2(N954), .ZN(N44705));
    INVX1 U31834 (.I(n16710), .ZN(N44706));
    INVX1 U31835 (.I(N11324), .ZN(N44707));
    INVX1 U31836 (.I(n18592), .ZN(n44708));
    NANDX1 U31837 (.A1(N3747), .A2(n19267), .ZN(N44709));
    NOR2X1 U31838 (.A1(N7774), .A2(n17516), .ZN(n44710));
    NANDX1 U31839 (.A1(n34652), .A2(N5338), .ZN(N44711));
    NANDX1 U31840 (.A1(n36494), .A2(n41261), .ZN(N44712));
    NANDX1 U31841 (.A1(n17346), .A2(n35475), .ZN(N44713));
    NANDX1 U31842 (.A1(n19866), .A2(n43427), .ZN(N44714));
    INVX1 U31843 (.I(n16386), .ZN(N44715));
    NOR2X1 U31844 (.A1(n18858), .A2(n31086), .ZN(N44716));
    INVX1 U31845 (.I(n19811), .ZN(N44717));
    INVX1 U31846 (.I(n16783), .ZN(N44718));
    NOR2X1 U31847 (.A1(N9814), .A2(n25469), .ZN(N44719));
    INVX1 U31848 (.I(n17096), .ZN(n44720));
    NANDX1 U31849 (.A1(n36690), .A2(n37652), .ZN(n44721));
    NANDX1 U31850 (.A1(N10733), .A2(n41051), .ZN(N44722));
    NOR2X1 U31851 (.A1(N5750), .A2(n29355), .ZN(N44723));
    NANDX1 U31852 (.A1(N3538), .A2(n40380), .ZN(N44724));
    NANDX1 U31853 (.A1(n39012), .A2(N6914), .ZN(N44725));
    INVX1 U31854 (.I(n28646), .ZN(N44726));
    INVX1 U31855 (.I(n33505), .ZN(n44727));
    NANDX1 U31856 (.A1(n39614), .A2(N10798), .ZN(N44728));
    NOR2X1 U31857 (.A1(N5632), .A2(N9288), .ZN(N44729));
    NANDX1 U31858 (.A1(n14784), .A2(n19101), .ZN(N44730));
    INVX1 U31859 (.I(n32207), .ZN(n44731));
    NOR2X1 U31860 (.A1(N10169), .A2(n25424), .ZN(N44732));
    NANDX1 U31861 (.A1(n36837), .A2(n25836), .ZN(N44733));
    NOR2X1 U31862 (.A1(N892), .A2(n31585), .ZN(N44734));
    NOR2X1 U31863 (.A1(n34592), .A2(n35122), .ZN(N44735));
    INVX1 U31864 (.I(n42166), .ZN(N44736));
    INVX1 U31865 (.I(n30167), .ZN(N44737));
    INVX1 U31866 (.I(n38666), .ZN(N44738));
    INVX1 U31867 (.I(N5845), .ZN(N44739));
    INVX1 U31868 (.I(n13912), .ZN(N44740));
    INVX1 U31869 (.I(N753), .ZN(N44741));
    INVX1 U31870 (.I(n25930), .ZN(N44742));
    NANDX1 U31871 (.A1(n24006), .A2(n34710), .ZN(N44743));
    NANDX1 U31872 (.A1(N12740), .A2(n17113), .ZN(N44744));
    NOR2X1 U31873 (.A1(n27843), .A2(n26847), .ZN(N44745));
    NANDX1 U31874 (.A1(N10206), .A2(n34159), .ZN(N44746));
    NOR2X1 U31875 (.A1(n31470), .A2(n27354), .ZN(n44747));
    INVX1 U31876 (.I(n23119), .ZN(N44748));
    NOR2X1 U31877 (.A1(n41206), .A2(n33139), .ZN(N44749));
    INVX1 U31878 (.I(N3226), .ZN(N44750));
    INVX1 U31879 (.I(N11600), .ZN(N44751));
    INVX1 U31880 (.I(n26269), .ZN(N44752));
    NOR2X1 U31881 (.A1(n15393), .A2(n16701), .ZN(N44753));
    INVX1 U31882 (.I(n31002), .ZN(N44754));
    INVX1 U31883 (.I(N4948), .ZN(N44755));
    INVX1 U31884 (.I(n40548), .ZN(N44756));
    NANDX1 U31885 (.A1(n29031), .A2(n31381), .ZN(N44757));
    NOR2X1 U31886 (.A1(N12405), .A2(N5258), .ZN(N44758));
    NOR2X1 U31887 (.A1(n36243), .A2(n13178), .ZN(N44759));
    NOR2X1 U31888 (.A1(n20124), .A2(N1898), .ZN(N44760));
    INVX1 U31889 (.I(n27259), .ZN(N44761));
    NOR2X1 U31890 (.A1(n15238), .A2(n21088), .ZN(N44762));
    INVX1 U31891 (.I(N97), .ZN(N44763));
    NOR2X1 U31892 (.A1(N1606), .A2(n16045), .ZN(N44764));
    NANDX1 U31893 (.A1(N6678), .A2(n32746), .ZN(n44765));
    NOR2X1 U31894 (.A1(n37679), .A2(n38837), .ZN(n44766));
    NANDX1 U31895 (.A1(N6125), .A2(n35912), .ZN(n44767));
    INVX1 U31896 (.I(n24835), .ZN(N44768));
    INVX1 U31897 (.I(N12230), .ZN(N44769));
    NANDX1 U31898 (.A1(n18758), .A2(n37005), .ZN(N44770));
    NOR2X1 U31899 (.A1(n31936), .A2(n16625), .ZN(N44771));
    INVX1 U31900 (.I(n23513), .ZN(N44772));
    INVX1 U31901 (.I(n13279), .ZN(N44773));
    NANDX1 U31902 (.A1(n13960), .A2(n34366), .ZN(N44774));
    NANDX1 U31903 (.A1(N3737), .A2(N2941), .ZN(N44775));
    INVX1 U31904 (.I(n19781), .ZN(N44776));
    NOR2X1 U31905 (.A1(N3321), .A2(N9054), .ZN(N44777));
    NANDX1 U31906 (.A1(n30680), .A2(N4418), .ZN(N44778));
    INVX1 U31907 (.I(n26484), .ZN(N44779));
    NANDX1 U31908 (.A1(N5672), .A2(N7847), .ZN(N44780));
    NANDX1 U31909 (.A1(N7581), .A2(n34765), .ZN(N44781));
    NOR2X1 U31910 (.A1(N1113), .A2(N10982), .ZN(N44782));
    INVX1 U31911 (.I(N7417), .ZN(N44783));
    NOR2X1 U31912 (.A1(n20450), .A2(n39292), .ZN(N44784));
    INVX1 U31913 (.I(n33272), .ZN(N44785));
    INVX1 U31914 (.I(n24007), .ZN(N44786));
    NOR2X1 U31915 (.A1(n13515), .A2(n26947), .ZN(N44787));
    INVX1 U31916 (.I(n33296), .ZN(N44788));
    NOR2X1 U31917 (.A1(n17953), .A2(n32029), .ZN(N44789));
    NOR2X1 U31918 (.A1(N5160), .A2(n26127), .ZN(n44790));
    INVX1 U31919 (.I(n21324), .ZN(N44791));
    NOR2X1 U31920 (.A1(n42858), .A2(n29170), .ZN(N44792));
    NANDX1 U31921 (.A1(N6967), .A2(N10142), .ZN(N44793));
    NANDX1 U31922 (.A1(n41231), .A2(N10804), .ZN(n44794));
    NOR2X1 U31923 (.A1(N5176), .A2(n40958), .ZN(N44795));
    NOR2X1 U31924 (.A1(N995), .A2(n40918), .ZN(n44796));
    INVX1 U31925 (.I(N453), .ZN(N44797));
    NOR2X1 U31926 (.A1(N2879), .A2(N3648), .ZN(N44798));
    NOR2X1 U31927 (.A1(n27831), .A2(n36943), .ZN(N44799));
    NOR2X1 U31928 (.A1(N2311), .A2(n15179), .ZN(n44800));
    NOR2X1 U31929 (.A1(n40623), .A2(n30985), .ZN(N44801));
    NOR2X1 U31930 (.A1(n18474), .A2(n33328), .ZN(N44802));
    NOR2X1 U31931 (.A1(n37323), .A2(n35708), .ZN(N44803));
    NANDX1 U31932 (.A1(N3992), .A2(n13411), .ZN(N44804));
    NANDX1 U31933 (.A1(N4475), .A2(n31523), .ZN(N44805));
    NANDX1 U31934 (.A1(N1960), .A2(n16292), .ZN(N44806));
    NANDX1 U31935 (.A1(n42878), .A2(n24013), .ZN(N44807));
    NOR2X1 U31936 (.A1(n20857), .A2(n26891), .ZN(N44808));
    INVX1 U31937 (.I(n25783), .ZN(N44809));
    NANDX1 U31938 (.A1(n18357), .A2(N888), .ZN(N44810));
    INVX1 U31939 (.I(n23215), .ZN(N44811));
    INVX1 U31940 (.I(n33542), .ZN(N44812));
    INVX1 U31941 (.I(N3164), .ZN(N44813));
    NOR2X1 U31942 (.A1(N583), .A2(N545), .ZN(N44814));
    NANDX1 U31943 (.A1(n36291), .A2(n38044), .ZN(N44815));
    NANDX1 U31944 (.A1(N6229), .A2(n40150), .ZN(N44816));
    NOR2X1 U31945 (.A1(n27431), .A2(n37110), .ZN(N44817));
    INVX1 U31946 (.I(n33402), .ZN(N44818));
    INVX1 U31947 (.I(n24735), .ZN(N44819));
    NANDX1 U31948 (.A1(N2512), .A2(n35272), .ZN(N44820));
    NOR2X1 U31949 (.A1(n37718), .A2(N7262), .ZN(N44821));
    NANDX1 U31950 (.A1(N2282), .A2(n41301), .ZN(n44822));
    NANDX1 U31951 (.A1(n25496), .A2(n36149), .ZN(N44823));
    INVX1 U31952 (.I(n36223), .ZN(N44824));
    NOR2X1 U31953 (.A1(n35484), .A2(n26486), .ZN(N44825));
    INVX1 U31954 (.I(n27556), .ZN(N44826));
    INVX1 U31955 (.I(n13788), .ZN(N44827));
    NOR2X1 U31956 (.A1(n15212), .A2(N10465), .ZN(N44828));
    NOR2X1 U31957 (.A1(n32322), .A2(n37255), .ZN(N44829));
    INVX1 U31958 (.I(N11931), .ZN(N44830));
    NOR2X1 U31959 (.A1(n32941), .A2(n15553), .ZN(N44831));
    INVX1 U31960 (.I(n14420), .ZN(N44832));
    NOR2X1 U31961 (.A1(n27795), .A2(n21681), .ZN(N44833));
    NANDX1 U31962 (.A1(n30076), .A2(n19509), .ZN(n44834));
    NOR2X1 U31963 (.A1(N1779), .A2(N1865), .ZN(N44835));
    INVX1 U31964 (.I(n38002), .ZN(N44836));
    INVX1 U31965 (.I(n36067), .ZN(N44837));
    NANDX1 U31966 (.A1(n39753), .A2(n20150), .ZN(N44838));
    NANDX1 U31967 (.A1(N10068), .A2(n23128), .ZN(N44839));
    INVX1 U31968 (.I(N10213), .ZN(N44840));
    NOR2X1 U31969 (.A1(n13418), .A2(n37147), .ZN(N44841));
    INVX1 U31970 (.I(n15028), .ZN(N44842));
    NANDX1 U31971 (.A1(N3679), .A2(n30581), .ZN(N44843));
    NANDX1 U31972 (.A1(n18099), .A2(N12534), .ZN(N44844));
    NOR2X1 U31973 (.A1(n29459), .A2(n15608), .ZN(N44845));
    NOR2X1 U31974 (.A1(N5496), .A2(n22402), .ZN(N44846));
    NOR2X1 U31975 (.A1(n40512), .A2(n22985), .ZN(N44847));
    NANDX1 U31976 (.A1(n17576), .A2(N5259), .ZN(N44848));
    NOR2X1 U31977 (.A1(n13856), .A2(n15088), .ZN(n44849));
    INVX1 U31978 (.I(n23924), .ZN(N44850));
    NOR2X1 U31979 (.A1(n26641), .A2(n23816), .ZN(N44851));
    NOR2X1 U31980 (.A1(n29738), .A2(n17490), .ZN(N44852));
    NOR2X1 U31981 (.A1(N1294), .A2(n42202), .ZN(N44853));
    INVX1 U31982 (.I(n21554), .ZN(N44854));
    NANDX1 U31983 (.A1(n16094), .A2(n34087), .ZN(N44855));
    NANDX1 U31984 (.A1(N2080), .A2(n39374), .ZN(N44856));
    INVX1 U31985 (.I(n40727), .ZN(N44857));
    NOR2X1 U31986 (.A1(n37436), .A2(n37767), .ZN(N44858));
    NANDX1 U31987 (.A1(n19458), .A2(N1550), .ZN(N44859));
    INVX1 U31988 (.I(N1853), .ZN(N44860));
    INVX1 U31989 (.I(n40992), .ZN(N44861));
    INVX1 U31990 (.I(n29009), .ZN(N44862));
    NOR2X1 U31991 (.A1(n30566), .A2(N9352), .ZN(N44863));
    NOR2X1 U31992 (.A1(n16832), .A2(n16521), .ZN(N44864));
    NANDX1 U31993 (.A1(N7805), .A2(n15250), .ZN(N44865));
    NANDX1 U31994 (.A1(n29358), .A2(n39088), .ZN(N44866));
    NOR2X1 U31995 (.A1(N9652), .A2(n39205), .ZN(N44867));
    INVX1 U31996 (.I(N5553), .ZN(N44868));
    NANDX1 U31997 (.A1(N2939), .A2(n13535), .ZN(N44869));
    NANDX1 U31998 (.A1(n30385), .A2(N1029), .ZN(N44870));
    INVX1 U31999 (.I(n31935), .ZN(N44871));
    INVX1 U32000 (.I(n19669), .ZN(N44872));
    NANDX1 U32001 (.A1(n24452), .A2(n13274), .ZN(N44873));
    NOR2X1 U32002 (.A1(N6393), .A2(N367), .ZN(N44874));
    NANDX1 U32003 (.A1(N11913), .A2(N6878), .ZN(N44875));
    NOR2X1 U32004 (.A1(n32390), .A2(n14682), .ZN(N44876));
    NOR2X1 U32005 (.A1(n40541), .A2(n33719), .ZN(N44877));
    NOR2X1 U32006 (.A1(n21314), .A2(n43370), .ZN(N44878));
    INVX1 U32007 (.I(n26998), .ZN(N44879));
    NANDX1 U32008 (.A1(N5626), .A2(n29936), .ZN(N44880));
    NOR2X1 U32009 (.A1(n14304), .A2(n16849), .ZN(N44881));
    NOR2X1 U32010 (.A1(n32120), .A2(N5311), .ZN(N44882));
    NOR2X1 U32011 (.A1(n41468), .A2(N9178), .ZN(N44883));
    NOR2X1 U32012 (.A1(N11269), .A2(n31733), .ZN(N44884));
    NOR2X1 U32013 (.A1(N1315), .A2(N9847), .ZN(N44885));
    INVX1 U32014 (.I(n41345), .ZN(N44886));
    INVX1 U32015 (.I(n37337), .ZN(n44887));
    NOR2X1 U32016 (.A1(n14364), .A2(n24086), .ZN(N44888));
    INVX1 U32017 (.I(n42694), .ZN(N44889));
    NANDX1 U32018 (.A1(n35850), .A2(n23284), .ZN(N44890));
    NOR2X1 U32019 (.A1(n30980), .A2(n28909), .ZN(N44891));
    INVX1 U32020 (.I(N6491), .ZN(n44892));
    INVX1 U32021 (.I(n21915), .ZN(N44893));
    INVX1 U32022 (.I(N11219), .ZN(N44894));
    NOR2X1 U32023 (.A1(n32166), .A2(N9214), .ZN(n44895));
    NOR2X1 U32024 (.A1(n39449), .A2(N10162), .ZN(N44896));
    NOR2X1 U32025 (.A1(n32484), .A2(N1157), .ZN(N44897));
    INVX1 U32026 (.I(n37431), .ZN(N44898));
    NOR2X1 U32027 (.A1(N8028), .A2(n31296), .ZN(N44899));
    NANDX1 U32028 (.A1(N12071), .A2(N11909), .ZN(N44900));
    NANDX1 U32029 (.A1(N11292), .A2(N3515), .ZN(N44901));
    INVX1 U32030 (.I(n34575), .ZN(N44902));
    INVX1 U32031 (.I(N6779), .ZN(N44903));
    NOR2X1 U32032 (.A1(n16864), .A2(N2949), .ZN(N44904));
    INVX1 U32033 (.I(n28459), .ZN(N44905));
    INVX1 U32034 (.I(N10329), .ZN(N44906));
    NOR2X1 U32035 (.A1(n40977), .A2(N9223), .ZN(N44907));
    INVX1 U32036 (.I(n36953), .ZN(N44908));
    INVX1 U32037 (.I(N1034), .ZN(N44909));
    NOR2X1 U32038 (.A1(n20540), .A2(N4582), .ZN(N44910));
    INVX1 U32039 (.I(N9248), .ZN(N44911));
    INVX1 U32040 (.I(n40897), .ZN(N44912));
    NOR2X1 U32041 (.A1(n24680), .A2(n42485), .ZN(N44913));
    INVX1 U32042 (.I(n25651), .ZN(N44914));
    NANDX1 U32043 (.A1(n13202), .A2(n16754), .ZN(N44915));
    NOR2X1 U32044 (.A1(n19980), .A2(n26444), .ZN(N44916));
    NANDX1 U32045 (.A1(n22929), .A2(n15234), .ZN(N44917));
    NOR2X1 U32046 (.A1(n31739), .A2(n25563), .ZN(N44918));
    NOR2X1 U32047 (.A1(n29243), .A2(n34785), .ZN(N44919));
    NOR2X1 U32048 (.A1(N12403), .A2(N376), .ZN(N44920));
    NOR2X1 U32049 (.A1(n28046), .A2(N10596), .ZN(N44921));
    INVX1 U32050 (.I(n27328), .ZN(N44922));
    INVX1 U32051 (.I(N2339), .ZN(N44923));
    INVX1 U32052 (.I(n20032), .ZN(N44924));
    NOR2X1 U32053 (.A1(n13445), .A2(n13963), .ZN(N44925));
    NOR2X1 U32054 (.A1(N5651), .A2(n27164), .ZN(N44926));
    NOR2X1 U32055 (.A1(n19975), .A2(N3672), .ZN(N44927));
    NOR2X1 U32056 (.A1(n40842), .A2(n26600), .ZN(N44928));
    INVX1 U32057 (.I(N3223), .ZN(N44929));
    NANDX1 U32058 (.A1(n18757), .A2(N646), .ZN(N44930));
    INVX1 U32059 (.I(n43221), .ZN(N44931));
    NOR2X1 U32060 (.A1(n35871), .A2(N124), .ZN(N44932));
    NANDX1 U32061 (.A1(N10125), .A2(N399), .ZN(N44933));
    NOR2X1 U32062 (.A1(n37452), .A2(N9922), .ZN(N44934));
    INVX1 U32063 (.I(N8411), .ZN(N44935));
    INVX1 U32064 (.I(N9637), .ZN(N44936));
    NOR2X1 U32065 (.A1(n33595), .A2(N8513), .ZN(n44937));
    NANDX1 U32066 (.A1(n17287), .A2(n24142), .ZN(N44938));
    INVX1 U32067 (.I(N10638), .ZN(N44939));
    NOR2X1 U32068 (.A1(n34529), .A2(n26917), .ZN(N44940));
    NOR2X1 U32069 (.A1(n27431), .A2(n31462), .ZN(N44941));
    NOR2X1 U32070 (.A1(n17756), .A2(N11458), .ZN(N44942));
    INVX1 U32071 (.I(N12837), .ZN(N44943));
    NANDX1 U32072 (.A1(n13924), .A2(N3387), .ZN(n44944));
    INVX1 U32073 (.I(N4002), .ZN(N44945));
    NOR2X1 U32074 (.A1(n41112), .A2(N3603), .ZN(N44946));
    INVX1 U32075 (.I(n39202), .ZN(N44947));
    INVX1 U32076 (.I(n40034), .ZN(N44948));
    INVX1 U32077 (.I(n13358), .ZN(N44949));
    NOR2X1 U32078 (.A1(n34770), .A2(n20324), .ZN(N44950));
    NOR2X1 U32079 (.A1(n28457), .A2(n30961), .ZN(n44951));
    NANDX1 U32080 (.A1(N9193), .A2(n14405), .ZN(N44952));
    NOR2X1 U32081 (.A1(n26303), .A2(N2395), .ZN(N44953));
    NOR2X1 U32082 (.A1(N586), .A2(N3532), .ZN(N44954));
    NANDX1 U32083 (.A1(N3103), .A2(n40540), .ZN(N44955));
    INVX1 U32084 (.I(n39641), .ZN(N44956));
    NOR2X1 U32085 (.A1(n41427), .A2(n23308), .ZN(N44957));
    NOR2X1 U32086 (.A1(n34710), .A2(n43385), .ZN(N44958));
    INVX1 U32087 (.I(n14473), .ZN(N44959));
    NOR2X1 U32088 (.A1(n34513), .A2(n17510), .ZN(N44960));
    NANDX1 U32089 (.A1(n25810), .A2(n37834), .ZN(N44961));
    INVX1 U32090 (.I(N10794), .ZN(N44962));
    NANDX1 U32091 (.A1(n33308), .A2(N9666), .ZN(N44963));
    NOR2X1 U32092 (.A1(n39279), .A2(n35968), .ZN(N44964));
    NOR2X1 U32093 (.A1(n15830), .A2(n26233), .ZN(N44965));
    NANDX1 U32094 (.A1(N6180), .A2(n29335), .ZN(N44966));
    NANDX1 U32095 (.A1(N133), .A2(n15184), .ZN(n44967));
    NANDX1 U32096 (.A1(n31239), .A2(n38491), .ZN(N44968));
    NANDX1 U32097 (.A1(n22476), .A2(n28083), .ZN(N44969));
    NOR2X1 U32098 (.A1(n26628), .A2(n14236), .ZN(n44970));
    INVX1 U32099 (.I(N666), .ZN(N44971));
    NOR2X1 U32100 (.A1(n34311), .A2(n28179), .ZN(N44972));
    INVX1 U32101 (.I(n34784), .ZN(N44973));
    NOR2X1 U32102 (.A1(N7609), .A2(N977), .ZN(N44974));
    NANDX1 U32103 (.A1(n36568), .A2(n36944), .ZN(n44975));
    NANDX1 U32104 (.A1(n42077), .A2(n19704), .ZN(N44976));
    INVX1 U32105 (.I(N4784), .ZN(N44977));
    NANDX1 U32106 (.A1(N10741), .A2(n38068), .ZN(N44978));
    INVX1 U32107 (.I(n23227), .ZN(N44979));
    INVX1 U32108 (.I(n38600), .ZN(N44980));
    NANDX1 U32109 (.A1(n27670), .A2(n23210), .ZN(N44981));
    INVX1 U32110 (.I(N505), .ZN(N44982));
    INVX1 U32111 (.I(n39402), .ZN(N44983));
    NANDX1 U32112 (.A1(N11946), .A2(n30240), .ZN(N44984));
    NANDX1 U32113 (.A1(n29719), .A2(n21551), .ZN(N44985));
    NOR2X1 U32114 (.A1(n27007), .A2(n22527), .ZN(N44986));
    INVX1 U32115 (.I(n20102), .ZN(n44987));
    NOR2X1 U32116 (.A1(N1179), .A2(n18706), .ZN(n44988));
    INVX1 U32117 (.I(n33312), .ZN(N44989));
    NANDX1 U32118 (.A1(n20628), .A2(n33732), .ZN(N44990));
    NOR2X1 U32119 (.A1(n20737), .A2(n13486), .ZN(N44991));
    NANDX1 U32120 (.A1(N5544), .A2(n26926), .ZN(N44992));
    INVX1 U32121 (.I(n28753), .ZN(N44993));
    INVX1 U32122 (.I(n20491), .ZN(N44994));
    INVX1 U32123 (.I(n43436), .ZN(N44995));
    NOR2X1 U32124 (.A1(n24350), .A2(n19883), .ZN(N44996));
    INVX1 U32125 (.I(N276), .ZN(N44997));
    NANDX1 U32126 (.A1(n28463), .A2(n27282), .ZN(N44998));
    NOR2X1 U32127 (.A1(N12200), .A2(n37064), .ZN(N44999));
    NOR2X1 U32128 (.A1(n13378), .A2(N1977), .ZN(N45000));
    NOR2X1 U32129 (.A1(n36369), .A2(N4826), .ZN(N45001));
    NANDX1 U32130 (.A1(n26628), .A2(n35421), .ZN(N45002));
    NANDX1 U32131 (.A1(n40113), .A2(n38058), .ZN(N45003));
    INVX1 U32132 (.I(n13246), .ZN(N45004));
    NOR2X1 U32133 (.A1(n32133), .A2(N6960), .ZN(N45005));
    NOR2X1 U32134 (.A1(N1065), .A2(N6923), .ZN(N45006));
    NANDX1 U32135 (.A1(n15094), .A2(n16485), .ZN(N45007));
    NOR2X1 U32136 (.A1(N5049), .A2(N4126), .ZN(N45008));
    INVX1 U32137 (.I(n22010), .ZN(N45009));
    NOR2X1 U32138 (.A1(N12040), .A2(n15601), .ZN(N45010));
    NANDX1 U32139 (.A1(n25417), .A2(N7258), .ZN(N45011));
    NANDX1 U32140 (.A1(n18313), .A2(N12083), .ZN(N45012));
    NOR2X1 U32141 (.A1(n34620), .A2(n37183), .ZN(N45013));
    NANDX1 U32142 (.A1(n20940), .A2(n21449), .ZN(N45014));
    NANDX1 U32143 (.A1(n23866), .A2(n25700), .ZN(N45015));
    NOR2X1 U32144 (.A1(n30825), .A2(n40122), .ZN(N45016));
    NANDX1 U32145 (.A1(n27427), .A2(N12092), .ZN(N45017));
    NANDX1 U32146 (.A1(N439), .A2(n37262), .ZN(N45018));
    NOR2X1 U32147 (.A1(N4565), .A2(n37102), .ZN(n45019));
    NOR2X1 U32148 (.A1(N8538), .A2(N5669), .ZN(N45020));
    INVX1 U32149 (.I(N7716), .ZN(N45021));
    NANDX1 U32150 (.A1(n19663), .A2(n37800), .ZN(N45022));
    NANDX1 U32151 (.A1(n21425), .A2(N11833), .ZN(N45023));
    NOR2X1 U32152 (.A1(n15135), .A2(n37495), .ZN(N45024));
    NOR2X1 U32153 (.A1(n26263), .A2(n23065), .ZN(N45025));
    NOR2X1 U32154 (.A1(N8491), .A2(N7615), .ZN(N45026));
    NOR2X1 U32155 (.A1(N5140), .A2(n16061), .ZN(N45027));
    NANDX1 U32156 (.A1(N6912), .A2(n39600), .ZN(N45028));
    INVX1 U32157 (.I(N701), .ZN(N45029));
    INVX1 U32158 (.I(n30697), .ZN(N45030));
    NANDX1 U32159 (.A1(n31839), .A2(n28914), .ZN(N45031));
    NOR2X1 U32160 (.A1(n33924), .A2(n26309), .ZN(N45032));
    NANDX1 U32161 (.A1(N10114), .A2(n20636), .ZN(N45033));
    NOR2X1 U32162 (.A1(n21218), .A2(n22148), .ZN(N45034));
    NANDX1 U32163 (.A1(n26033), .A2(N5850), .ZN(n45035));
    INVX1 U32164 (.I(N8823), .ZN(N45036));
    NANDX1 U32165 (.A1(n23915), .A2(N6993), .ZN(N45037));
    INVX1 U32166 (.I(n22182), .ZN(N45038));
    NOR2X1 U32167 (.A1(n42268), .A2(N4404), .ZN(N45039));
    INVX1 U32168 (.I(n38395), .ZN(N45040));
    NANDX1 U32169 (.A1(N9424), .A2(N9317), .ZN(N45041));
    NOR2X1 U32170 (.A1(n36905), .A2(n30835), .ZN(N45042));
    INVX1 U32171 (.I(n26582), .ZN(N45043));
    INVX1 U32172 (.I(N8869), .ZN(N45044));
    NOR2X1 U32173 (.A1(n21080), .A2(n19184), .ZN(N45045));
    NANDX1 U32174 (.A1(n42298), .A2(n31011), .ZN(N45046));
    NOR2X1 U32175 (.A1(n14538), .A2(n36860), .ZN(N45047));
    INVX1 U32176 (.I(n23360), .ZN(N45048));
    NANDX1 U32177 (.A1(n21176), .A2(n20033), .ZN(n45049));
    NANDX1 U32178 (.A1(n43358), .A2(n21845), .ZN(N45050));
    NOR2X1 U32179 (.A1(n37441), .A2(n30568), .ZN(N45051));
    NANDX1 U32180 (.A1(n24504), .A2(n29671), .ZN(N45052));
    INVX1 U32181 (.I(n21623), .ZN(N45053));
    INVX1 U32182 (.I(N7943), .ZN(N45054));
    NANDX1 U32183 (.A1(n39364), .A2(n18909), .ZN(N45055));
    NANDX1 U32184 (.A1(n32914), .A2(n39989), .ZN(N45056));
    NOR2X1 U32185 (.A1(N11869), .A2(n28494), .ZN(N45057));
    INVX1 U32186 (.I(n16772), .ZN(N45058));
    INVX1 U32187 (.I(n35991), .ZN(N45059));
    NOR2X1 U32188 (.A1(N12598), .A2(N4499), .ZN(N45060));
    INVX1 U32189 (.I(n32630), .ZN(N45061));
    NOR2X1 U32190 (.A1(n24774), .A2(N11002), .ZN(n45062));
    NOR2X1 U32191 (.A1(N8422), .A2(n31249), .ZN(N45063));
    INVX1 U32192 (.I(n22605), .ZN(N45064));
    NANDX1 U32193 (.A1(n37080), .A2(N755), .ZN(N45065));
    NANDX1 U32194 (.A1(n34702), .A2(n38089), .ZN(N45066));
    NOR2X1 U32195 (.A1(n43291), .A2(n40819), .ZN(N45067));
    INVX1 U32196 (.I(n39807), .ZN(N45068));
    NOR2X1 U32197 (.A1(N6789), .A2(n24828), .ZN(N45069));
    NOR2X1 U32198 (.A1(n13240), .A2(n14066), .ZN(N45070));
    NOR2X1 U32199 (.A1(n16953), .A2(n26663), .ZN(N45071));
    INVX1 U32200 (.I(n41841), .ZN(N45072));
    NANDX1 U32201 (.A1(n16812), .A2(N12822), .ZN(N45073));
    NANDX1 U32202 (.A1(n22047), .A2(n21243), .ZN(N45074));
    NOR2X1 U32203 (.A1(n28226), .A2(N375), .ZN(N45075));
    INVX1 U32204 (.I(N11513), .ZN(N45076));
    INVX1 U32205 (.I(n20994), .ZN(n45077));
    INVX1 U32206 (.I(n28897), .ZN(N45078));
    NOR2X1 U32207 (.A1(n35712), .A2(n26243), .ZN(N45079));
    INVX1 U32208 (.I(n32046), .ZN(N45080));
    INVX1 U32209 (.I(n17862), .ZN(N45081));
    NOR2X1 U32210 (.A1(n32932), .A2(n31102), .ZN(N45082));
    NOR2X1 U32211 (.A1(n23200), .A2(N4582), .ZN(n45083));
    NANDX1 U32212 (.A1(N7646), .A2(N2950), .ZN(N45084));
    NOR2X1 U32213 (.A1(n14137), .A2(n15771), .ZN(N45085));
    NANDX1 U32214 (.A1(n25863), .A2(n26693), .ZN(N45086));
    INVX1 U32215 (.I(N10616), .ZN(N45087));
    INVX1 U32216 (.I(n29893), .ZN(N45088));
    INVX1 U32217 (.I(n17875), .ZN(N45089));
    NOR2X1 U32218 (.A1(n14549), .A2(N3299), .ZN(N45090));
    NOR2X1 U32219 (.A1(n39941), .A2(n19221), .ZN(N45091));
    NOR2X1 U32220 (.A1(n28514), .A2(N610), .ZN(N45092));
    INVX1 U32221 (.I(n21275), .ZN(N45093));
    INVX1 U32222 (.I(n29810), .ZN(N45094));
    INVX1 U32223 (.I(N2948), .ZN(N45095));
    NANDX1 U32224 (.A1(n18116), .A2(N273), .ZN(N45096));
    NOR2X1 U32225 (.A1(N3312), .A2(n14409), .ZN(N45097));
    NANDX1 U32226 (.A1(N5010), .A2(n29951), .ZN(N45098));
    INVX1 U32227 (.I(n33817), .ZN(N45099));
    NOR2X1 U32228 (.A1(n32436), .A2(N9917), .ZN(N45100));
    INVX1 U32229 (.I(N6838), .ZN(N45101));
    INVX1 U32230 (.I(n13129), .ZN(N45102));
    INVX1 U32231 (.I(n20256), .ZN(N45103));
    NOR2X1 U32232 (.A1(n19036), .A2(N1102), .ZN(n45104));
    NOR2X1 U32233 (.A1(n19645), .A2(n43282), .ZN(N45105));
    INVX1 U32234 (.I(n42865), .ZN(N45106));
    NOR2X1 U32235 (.A1(n23372), .A2(N2340), .ZN(N45107));
    INVX1 U32236 (.I(n31168), .ZN(N45108));
    INVX1 U32237 (.I(n26916), .ZN(N45109));
    NANDX1 U32238 (.A1(N6700), .A2(n15913), .ZN(N45110));
    NANDX1 U32239 (.A1(n26330), .A2(n21282), .ZN(N45111));
    NANDX1 U32240 (.A1(n13103), .A2(N10245), .ZN(n45112));
    NOR2X1 U32241 (.A1(N11683), .A2(N6762), .ZN(N45113));
    NANDX1 U32242 (.A1(n14491), .A2(N6577), .ZN(N45114));
    NOR2X1 U32243 (.A1(n13768), .A2(n15292), .ZN(N45115));
    INVX1 U32244 (.I(n31238), .ZN(N45116));
    INVX1 U32245 (.I(n26645), .ZN(N45117));
    INVX1 U32246 (.I(n24008), .ZN(N45118));
    NOR2X1 U32247 (.A1(N6409), .A2(n16027), .ZN(N45119));
    NANDX1 U32248 (.A1(n27256), .A2(N8318), .ZN(N45120));
    NANDX1 U32249 (.A1(n18263), .A2(n15017), .ZN(N45121));
    NANDX1 U32250 (.A1(N3958), .A2(n41346), .ZN(N45122));
    INVX1 U32251 (.I(n23470), .ZN(N45123));
    INVX1 U32252 (.I(N12610), .ZN(N45124));
    NANDX1 U32253 (.A1(N12338), .A2(N9051), .ZN(N45125));
    NOR2X1 U32254 (.A1(n26829), .A2(n15628), .ZN(n45126));
    NANDX1 U32255 (.A1(n30276), .A2(n20599), .ZN(N45127));
    NANDX1 U32256 (.A1(n18041), .A2(N1743), .ZN(N45128));
    NANDX1 U32257 (.A1(N1078), .A2(n15430), .ZN(N45129));
    NANDX1 U32258 (.A1(n40638), .A2(n31457), .ZN(N45130));
    NOR2X1 U32259 (.A1(n24422), .A2(n39774), .ZN(N45131));
    NANDX1 U32260 (.A1(n32364), .A2(N999), .ZN(N45132));
    NOR2X1 U32261 (.A1(n36321), .A2(n32024), .ZN(N45133));
    INVX1 U32262 (.I(n16319), .ZN(n45134));
    NOR2X1 U32263 (.A1(n39541), .A2(n15425), .ZN(N45135));
    NANDX1 U32264 (.A1(N5119), .A2(n30329), .ZN(N45136));
    NANDX1 U32265 (.A1(n20746), .A2(N4662), .ZN(n45137));
    NANDX1 U32266 (.A1(n31025), .A2(n38981), .ZN(N45138));
    NANDX1 U32267 (.A1(n32767), .A2(n13001), .ZN(N45139));
    NOR2X1 U32268 (.A1(N4724), .A2(N12323), .ZN(n45140));
    NOR2X1 U32269 (.A1(n25860), .A2(N3692), .ZN(n45141));
    INVX1 U32270 (.I(n22162), .ZN(N45142));
    NANDX1 U32271 (.A1(n36643), .A2(N12840), .ZN(N45143));
    NANDX1 U32272 (.A1(n29491), .A2(N1391), .ZN(N45144));
    NANDX1 U32273 (.A1(n35489), .A2(n23750), .ZN(N45145));
    INVX1 U32274 (.I(n40593), .ZN(N45146));
    NOR2X1 U32275 (.A1(N403), .A2(n27449), .ZN(N45147));
    INVX1 U32276 (.I(N10829), .ZN(N45148));
    INVX1 U32277 (.I(N6923), .ZN(N45149));
    INVX1 U32278 (.I(n17299), .ZN(N45150));
    NOR2X1 U32279 (.A1(n20827), .A2(n19979), .ZN(N45151));
    NOR2X1 U32280 (.A1(n15230), .A2(n21981), .ZN(n45152));
    NOR2X1 U32281 (.A1(n41090), .A2(n25672), .ZN(N45153));
    NOR2X1 U32282 (.A1(N9459), .A2(n39694), .ZN(N45154));
    NANDX1 U32283 (.A1(n22298), .A2(N1659), .ZN(N45155));
    INVX1 U32284 (.I(n13368), .ZN(n45156));
    NANDX1 U32285 (.A1(n34157), .A2(n37118), .ZN(N45157));
    NOR2X1 U32286 (.A1(n20957), .A2(n41772), .ZN(N45158));
    NOR2X1 U32287 (.A1(n38086), .A2(n21006), .ZN(N45159));
    NANDX1 U32288 (.A1(N6083), .A2(n27928), .ZN(N45160));
    NANDX1 U32289 (.A1(n13061), .A2(n37106), .ZN(N45161));
    NOR2X1 U32290 (.A1(n33039), .A2(n39296), .ZN(N45162));
    NANDX1 U32291 (.A1(N1227), .A2(n21344), .ZN(N45163));
    NANDX1 U32292 (.A1(n26898), .A2(n17991), .ZN(N45164));
    NANDX1 U32293 (.A1(n23120), .A2(n30640), .ZN(N45165));
    INVX1 U32294 (.I(n14458), .ZN(N45166));
    NANDX1 U32295 (.A1(n24837), .A2(n38165), .ZN(N45167));
    INVX1 U32296 (.I(N8162), .ZN(N45168));
    NANDX1 U32297 (.A1(n20308), .A2(N6461), .ZN(N45169));
    INVX1 U32298 (.I(n14921), .ZN(N45170));
    NANDX1 U32299 (.A1(N11697), .A2(N10683), .ZN(N45171));
    INVX1 U32300 (.I(N9338), .ZN(N45172));
    INVX1 U32301 (.I(n28387), .ZN(N45173));
    INVX1 U32302 (.I(N2990), .ZN(N45174));
    NANDX1 U32303 (.A1(n20222), .A2(N4217), .ZN(N45175));
    NOR2X1 U32304 (.A1(N10255), .A2(n31114), .ZN(N45176));
    NANDX1 U32305 (.A1(N9747), .A2(N441), .ZN(n45177));
    INVX1 U32306 (.I(n21215), .ZN(N45178));
    INVX1 U32307 (.I(n15904), .ZN(N45179));
    INVX1 U32308 (.I(n32423), .ZN(N45180));
    INVX1 U32309 (.I(N420), .ZN(N45181));
    INVX1 U32310 (.I(n35562), .ZN(N45182));
    INVX1 U32311 (.I(n37901), .ZN(N45183));
    INVX1 U32312 (.I(n24026), .ZN(n45184));
    NANDX1 U32313 (.A1(N7372), .A2(n25627), .ZN(N45185));
    INVX1 U32314 (.I(n20795), .ZN(N45186));
    NOR2X1 U32315 (.A1(N12307), .A2(n23785), .ZN(N45187));
    INVX1 U32316 (.I(n22208), .ZN(N45188));
    NANDX1 U32317 (.A1(n16190), .A2(n32463), .ZN(N45189));
    NOR2X1 U32318 (.A1(n15620), .A2(n31889), .ZN(N45190));
    NANDX1 U32319 (.A1(n35369), .A2(N9631), .ZN(N45191));
    NOR2X1 U32320 (.A1(n40952), .A2(N1890), .ZN(N45192));
    NANDX1 U32321 (.A1(N12734), .A2(N2309), .ZN(N45193));
    NOR2X1 U32322 (.A1(n37975), .A2(n42341), .ZN(N45194));
    NANDX1 U32323 (.A1(n34664), .A2(n22894), .ZN(N45195));
    NANDX1 U32324 (.A1(n31716), .A2(n38200), .ZN(N45196));
    NANDX1 U32325 (.A1(N9038), .A2(n38420), .ZN(N45197));
    NOR2X1 U32326 (.A1(n22502), .A2(N9057), .ZN(N45198));
    NANDX1 U32327 (.A1(n40182), .A2(n14926), .ZN(N45199));
    NANDX1 U32328 (.A1(n35184), .A2(n20225), .ZN(N45200));
    NANDX1 U32329 (.A1(n20306), .A2(N12121), .ZN(N45201));
    NANDX1 U32330 (.A1(N10006), .A2(n42752), .ZN(N45202));
    NANDX1 U32331 (.A1(n21808), .A2(N12014), .ZN(N45203));
    INVX1 U32332 (.I(n25922), .ZN(n45204));
    INVX1 U32333 (.I(n15978), .ZN(N45205));
    INVX1 U32334 (.I(n30860), .ZN(N45206));
    NANDX1 U32335 (.A1(N8492), .A2(N8783), .ZN(n45207));
    INVX1 U32336 (.I(n41133), .ZN(N45208));
    INVX1 U32337 (.I(n18225), .ZN(N45209));
    NOR2X1 U32338 (.A1(n19682), .A2(n16961), .ZN(N45210));
    NANDX1 U32339 (.A1(n16391), .A2(n31886), .ZN(n45211));
    NOR2X1 U32340 (.A1(n41254), .A2(n41790), .ZN(N45212));
    INVX1 U32341 (.I(N7767), .ZN(N45213));
    NANDX1 U32342 (.A1(n41365), .A2(N7452), .ZN(N45214));
    NOR2X1 U32343 (.A1(n23013), .A2(n29259), .ZN(N45215));
    NOR2X1 U32344 (.A1(n40122), .A2(N1389), .ZN(N45216));
    NANDX1 U32345 (.A1(N12627), .A2(n15533), .ZN(N45217));
    NANDX1 U32346 (.A1(n41177), .A2(n13704), .ZN(n45218));
    NANDX1 U32347 (.A1(n20982), .A2(N11364), .ZN(N45219));
    NANDX1 U32348 (.A1(n28886), .A2(N179), .ZN(N45220));
    NOR2X1 U32349 (.A1(N2374), .A2(n35510), .ZN(N45221));
    NOR2X1 U32350 (.A1(n23939), .A2(n29721), .ZN(N45222));
    INVX1 U32351 (.I(n22256), .ZN(N45223));
    INVX1 U32352 (.I(N11614), .ZN(N45224));
    NOR2X1 U32353 (.A1(n35426), .A2(n19065), .ZN(N45225));
    NOR2X1 U32354 (.A1(n14966), .A2(n38004), .ZN(n45226));
    NOR2X1 U32355 (.A1(N1296), .A2(n39392), .ZN(N45227));
    NANDX1 U32356 (.A1(n13922), .A2(N1132), .ZN(N45228));
    INVX1 U32357 (.I(N11627), .ZN(N45229));
    NOR2X1 U32358 (.A1(n21102), .A2(n22288), .ZN(N45230));
    NOR2X1 U32359 (.A1(N1416), .A2(N7702), .ZN(N45231));
    INVX1 U32360 (.I(N11730), .ZN(N45232));
    INVX1 U32361 (.I(n41245), .ZN(N45233));
    INVX1 U32362 (.I(n34014), .ZN(N45234));
    NANDX1 U32363 (.A1(n21642), .A2(N2477), .ZN(N45235));
    NOR2X1 U32364 (.A1(n22935), .A2(n14530), .ZN(N45236));
    INVX1 U32365 (.I(n41999), .ZN(N45237));
    NANDX1 U32366 (.A1(N7833), .A2(n36530), .ZN(N45238));
    NANDX1 U32367 (.A1(N9128), .A2(n22129), .ZN(n45239));
    INVX1 U32368 (.I(n23050), .ZN(n45240));
    INVX1 U32369 (.I(n42836), .ZN(n45241));
    NOR2X1 U32370 (.A1(n17454), .A2(n20466), .ZN(N45242));
    NOR2X1 U32371 (.A1(n23011), .A2(n21881), .ZN(N45243));
    NANDX1 U32372 (.A1(n28747), .A2(n23290), .ZN(N45244));
    NOR2X1 U32373 (.A1(n16199), .A2(n30765), .ZN(N45245));
    NANDX1 U32374 (.A1(n23052), .A2(N8934), .ZN(N45246));
    NOR2X1 U32375 (.A1(n34286), .A2(n21548), .ZN(N45247));
    INVX1 U32376 (.I(n37473), .ZN(N45248));
    NOR2X1 U32377 (.A1(n23511), .A2(N1834), .ZN(N45249));
    INVX1 U32378 (.I(n18556), .ZN(N45250));
    NANDX1 U32379 (.A1(n14620), .A2(n23424), .ZN(N45251));
    INVX1 U32380 (.I(n27560), .ZN(N45252));
    NOR2X1 U32381 (.A1(n37725), .A2(N1541), .ZN(N45253));
    INVX1 U32382 (.I(n30576), .ZN(N45254));
    INVX1 U32383 (.I(N1020), .ZN(N45255));
    NOR2X1 U32384 (.A1(n42978), .A2(n13990), .ZN(N45256));
    NOR2X1 U32385 (.A1(n15704), .A2(N1282), .ZN(N45257));
    NANDX1 U32386 (.A1(n28436), .A2(n43367), .ZN(N45258));
    NANDX1 U32387 (.A1(n19249), .A2(n21442), .ZN(N45259));
    NANDX1 U32388 (.A1(N2930), .A2(n31195), .ZN(N45260));
    INVX1 U32389 (.I(N4763), .ZN(N45261));
    INVX1 U32390 (.I(n24242), .ZN(N45262));
    INVX1 U32391 (.I(n38306), .ZN(N45263));
    NOR2X1 U32392 (.A1(n18773), .A2(n22393), .ZN(n45264));
    NANDX1 U32393 (.A1(N2705), .A2(n13613), .ZN(n45265));
    INVX1 U32394 (.I(n33280), .ZN(n45266));
    INVX1 U32395 (.I(N7138), .ZN(N45267));
    NANDX1 U32396 (.A1(n37669), .A2(n21127), .ZN(n45268));
    NANDX1 U32397 (.A1(n43053), .A2(n22408), .ZN(N45269));
    INVX1 U32398 (.I(n28016), .ZN(N45270));
    NANDX1 U32399 (.A1(N5498), .A2(n36944), .ZN(N45271));
    NANDX1 U32400 (.A1(n41465), .A2(n39873), .ZN(N45272));
    NANDX1 U32401 (.A1(N3679), .A2(n34315), .ZN(N45273));
    NOR2X1 U32402 (.A1(n17600), .A2(n29398), .ZN(N45274));
    INVX1 U32403 (.I(n21792), .ZN(N45275));
    NOR2X1 U32404 (.A1(n41416), .A2(n38451), .ZN(N45276));
    INVX1 U32405 (.I(N1237), .ZN(N45277));
    NANDX1 U32406 (.A1(n30362), .A2(n39400), .ZN(N45278));
    INVX1 U32407 (.I(n40976), .ZN(N45279));
    NANDX1 U32408 (.A1(n19041), .A2(n39550), .ZN(N45280));
    NANDX1 U32409 (.A1(n41448), .A2(N6612), .ZN(N45281));
    NOR2X1 U32410 (.A1(N9958), .A2(N1789), .ZN(N45282));
    NANDX1 U32411 (.A1(n33060), .A2(n32934), .ZN(N45283));
    NANDX1 U32412 (.A1(N10733), .A2(n26292), .ZN(N45284));
    INVX1 U32413 (.I(n34924), .ZN(N45285));
    INVX1 U32414 (.I(n30023), .ZN(N45286));
    NOR2X1 U32415 (.A1(n22211), .A2(n24400), .ZN(N45287));
    NOR2X1 U32416 (.A1(N6869), .A2(n21482), .ZN(N45288));
    NOR2X1 U32417 (.A1(N7965), .A2(n41523), .ZN(N45289));
    INVX1 U32418 (.I(N5879), .ZN(N45290));
    NOR2X1 U32419 (.A1(N8218), .A2(n24919), .ZN(N45291));
    NOR2X1 U32420 (.A1(n20754), .A2(N12574), .ZN(N45292));
    NOR2X1 U32421 (.A1(N7513), .A2(N12211), .ZN(N45293));
    INVX1 U32422 (.I(n20896), .ZN(N45294));
    INVX1 U32423 (.I(N12324), .ZN(N45295));
    INVX1 U32424 (.I(N2211), .ZN(N45296));
    NANDX1 U32425 (.A1(n31304), .A2(n37134), .ZN(N45297));
    NANDX1 U32426 (.A1(n17855), .A2(N4137), .ZN(N45298));
    INVX1 U32427 (.I(n31934), .ZN(N45299));
    NANDX1 U32428 (.A1(n14322), .A2(N9943), .ZN(N45300));
    NANDX1 U32429 (.A1(N11966), .A2(N7993), .ZN(N45301));
    NOR2X1 U32430 (.A1(N7524), .A2(n36698), .ZN(n45302));
    NOR2X1 U32431 (.A1(n22122), .A2(n18009), .ZN(N45303));
    NOR2X1 U32432 (.A1(n34696), .A2(n39083), .ZN(N45304));
    INVX1 U32433 (.I(n36586), .ZN(N45305));
    INVX1 U32434 (.I(N417), .ZN(n45306));
    NANDX1 U32435 (.A1(n30797), .A2(n31095), .ZN(N45307));
    NOR2X1 U32436 (.A1(n25940), .A2(n18926), .ZN(N45308));
    INVX1 U32437 (.I(n21502), .ZN(N45309));
    NANDX1 U32438 (.A1(n28072), .A2(n18634), .ZN(N45310));
    NOR2X1 U32439 (.A1(n30306), .A2(n32955), .ZN(N45311));
    NANDX1 U32440 (.A1(n31874), .A2(n34601), .ZN(N45312));
    NOR2X1 U32441 (.A1(n28704), .A2(n42124), .ZN(N45313));
    NANDX1 U32442 (.A1(n23431), .A2(n20774), .ZN(N45314));
    INVX1 U32443 (.I(N5759), .ZN(n45315));
    NOR2X1 U32444 (.A1(N8740), .A2(n18432), .ZN(N45316));
    INVX1 U32445 (.I(n27213), .ZN(N45317));
    NOR2X1 U32446 (.A1(n22854), .A2(n14537), .ZN(N45318));
    INVX1 U32447 (.I(N9656), .ZN(N45319));
    NANDX1 U32448 (.A1(n15076), .A2(n33591), .ZN(N45320));
    NOR2X1 U32449 (.A1(n31215), .A2(N7871), .ZN(N45321));
    INVX1 U32450 (.I(N2664), .ZN(N45322));
    NANDX1 U32451 (.A1(N5981), .A2(N6888), .ZN(N45323));
    INVX1 U32452 (.I(n40581), .ZN(N45324));
    NOR2X1 U32453 (.A1(N1489), .A2(n39232), .ZN(N45325));
    INVX1 U32454 (.I(n24919), .ZN(N45326));
    NOR2X1 U32455 (.A1(n37675), .A2(n20357), .ZN(N45327));
    NANDX1 U32456 (.A1(N2942), .A2(n38789), .ZN(N45328));
    INVX1 U32457 (.I(n19834), .ZN(N45329));
    NANDX1 U32458 (.A1(n15212), .A2(n34370), .ZN(N45330));
    NOR2X1 U32459 (.A1(n24867), .A2(n21053), .ZN(N45331));
    NOR2X1 U32460 (.A1(N4665), .A2(n18917), .ZN(N45332));
    INVX1 U32461 (.I(N12535), .ZN(N45333));
    NANDX1 U32462 (.A1(n28307), .A2(n40391), .ZN(n45334));
    NOR2X1 U32463 (.A1(n35194), .A2(n13176), .ZN(N45335));
    NOR2X1 U32464 (.A1(N505), .A2(N4344), .ZN(N45336));
    INVX1 U32465 (.I(n14729), .ZN(N45337));
    NANDX1 U32466 (.A1(n19835), .A2(N8931), .ZN(N45338));
    NOR2X1 U32467 (.A1(n27723), .A2(N1553), .ZN(N45339));
    NANDX1 U32468 (.A1(n20081), .A2(N11066), .ZN(N45340));
    INVX1 U32469 (.I(n35292), .ZN(N45341));
    INVX1 U32470 (.I(N7491), .ZN(N45342));
    NOR2X1 U32471 (.A1(N12696), .A2(N1919), .ZN(N45343));
    NOR2X1 U32472 (.A1(n31613), .A2(n37881), .ZN(N45344));
    NANDX1 U32473 (.A1(n13235), .A2(N12395), .ZN(N45345));
    NANDX1 U32474 (.A1(N837), .A2(N4116), .ZN(N45346));
    INVX1 U32475 (.I(n29019), .ZN(N45347));
    NOR2X1 U32476 (.A1(n17361), .A2(n42640), .ZN(N45348));
    INVX1 U32477 (.I(n36302), .ZN(N45349));
    INVX1 U32478 (.I(N7639), .ZN(n45350));
    NOR2X1 U32479 (.A1(n36405), .A2(N9191), .ZN(n45351));
    INVX1 U32480 (.I(n13013), .ZN(N45352));
    NANDX1 U32481 (.A1(n43278), .A2(n37985), .ZN(N45353));
    NANDX1 U32482 (.A1(n40448), .A2(n34030), .ZN(N45354));
    NOR2X1 U32483 (.A1(n42366), .A2(N1588), .ZN(N45355));
    INVX1 U32484 (.I(n36775), .ZN(N45356));
    INVX1 U32485 (.I(N5329), .ZN(N45357));
    NANDX1 U32486 (.A1(n24995), .A2(N6165), .ZN(N45358));
    NOR2X1 U32487 (.A1(n38013), .A2(n35183), .ZN(N45359));
    NANDX1 U32488 (.A1(N1581), .A2(n24031), .ZN(N45360));
    NANDX1 U32489 (.A1(n37883), .A2(n43032), .ZN(N45361));
    NOR2X1 U32490 (.A1(N5898), .A2(n35964), .ZN(N45362));
    INVX1 U32491 (.I(n31358), .ZN(N45363));
    INVX1 U32492 (.I(N8945), .ZN(N45364));
    INVX1 U32493 (.I(n33169), .ZN(N45365));
    INVX1 U32494 (.I(n17819), .ZN(N45366));
    NOR2X1 U32495 (.A1(n24799), .A2(n16713), .ZN(N45367));
    NANDX1 U32496 (.A1(N6573), .A2(n43167), .ZN(n45368));
    NOR2X1 U32497 (.A1(N11902), .A2(n38543), .ZN(N45369));
    NANDX1 U32498 (.A1(N7746), .A2(n17395), .ZN(N45370));
    NANDX1 U32499 (.A1(n32609), .A2(N867), .ZN(n45371));
    NANDX1 U32500 (.A1(n13167), .A2(n36838), .ZN(N45372));
    NANDX1 U32501 (.A1(N2406), .A2(n36976), .ZN(N45373));
    NANDX1 U32502 (.A1(n38370), .A2(n35985), .ZN(N45374));
    NANDX1 U32503 (.A1(n23234), .A2(n34609), .ZN(N45375));
    NOR2X1 U32504 (.A1(N2610), .A2(N1661), .ZN(N45376));
    NOR2X1 U32505 (.A1(n16015), .A2(n16139), .ZN(N45377));
    NOR2X1 U32506 (.A1(n31008), .A2(n22711), .ZN(N45378));
    INVX1 U32507 (.I(N7041), .ZN(N45379));
    NOR2X1 U32508 (.A1(N6711), .A2(n41221), .ZN(N45380));
    INVX1 U32509 (.I(n24106), .ZN(N45381));
    NOR2X1 U32510 (.A1(n21174), .A2(n24972), .ZN(N45382));
    NANDX1 U32511 (.A1(n24020), .A2(n18337), .ZN(N45383));
    INVX1 U32512 (.I(n26425), .ZN(N45384));
    NANDX1 U32513 (.A1(N6693), .A2(N11002), .ZN(N45385));
    INVX1 U32514 (.I(n37698), .ZN(N45386));
    NANDX1 U32515 (.A1(n18321), .A2(N2601), .ZN(N45387));
    NOR2X1 U32516 (.A1(N9661), .A2(n18475), .ZN(N45388));
    NANDX1 U32517 (.A1(n25799), .A2(n40741), .ZN(N45389));
    INVX1 U32518 (.I(N5038), .ZN(N45390));
    INVX1 U32519 (.I(n26795), .ZN(N45391));
    NANDX1 U32520 (.A1(n25940), .A2(n14223), .ZN(n45392));
    NOR2X1 U32521 (.A1(N6573), .A2(n20050), .ZN(N45393));
    NANDX1 U32522 (.A1(n21224), .A2(N12706), .ZN(N45394));
    NANDX1 U32523 (.A1(n29240), .A2(N9431), .ZN(N45395));
    NOR2X1 U32524 (.A1(n20440), .A2(N5804), .ZN(N45396));
    NANDX1 U32525 (.A1(N4152), .A2(N29), .ZN(N45397));
    INVX1 U32526 (.I(N12153), .ZN(N45398));
    NOR2X1 U32527 (.A1(n22726), .A2(N11493), .ZN(N45399));
    NANDX1 U32528 (.A1(N11472), .A2(n37292), .ZN(n45400));
    NANDX1 U32529 (.A1(n31226), .A2(n32009), .ZN(n45401));
    INVX1 U32530 (.I(n14548), .ZN(N45402));
    NOR2X1 U32531 (.A1(n22260), .A2(n18450), .ZN(N45403));
    NOR2X1 U32532 (.A1(n18512), .A2(n38499), .ZN(n45404));
    NANDX1 U32533 (.A1(n39735), .A2(n40884), .ZN(N45405));
    NANDX1 U32534 (.A1(n15182), .A2(N6843), .ZN(N45406));
    NANDX1 U32535 (.A1(n35622), .A2(N2326), .ZN(N45407));
    NOR2X1 U32536 (.A1(n29453), .A2(n35506), .ZN(N45408));
    INVX1 U32537 (.I(n41605), .ZN(N45409));
    NOR2X1 U32538 (.A1(n30684), .A2(N9626), .ZN(N45410));
    INVX1 U32539 (.I(n42155), .ZN(N45411));
    NOR2X1 U32540 (.A1(N5369), .A2(n29908), .ZN(N45412));
    INVX1 U32541 (.I(N1689), .ZN(N45413));
    INVX1 U32542 (.I(n22357), .ZN(N45414));
    NOR2X1 U32543 (.A1(N9112), .A2(n27155), .ZN(N45415));
    NOR2X1 U32544 (.A1(n37291), .A2(N6908), .ZN(N45416));
    INVX1 U32545 (.I(n34702), .ZN(N45417));
    INVX1 U32546 (.I(N110), .ZN(N45418));
    NOR2X1 U32547 (.A1(n25102), .A2(n25411), .ZN(N45419));
    NOR2X1 U32548 (.A1(N3705), .A2(N11392), .ZN(N45420));
    NANDX1 U32549 (.A1(N11663), .A2(n42676), .ZN(N45421));
    NOR2X1 U32550 (.A1(n42346), .A2(n41981), .ZN(N45422));
    NOR2X1 U32551 (.A1(n30708), .A2(n35105), .ZN(N45423));
    INVX1 U32552 (.I(n17144), .ZN(N45424));
    INVX1 U32553 (.I(N3976), .ZN(N45425));
    NOR2X1 U32554 (.A1(n18482), .A2(n17603), .ZN(N45426));
    NOR2X1 U32555 (.A1(N2164), .A2(N6269), .ZN(N45427));
    INVX1 U32556 (.I(n42223), .ZN(n45428));
    NANDX1 U32557 (.A1(n24797), .A2(n40368), .ZN(N45429));
    NANDX1 U32558 (.A1(N12549), .A2(n21997), .ZN(N45430));
    NANDX1 U32559 (.A1(N2625), .A2(n15382), .ZN(N45431));
    INVX1 U32560 (.I(n17887), .ZN(n45432));
    NANDX1 U32561 (.A1(N6672), .A2(N7170), .ZN(N45433));
    NOR2X1 U32562 (.A1(N5180), .A2(N4089), .ZN(N45434));
    NANDX1 U32563 (.A1(n40285), .A2(n39529), .ZN(N45435));
    NOR2X1 U32564 (.A1(n36409), .A2(n33184), .ZN(N45436));
    NOR2X1 U32565 (.A1(N1098), .A2(N7315), .ZN(n45437));
    NOR2X1 U32566 (.A1(n36414), .A2(n13583), .ZN(N45438));
    INVX1 U32567 (.I(n35164), .ZN(N45439));
    NOR2X1 U32568 (.A1(n18309), .A2(n21740), .ZN(N45440));
    INVX1 U32569 (.I(n30857), .ZN(N45441));
    NOR2X1 U32570 (.A1(n14994), .A2(n23162), .ZN(N45442));
    INVX1 U32571 (.I(n22462), .ZN(N45443));
    NOR2X1 U32572 (.A1(n32368), .A2(n29133), .ZN(N45444));
    NANDX1 U32573 (.A1(N4492), .A2(n23992), .ZN(N45445));
    NOR2X1 U32574 (.A1(N7324), .A2(N10484), .ZN(n45446));
    INVX1 U32575 (.I(n16978), .ZN(N45447));
    NOR2X1 U32576 (.A1(N7113), .A2(n24118), .ZN(N45448));
    NOR2X1 U32577 (.A1(n14427), .A2(n27535), .ZN(N45449));
    NANDX1 U32578 (.A1(n17689), .A2(n21047), .ZN(N45450));
    NANDX1 U32579 (.A1(N12148), .A2(n39356), .ZN(N45451));
    NOR2X1 U32580 (.A1(n20745), .A2(n26740), .ZN(N45452));
    NANDX1 U32581 (.A1(n25419), .A2(N6429), .ZN(n45453));
    NOR2X1 U32582 (.A1(n37560), .A2(n26836), .ZN(n45454));
    NANDX1 U32583 (.A1(n23220), .A2(N10940), .ZN(n45455));
    NANDX1 U32584 (.A1(N3739), .A2(n32285), .ZN(n45456));
    NOR2X1 U32585 (.A1(n14223), .A2(N6213), .ZN(n45457));
    INVX1 U32586 (.I(N7323), .ZN(N45458));
    NOR2X1 U32587 (.A1(n29515), .A2(N1520), .ZN(N45459));
    NANDX1 U32588 (.A1(N3257), .A2(n32131), .ZN(N45460));
    INVX1 U32589 (.I(n24304), .ZN(N45461));
    NOR2X1 U32590 (.A1(n36947), .A2(n20187), .ZN(N45462));
    NANDX1 U32591 (.A1(N3900), .A2(n36606), .ZN(n45463));
    NOR2X1 U32592 (.A1(n18998), .A2(n32715), .ZN(N45464));
    NOR2X1 U32593 (.A1(n13085), .A2(n16078), .ZN(N45465));
    NANDX1 U32594 (.A1(n25984), .A2(n27018), .ZN(N45466));
    INVX1 U32595 (.I(n29722), .ZN(N45467));
    INVX1 U32596 (.I(n30943), .ZN(N45468));
    INVX1 U32597 (.I(N11722), .ZN(N45469));
    INVX1 U32598 (.I(n30626), .ZN(n45470));
    INVX1 U32599 (.I(N12061), .ZN(N45471));
    NOR2X1 U32600 (.A1(n32157), .A2(N4998), .ZN(N45472));
    INVX1 U32601 (.I(n13484), .ZN(N45473));
    INVX1 U32602 (.I(N11124), .ZN(N45474));
    INVX1 U32603 (.I(n39167), .ZN(N45475));
    INVX1 U32604 (.I(n33690), .ZN(N45476));
    NOR2X1 U32605 (.A1(N6246), .A2(N9215), .ZN(N45477));
    NOR2X1 U32606 (.A1(n39469), .A2(n22299), .ZN(N45478));
    NOR2X1 U32607 (.A1(n26464), .A2(n37962), .ZN(N45479));
    NANDX1 U32608 (.A1(n15195), .A2(n24211), .ZN(N45480));
    NOR2X1 U32609 (.A1(n35817), .A2(N4043), .ZN(N45481));
    NOR2X1 U32610 (.A1(n18363), .A2(n24348), .ZN(n45482));
    INVX1 U32611 (.I(n20104), .ZN(N45483));
    NOR2X1 U32612 (.A1(N10846), .A2(n25101), .ZN(N45484));
    INVX1 U32613 (.I(n24329), .ZN(N45485));
    NOR2X1 U32614 (.A1(n24307), .A2(n20967), .ZN(N45486));
    NANDX1 U32615 (.A1(n15999), .A2(N864), .ZN(N45487));
    NANDX1 U32616 (.A1(n22245), .A2(N10078), .ZN(N45488));
    NANDX1 U32617 (.A1(n18241), .A2(n22056), .ZN(N45489));
    NANDX1 U32618 (.A1(N1232), .A2(n16545), .ZN(N45490));
    NOR2X1 U32619 (.A1(N6106), .A2(n30436), .ZN(N45491));
    NOR2X1 U32620 (.A1(n31602), .A2(n24158), .ZN(N45492));
    NOR2X1 U32621 (.A1(n39644), .A2(N5033), .ZN(N45493));
    INVX1 U32622 (.I(N5955), .ZN(N45494));
    NOR2X1 U32623 (.A1(n39688), .A2(n20735), .ZN(N45495));
    NOR2X1 U32624 (.A1(n20544), .A2(n21343), .ZN(N45496));
    INVX1 U32625 (.I(n31191), .ZN(N45497));
    INVX1 U32626 (.I(N7430), .ZN(N45498));
    NANDX1 U32627 (.A1(n25607), .A2(n29674), .ZN(N45499));
    INVX1 U32628 (.I(N1318), .ZN(N45500));
    NOR2X1 U32629 (.A1(N10395), .A2(N4328), .ZN(N45501));
    INVX1 U32630 (.I(n16620), .ZN(N45502));
    NOR2X1 U32631 (.A1(n34610), .A2(N3583), .ZN(N45503));
    NOR2X1 U32632 (.A1(n22739), .A2(n27740), .ZN(N45504));
    NANDX1 U32633 (.A1(n18911), .A2(n22452), .ZN(N45505));
    NOR2X1 U32634 (.A1(n24865), .A2(n30185), .ZN(N45506));
    NANDX1 U32635 (.A1(N2128), .A2(n40782), .ZN(N45507));
    NOR2X1 U32636 (.A1(n13150), .A2(n32213), .ZN(N45508));
    INVX1 U32637 (.I(n20475), .ZN(N45509));
    NANDX1 U32638 (.A1(N4730), .A2(n35761), .ZN(n45510));
    INVX1 U32639 (.I(n36541), .ZN(N45511));
    NANDX1 U32640 (.A1(n19965), .A2(n36616), .ZN(n45512));
    INVX1 U32641 (.I(n15318), .ZN(N45513));
    NOR2X1 U32642 (.A1(n18306), .A2(n39607), .ZN(N45514));
    INVX1 U32643 (.I(N4774), .ZN(N45515));
    NOR2X1 U32644 (.A1(n30764), .A2(n31075), .ZN(N45516));
    NOR2X1 U32645 (.A1(N9743), .A2(N9595), .ZN(N45517));
    NOR2X1 U32646 (.A1(n29608), .A2(n27801), .ZN(N45518));
    NOR2X1 U32647 (.A1(n16597), .A2(N12759), .ZN(N45519));
    NANDX1 U32648 (.A1(N5337), .A2(n28907), .ZN(N45520));
    NANDX1 U32649 (.A1(n34658), .A2(n23317), .ZN(N45521));
    INVX1 U32650 (.I(n17029), .ZN(N45522));
    NANDX1 U32651 (.A1(n32692), .A2(n26674), .ZN(N45523));
    NANDX1 U32652 (.A1(N9984), .A2(n31671), .ZN(N45524));
    INVX1 U32653 (.I(n17969), .ZN(N45525));
    INVX1 U32654 (.I(n22314), .ZN(N45526));
    INVX1 U32655 (.I(N3206), .ZN(N45527));
    NANDX1 U32656 (.A1(N24), .A2(n20349), .ZN(n45528));
    NANDX1 U32657 (.A1(N9618), .A2(n18885), .ZN(n45529));
    NOR2X1 U32658 (.A1(n27099), .A2(N9227), .ZN(N45530));
    NANDX1 U32659 (.A1(n39857), .A2(N2399), .ZN(N45531));
    NOR2X1 U32660 (.A1(n25292), .A2(n16045), .ZN(N45532));
    NANDX1 U32661 (.A1(N5136), .A2(N11659), .ZN(N45533));
    NOR2X1 U32662 (.A1(N11200), .A2(n34030), .ZN(n45534));
    INVX1 U32663 (.I(N10408), .ZN(N45535));
    NANDX1 U32664 (.A1(N9220), .A2(n29697), .ZN(N45536));
    NANDX1 U32665 (.A1(n26704), .A2(N8539), .ZN(N45537));
    NANDX1 U32666 (.A1(n19590), .A2(N7823), .ZN(N45538));
    NANDX1 U32667 (.A1(n39938), .A2(N6530), .ZN(N45539));
    INVX1 U32668 (.I(n15350), .ZN(N45540));
    NOR2X1 U32669 (.A1(N3557), .A2(n14257), .ZN(N45541));
    NANDX1 U32670 (.A1(n33094), .A2(n16655), .ZN(N45542));
    INVX1 U32671 (.I(N4593), .ZN(N45543));
    INVX1 U32672 (.I(n43208), .ZN(N45544));
    INVX1 U32673 (.I(n34038), .ZN(N45545));
    NOR2X1 U32674 (.A1(N10607), .A2(n14276), .ZN(n45546));
    NOR2X1 U32675 (.A1(n21014), .A2(N4496), .ZN(N45547));
    INVX1 U32676 (.I(n40391), .ZN(N45548));
    INVX1 U32677 (.I(n40707), .ZN(N45549));
    NOR2X1 U32678 (.A1(N12654), .A2(n16824), .ZN(N45550));
    INVX1 U32679 (.I(n22967), .ZN(N45551));
    NOR2X1 U32680 (.A1(n42641), .A2(n32578), .ZN(N45552));
    INVX1 U32681 (.I(n34012), .ZN(N45553));
    NOR2X1 U32682 (.A1(n22255), .A2(N6182), .ZN(N45554));
    NANDX1 U32683 (.A1(n28590), .A2(n18277), .ZN(N45555));
    NOR2X1 U32684 (.A1(N7497), .A2(n18012), .ZN(N45556));
    NOR2X1 U32685 (.A1(n31214), .A2(N12095), .ZN(N45557));
    INVX1 U32686 (.I(N2017), .ZN(N45558));
    NANDX1 U32687 (.A1(n40734), .A2(n39665), .ZN(N45559));
    NOR2X1 U32688 (.A1(n37652), .A2(n31709), .ZN(n45560));
    NANDX1 U32689 (.A1(n22468), .A2(N890), .ZN(N45561));
    NOR2X1 U32690 (.A1(n25427), .A2(n13537), .ZN(N45562));
    NOR2X1 U32691 (.A1(n24595), .A2(N2642), .ZN(N45563));
    NANDX1 U32692 (.A1(N4814), .A2(n28455), .ZN(N45564));
    NOR2X1 U32693 (.A1(N675), .A2(N418), .ZN(n45565));
    NOR2X1 U32694 (.A1(n18952), .A2(n20444), .ZN(N45566));
    INVX1 U32695 (.I(n36963), .ZN(N45567));
    NANDX1 U32696 (.A1(n27557), .A2(n38738), .ZN(N45568));
    NOR2X1 U32697 (.A1(n19253), .A2(N12144), .ZN(N45569));
    INVX1 U32698 (.I(N5125), .ZN(N45570));
    NOR2X1 U32699 (.A1(n30399), .A2(n36833), .ZN(N45571));
    INVX1 U32700 (.I(N9394), .ZN(N45572));
    NOR2X1 U32701 (.A1(N10689), .A2(n24500), .ZN(N45573));
    NOR2X1 U32702 (.A1(n37958), .A2(n38774), .ZN(N45574));
    NOR2X1 U32703 (.A1(n29753), .A2(n33268), .ZN(N45575));
    NANDX1 U32704 (.A1(n33482), .A2(n33942), .ZN(N45576));
    INVX1 U32705 (.I(n32649), .ZN(N45577));
    NOR2X1 U32706 (.A1(n28783), .A2(n28991), .ZN(N45578));
    NANDX1 U32707 (.A1(N4548), .A2(N2755), .ZN(N45579));
    NANDX1 U32708 (.A1(N10353), .A2(N11688), .ZN(N45580));
    INVX1 U32709 (.I(n13419), .ZN(N45581));
    INVX1 U32710 (.I(N12065), .ZN(n45582));
    NOR2X1 U32711 (.A1(n43325), .A2(n41926), .ZN(n45583));
    INVX1 U32712 (.I(n27255), .ZN(N45584));
    NANDX1 U32713 (.A1(n13598), .A2(n14401), .ZN(N45585));
    NOR2X1 U32714 (.A1(n42052), .A2(N4188), .ZN(N45586));
    INVX1 U32715 (.I(n31847), .ZN(N45587));
    NANDX1 U32716 (.A1(N2749), .A2(n22316), .ZN(N45588));
    NOR2X1 U32717 (.A1(n35397), .A2(n21417), .ZN(N45589));
    NANDX1 U32718 (.A1(N10596), .A2(n14008), .ZN(N45590));
    NANDX1 U32719 (.A1(N3030), .A2(n35016), .ZN(n45591));
    INVX1 U32720 (.I(n14717), .ZN(N45592));
    NANDX1 U32721 (.A1(n13435), .A2(n21209), .ZN(N45593));
    NOR2X1 U32722 (.A1(N3460), .A2(n21061), .ZN(n45594));
    NOR2X1 U32723 (.A1(n25710), .A2(n37995), .ZN(N45595));
    NANDX1 U32724 (.A1(n39307), .A2(n42075), .ZN(n45596));
    INVX1 U32725 (.I(n37886), .ZN(N45597));
    NOR2X1 U32726 (.A1(n29761), .A2(n15940), .ZN(n45598));
    NANDX1 U32727 (.A1(n32510), .A2(n38256), .ZN(N45599));
    INVX1 U32728 (.I(n14114), .ZN(N45600));
    NANDX1 U32729 (.A1(n20462), .A2(n24709), .ZN(N45601));
    INVX1 U32730 (.I(N10126), .ZN(N45602));
    NOR2X1 U32731 (.A1(N11430), .A2(N10142), .ZN(N45603));
    INVX1 U32732 (.I(n25804), .ZN(n45604));
    NOR2X1 U32733 (.A1(N9871), .A2(N8771), .ZN(N45605));
    INVX1 U32734 (.I(n20611), .ZN(N45606));
    NOR2X1 U32735 (.A1(n42425), .A2(n15133), .ZN(N45607));
    NANDX1 U32736 (.A1(n27939), .A2(n13735), .ZN(N45608));
    NOR2X1 U32737 (.A1(N12033), .A2(N6204), .ZN(N45609));
    INVX1 U32738 (.I(n27972), .ZN(N45610));
    INVX1 U32739 (.I(n29085), .ZN(N45611));
    NOR2X1 U32740 (.A1(n25486), .A2(n43199), .ZN(N45612));
    INVX1 U32741 (.I(n35628), .ZN(N45613));
    NOR2X1 U32742 (.A1(n27880), .A2(N2281), .ZN(N45614));
    NANDX1 U32743 (.A1(n39309), .A2(N12423), .ZN(N45615));
    NOR2X1 U32744 (.A1(N11321), .A2(n25679), .ZN(N45616));
    INVX1 U32745 (.I(n20091), .ZN(N45617));
    INVX1 U32746 (.I(n30037), .ZN(N45618));
    INVX1 U32747 (.I(n41346), .ZN(N45619));
    INVX1 U32748 (.I(N3548), .ZN(N45620));
    NOR2X1 U32749 (.A1(N5112), .A2(n13835), .ZN(N45621));
    INVX1 U32750 (.I(N995), .ZN(N45622));
    INVX1 U32751 (.I(N12024), .ZN(N45623));
    NOR2X1 U32752 (.A1(n39495), .A2(n24458), .ZN(n45624));
    NANDX1 U32753 (.A1(n39221), .A2(n42772), .ZN(N45625));
    NOR2X1 U32754 (.A1(n43015), .A2(n16859), .ZN(n45626));
    NANDX1 U32755 (.A1(n31076), .A2(N2376), .ZN(N45627));
    NOR2X1 U32756 (.A1(n40951), .A2(n13696), .ZN(N45628));
    NOR2X1 U32757 (.A1(N6904), .A2(n23466), .ZN(N45629));
    NOR2X1 U32758 (.A1(n36940), .A2(n23428), .ZN(N45630));
    NANDX1 U32759 (.A1(n28317), .A2(n16655), .ZN(N45631));
    NOR2X1 U32760 (.A1(n23108), .A2(n30489), .ZN(n45632));
    INVX1 U32761 (.I(n13782), .ZN(N45633));
    INVX1 U32762 (.I(n36877), .ZN(N45634));
    INVX1 U32763 (.I(n26600), .ZN(N45635));
    NOR2X1 U32764 (.A1(n42179), .A2(N12028), .ZN(N45636));
    NANDX1 U32765 (.A1(N7483), .A2(N11571), .ZN(N45637));
    NOR2X1 U32766 (.A1(N8219), .A2(n32326), .ZN(N45638));
    INVX1 U32767 (.I(n21378), .ZN(N45639));
    NANDX1 U32768 (.A1(n29450), .A2(N6422), .ZN(N45640));
    INVX1 U32769 (.I(N9444), .ZN(N45641));
    INVX1 U32770 (.I(n19855), .ZN(N45642));
    NOR2X1 U32771 (.A1(n15698), .A2(N4699), .ZN(N45643));
    NANDX1 U32772 (.A1(N2708), .A2(n17486), .ZN(n45644));
    NOR2X1 U32773 (.A1(n27562), .A2(n31267), .ZN(n45645));
    NOR2X1 U32774 (.A1(n20966), .A2(N3032), .ZN(N45646));
    NOR2X1 U32775 (.A1(n28508), .A2(n34890), .ZN(N45647));
    INVX1 U32776 (.I(n25029), .ZN(N45648));
    INVX1 U32777 (.I(n42883), .ZN(N45649));
    INVX1 U32778 (.I(n40271), .ZN(N45650));
    NANDX1 U32779 (.A1(N10691), .A2(N7856), .ZN(n45651));
    INVX1 U32780 (.I(n29821), .ZN(N45652));
    NOR2X1 U32781 (.A1(n34134), .A2(n28944), .ZN(N45653));
    INVX1 U32782 (.I(N10516), .ZN(N45654));
    NOR2X1 U32783 (.A1(N10042), .A2(N4894), .ZN(N45655));
    INVX1 U32784 (.I(N12749), .ZN(N45656));
    NANDX1 U32785 (.A1(n32166), .A2(n40310), .ZN(N45657));
    NANDX1 U32786 (.A1(n24851), .A2(N7484), .ZN(N45658));
    NOR2X1 U32787 (.A1(n33816), .A2(n25671), .ZN(N45659));
    NANDX1 U32788 (.A1(n21657), .A2(N7228), .ZN(N45660));
    NOR2X1 U32789 (.A1(N10747), .A2(n35316), .ZN(N45661));
    NANDX1 U32790 (.A1(n32163), .A2(n35686), .ZN(N45662));
    NANDX1 U32791 (.A1(n39909), .A2(n22034), .ZN(N45663));
    INVX1 U32792 (.I(n20250), .ZN(N45664));
    INVX1 U32793 (.I(n41819), .ZN(N45665));
    INVX1 U32794 (.I(n38358), .ZN(N45666));
    INVX1 U32795 (.I(n25338), .ZN(N45667));
    INVX1 U32796 (.I(N10816), .ZN(n45668));
    NOR2X1 U32797 (.A1(n32996), .A2(N7654), .ZN(N45669));
    NANDX1 U32798 (.A1(n14375), .A2(N4817), .ZN(n45670));
    INVX1 U32799 (.I(n37870), .ZN(N45671));
    NOR2X1 U32800 (.A1(N3474), .A2(n16054), .ZN(n45672));
    INVX1 U32801 (.I(n42339), .ZN(N45673));
    NANDX1 U32802 (.A1(n19237), .A2(n24210), .ZN(N45674));
    INVX1 U32803 (.I(N11451), .ZN(n45675));
    NANDX1 U32804 (.A1(n34759), .A2(n23164), .ZN(N45676));
    INVX1 U32805 (.I(N11537), .ZN(N45677));
    INVX1 U32806 (.I(N5965), .ZN(N45678));
    NANDX1 U32807 (.A1(N4914), .A2(N4032), .ZN(N45679));
    NOR2X1 U32808 (.A1(n16065), .A2(N4527), .ZN(N45680));
    NANDX1 U32809 (.A1(N5588), .A2(N12180), .ZN(N45681));
    INVX1 U32810 (.I(N9642), .ZN(N45682));
    NOR2X1 U32811 (.A1(N10718), .A2(N4040), .ZN(N45683));
    NOR2X1 U32812 (.A1(n14192), .A2(N9773), .ZN(n45684));
    INVX1 U32813 (.I(N2738), .ZN(N45685));
    NOR2X1 U32814 (.A1(n30001), .A2(n26948), .ZN(N45686));
    NOR2X1 U32815 (.A1(n41451), .A2(n40883), .ZN(N45687));
    NANDX1 U32816 (.A1(N10822), .A2(N5029), .ZN(N45688));
    NANDX1 U32817 (.A1(n31170), .A2(N673), .ZN(N45689));
    NOR2X1 U32818 (.A1(n36084), .A2(n37856), .ZN(N45690));
    NOR2X1 U32819 (.A1(n41828), .A2(n42383), .ZN(N45691));
    NOR2X1 U32820 (.A1(n37095), .A2(N770), .ZN(N45692));
    NOR2X1 U32821 (.A1(n36417), .A2(N7446), .ZN(N45693));
    NANDX1 U32822 (.A1(n30136), .A2(n34288), .ZN(N45694));
    NOR2X1 U32823 (.A1(n39908), .A2(N1579), .ZN(N45695));
    NOR2X1 U32824 (.A1(N12369), .A2(n21259), .ZN(N45696));
    NOR2X1 U32825 (.A1(n33471), .A2(N8917), .ZN(N45697));
    NOR2X1 U32826 (.A1(N2388), .A2(n19739), .ZN(N45698));
    INVX1 U32827 (.I(n26313), .ZN(N45699));
    INVX1 U32828 (.I(n21060), .ZN(n45700));
    INVX1 U32829 (.I(n33199), .ZN(N45701));
    NOR2X1 U32830 (.A1(N914), .A2(n21234), .ZN(N45702));
    NOR2X1 U32831 (.A1(N4003), .A2(N4537), .ZN(N45703));
    NANDX1 U32832 (.A1(N8638), .A2(n40953), .ZN(n45704));
    INVX1 U32833 (.I(n13670), .ZN(N45705));
    INVX1 U32834 (.I(n25895), .ZN(N45706));
    NANDX1 U32835 (.A1(n13731), .A2(n27473), .ZN(N45707));
    INVX1 U32836 (.I(n15779), .ZN(N45708));
    NOR2X1 U32837 (.A1(n29329), .A2(N5778), .ZN(N45709));
    NOR2X1 U32838 (.A1(N11535), .A2(N8165), .ZN(N45710));
    NOR2X1 U32839 (.A1(n31921), .A2(n24158), .ZN(N45711));
    NANDX1 U32840 (.A1(n42660), .A2(N9112), .ZN(N45712));
    NANDX1 U32841 (.A1(N4311), .A2(n43177), .ZN(N45713));
    NOR2X1 U32842 (.A1(N8343), .A2(N3708), .ZN(N45714));
    NANDX1 U32843 (.A1(N2825), .A2(N2025), .ZN(n45715));
    NOR2X1 U32844 (.A1(N4752), .A2(n15694), .ZN(N45716));
    INVX1 U32845 (.I(n30646), .ZN(N45717));
    NOR2X1 U32846 (.A1(n23431), .A2(N4327), .ZN(N45718));
    INVX1 U32847 (.I(n39210), .ZN(N45719));
    NANDX1 U32848 (.A1(n37694), .A2(N1515), .ZN(N45720));
    INVX1 U32849 (.I(n38908), .ZN(N45721));
    NOR2X1 U32850 (.A1(n26715), .A2(n27357), .ZN(N45722));
    NOR2X1 U32851 (.A1(n37104), .A2(n16224), .ZN(N45723));
    INVX1 U32852 (.I(n37219), .ZN(N45724));
    INVX1 U32853 (.I(n22012), .ZN(N45725));
    INVX1 U32854 (.I(n28877), .ZN(N45726));
    NOR2X1 U32855 (.A1(n20341), .A2(n21381), .ZN(N45727));
    NOR2X1 U32856 (.A1(n23066), .A2(n15813), .ZN(N45728));
    INVX1 U32857 (.I(n43086), .ZN(N45729));
    NANDX1 U32858 (.A1(n17589), .A2(n23045), .ZN(N45730));
    INVX1 U32859 (.I(n25954), .ZN(n45731));
    NANDX1 U32860 (.A1(n29409), .A2(n20176), .ZN(N45732));
    INVX1 U32861 (.I(n32530), .ZN(N45733));
    NANDX1 U32862 (.A1(n42486), .A2(N5452), .ZN(n45734));
    NANDX1 U32863 (.A1(n22530), .A2(n42555), .ZN(N45735));
    INVX1 U32864 (.I(n34516), .ZN(N45736));
    INVX1 U32865 (.I(n15612), .ZN(N45737));
    NOR2X1 U32866 (.A1(n30757), .A2(n34168), .ZN(n45738));
    NANDX1 U32867 (.A1(N7625), .A2(N12077), .ZN(N45739));
    NANDX1 U32868 (.A1(n20371), .A2(n27889), .ZN(N45740));
    NANDX1 U32869 (.A1(n19984), .A2(n20554), .ZN(N45741));
    NOR2X1 U32870 (.A1(n32708), .A2(n17546), .ZN(N45742));
    NANDX1 U32871 (.A1(n41169), .A2(N3482), .ZN(N45743));
    NOR2X1 U32872 (.A1(n40824), .A2(n25691), .ZN(N45744));
    INVX1 U32873 (.I(n29518), .ZN(N45745));
    INVX1 U32874 (.I(n19268), .ZN(N45746));
    NOR2X1 U32875 (.A1(n19904), .A2(n24666), .ZN(N45747));
    NANDX1 U32876 (.A1(N2413), .A2(n40277), .ZN(N45748));
    NANDX1 U32877 (.A1(n33169), .A2(n30973), .ZN(N45749));
    INVX1 U32878 (.I(n30473), .ZN(N45750));
    INVX1 U32879 (.I(N12568), .ZN(N45751));
    NOR2X1 U32880 (.A1(n17145), .A2(n27445), .ZN(N45752));
    NOR2X1 U32881 (.A1(n27378), .A2(N6119), .ZN(N45753));
    INVX1 U32882 (.I(n34603), .ZN(N45754));
    INVX1 U32883 (.I(n37119), .ZN(n45755));
    INVX1 U32884 (.I(N2396), .ZN(N45756));
    NOR2X1 U32885 (.A1(N9983), .A2(n32488), .ZN(N45757));
    NANDX1 U32886 (.A1(n30805), .A2(N8283), .ZN(N45758));
    NANDX1 U32887 (.A1(n40388), .A2(n22628), .ZN(N45759));
    INVX1 U32888 (.I(n42800), .ZN(N45760));
    NANDX1 U32889 (.A1(n33251), .A2(n22176), .ZN(N45761));
    NOR2X1 U32890 (.A1(n43415), .A2(n42329), .ZN(N45762));
    NOR2X1 U32891 (.A1(N12510), .A2(N6227), .ZN(N45763));
    NANDX1 U32892 (.A1(n29635), .A2(n12941), .ZN(N45764));
    INVX1 U32893 (.I(n35753), .ZN(N45765));
    INVX1 U32894 (.I(N881), .ZN(N45766));
    NOR2X1 U32895 (.A1(n35689), .A2(n18325), .ZN(n45767));
    NOR2X1 U32896 (.A1(n16366), .A2(n28307), .ZN(N45768));
    NOR2X1 U32897 (.A1(n26561), .A2(N5319), .ZN(N45769));
    INVX1 U32898 (.I(n24689), .ZN(N45770));
    INVX1 U32899 (.I(N4706), .ZN(N45771));
    NOR2X1 U32900 (.A1(n34714), .A2(n13818), .ZN(N45772));
    NOR2X1 U32901 (.A1(N3098), .A2(N110), .ZN(N45773));
    INVX1 U32902 (.I(N1954), .ZN(N45774));
    NANDX1 U32903 (.A1(N4025), .A2(n41332), .ZN(N45775));
    NOR2X1 U32904 (.A1(n23339), .A2(N481), .ZN(N45776));
    NANDX1 U32905 (.A1(n15619), .A2(N9371), .ZN(n45777));
    NANDX1 U32906 (.A1(n18644), .A2(N1587), .ZN(N45778));
    NANDX1 U32907 (.A1(N3424), .A2(n17952), .ZN(N45779));
    INVX1 U32908 (.I(n31012), .ZN(N45780));
    NANDX1 U32909 (.A1(n33121), .A2(n13090), .ZN(n45781));
    NOR2X1 U32910 (.A1(n25035), .A2(n17795), .ZN(N45782));
    NOR2X1 U32911 (.A1(N5956), .A2(n31613), .ZN(N45783));
    NOR2X1 U32912 (.A1(n42205), .A2(n31722), .ZN(N45784));
    NOR2X1 U32913 (.A1(n33838), .A2(n40532), .ZN(n45785));
    INVX1 U32914 (.I(n21378), .ZN(N45786));
    NOR2X1 U32915 (.A1(n37974), .A2(n21858), .ZN(N45787));
    NANDX1 U32916 (.A1(n43272), .A2(n31228), .ZN(n45788));
    NOR2X1 U32917 (.A1(N8124), .A2(n22494), .ZN(N45789));
    NANDX1 U32918 (.A1(N11547), .A2(n30125), .ZN(N45790));
    NOR2X1 U32919 (.A1(n42558), .A2(n20845), .ZN(N45791));
    NOR2X1 U32920 (.A1(N12175), .A2(n25933), .ZN(N45792));
    NOR2X1 U32921 (.A1(n19650), .A2(n32815), .ZN(N45793));
    NOR2X1 U32922 (.A1(N7790), .A2(N8438), .ZN(n45794));
    INVX1 U32923 (.I(n29191), .ZN(N45795));
    NANDX1 U32924 (.A1(n19887), .A2(n26250), .ZN(N45796));
    NOR2X1 U32925 (.A1(n41264), .A2(n24811), .ZN(N45797));
    NANDX1 U32926 (.A1(N9329), .A2(N3662), .ZN(N45798));
    NANDX1 U32927 (.A1(n40556), .A2(n17477), .ZN(N45799));
    INVX1 U32928 (.I(N9257), .ZN(N45800));
    NOR2X1 U32929 (.A1(n37333), .A2(n39382), .ZN(N45801));
    NOR2X1 U32930 (.A1(n26098), .A2(n16754), .ZN(N45802));
    NANDX1 U32931 (.A1(n38273), .A2(n32366), .ZN(N45803));
    NANDX1 U32932 (.A1(N4130), .A2(n21708), .ZN(N45804));
    NOR2X1 U32933 (.A1(N11919), .A2(n19826), .ZN(N45805));
    NOR2X1 U32934 (.A1(n41109), .A2(n38873), .ZN(N45806));
    INVX1 U32935 (.I(n23887), .ZN(N45807));
    NOR2X1 U32936 (.A1(n41909), .A2(n38377), .ZN(N45808));
    INVX1 U32937 (.I(N7765), .ZN(N45809));
    NANDX1 U32938 (.A1(N10817), .A2(n38001), .ZN(N45810));
    NOR2X1 U32939 (.A1(n26282), .A2(N3785), .ZN(N45811));
    INVX1 U32940 (.I(n20142), .ZN(N45812));
    NOR2X1 U32941 (.A1(n31780), .A2(N2768), .ZN(N45813));
    NOR2X1 U32942 (.A1(N4020), .A2(n30720), .ZN(N45814));
    NOR2X1 U32943 (.A1(n21732), .A2(n24529), .ZN(N45815));
    NOR2X1 U32944 (.A1(n26761), .A2(n36447), .ZN(N45816));
    INVX1 U32945 (.I(N7519), .ZN(N45817));
    INVX1 U32946 (.I(N993), .ZN(N45818));
    INVX1 U32947 (.I(n37329), .ZN(N45819));
    INVX1 U32948 (.I(N6600), .ZN(N45820));
    INVX1 U32949 (.I(N2589), .ZN(N45821));
    INVX1 U32950 (.I(n43311), .ZN(N45822));
    NANDX1 U32951 (.A1(n42044), .A2(N5560), .ZN(N45823));
    NOR2X1 U32952 (.A1(n35509), .A2(n42067), .ZN(N45824));
    INVX1 U32953 (.I(n35202), .ZN(N45825));
    INVX1 U32954 (.I(n31635), .ZN(N45826));
    INVX1 U32955 (.I(n24074), .ZN(N45827));
    INVX1 U32956 (.I(N5388), .ZN(N45828));
    INVX1 U32957 (.I(n33090), .ZN(N45829));
    NOR2X1 U32958 (.A1(N8454), .A2(n15744), .ZN(N45830));
    INVX1 U32959 (.I(n15972), .ZN(N45831));
    NANDX1 U32960 (.A1(N8060), .A2(n24135), .ZN(n45832));
    NANDX1 U32961 (.A1(n27815), .A2(n30734), .ZN(N45833));
    INVX1 U32962 (.I(n30403), .ZN(N45834));
    NANDX1 U32963 (.A1(n34474), .A2(n33488), .ZN(N45835));
    INVX1 U32964 (.I(n40033), .ZN(N45836));
    NANDX1 U32965 (.A1(n15065), .A2(n28308), .ZN(N45837));
    NANDX1 U32966 (.A1(n39947), .A2(n38042), .ZN(N45838));
    NANDX1 U32967 (.A1(n27483), .A2(N8323), .ZN(N45839));
    NANDX1 U32968 (.A1(n32870), .A2(N335), .ZN(N45840));
    NOR2X1 U32969 (.A1(n24025), .A2(n41940), .ZN(N45841));
    NOR2X1 U32970 (.A1(n31091), .A2(N4120), .ZN(N45842));
    INVX1 U32971 (.I(n39150), .ZN(N45843));
    NANDX1 U32972 (.A1(N5299), .A2(n13172), .ZN(N45844));
    NOR2X1 U32973 (.A1(n39934), .A2(n33255), .ZN(N45845));
    NANDX1 U32974 (.A1(n20615), .A2(n12950), .ZN(N45846));
    NANDX1 U32975 (.A1(N6855), .A2(n22011), .ZN(N45847));
    INVX1 U32976 (.I(n35162), .ZN(N45848));
    NANDX1 U32977 (.A1(N108), .A2(n19411), .ZN(N45849));
    INVX1 U32978 (.I(n17270), .ZN(N45850));
    NANDX1 U32979 (.A1(N587), .A2(n39819), .ZN(N45851));
    NANDX1 U32980 (.A1(n24857), .A2(n20371), .ZN(N45852));
    NOR2X1 U32981 (.A1(n21398), .A2(n41142), .ZN(N45853));
    NANDX1 U32982 (.A1(N3654), .A2(n36819), .ZN(N45854));
    NANDX1 U32983 (.A1(N8952), .A2(N6519), .ZN(N45855));
    INVX1 U32984 (.I(n38565), .ZN(N45856));
    INVX1 U32985 (.I(n31835), .ZN(N45857));
    NOR2X1 U32986 (.A1(n42402), .A2(n30723), .ZN(N45858));
    INVX1 U32987 (.I(n20940), .ZN(N45859));
    NOR2X1 U32988 (.A1(N3931), .A2(n37406), .ZN(N45860));
    NANDX1 U32989 (.A1(n23341), .A2(N3340), .ZN(N45861));
    NANDX1 U32990 (.A1(n40754), .A2(N3926), .ZN(N45862));
    NOR2X1 U32991 (.A1(n15029), .A2(n28782), .ZN(N45863));
    INVX1 U32992 (.I(n20923), .ZN(n45864));
    INVX1 U32993 (.I(N2006), .ZN(N45865));
    INVX1 U32994 (.I(N40), .ZN(N45866));
    INVX1 U32995 (.I(n38244), .ZN(N45867));
    NANDX1 U32996 (.A1(n24703), .A2(n40426), .ZN(N45868));
    INVX1 U32997 (.I(N10683), .ZN(N45869));
    INVX1 U32998 (.I(n42621), .ZN(N45870));
    NOR2X1 U32999 (.A1(N5718), .A2(N11390), .ZN(N45871));
    NANDX1 U33000 (.A1(n29754), .A2(N5000), .ZN(N45872));
    NOR2X1 U33001 (.A1(N10424), .A2(n18020), .ZN(N45873));
    NOR2X1 U33002 (.A1(n41516), .A2(n15301), .ZN(N45874));
    NANDX1 U33003 (.A1(n25482), .A2(n20009), .ZN(N45875));
    INVX1 U33004 (.I(n19498), .ZN(N45876));
    INVX1 U33005 (.I(n25956), .ZN(N45877));
    INVX1 U33006 (.I(N7756), .ZN(N45878));
    NOR2X1 U33007 (.A1(n39688), .A2(n35679), .ZN(N45879));
    NOR2X1 U33008 (.A1(n20918), .A2(n32632), .ZN(N45880));
    NOR2X1 U33009 (.A1(n21280), .A2(n17947), .ZN(N45881));
    INVX1 U33010 (.I(n30891), .ZN(N45882));
    INVX1 U33011 (.I(n41478), .ZN(N45883));
    NOR2X1 U33012 (.A1(n43097), .A2(n36157), .ZN(N45884));
    NOR2X1 U33013 (.A1(n43201), .A2(N10704), .ZN(N45885));
    NOR2X1 U33014 (.A1(n30924), .A2(n15685), .ZN(N45886));
    NANDX1 U33015 (.A1(N2613), .A2(n35693), .ZN(N45887));
    INVX1 U33016 (.I(n22110), .ZN(N45888));
    INVX1 U33017 (.I(n19002), .ZN(N45889));
    NANDX1 U33018 (.A1(n30587), .A2(n34676), .ZN(N45890));
    NANDX1 U33019 (.A1(n22793), .A2(N5549), .ZN(N45891));
    NOR2X1 U33020 (.A1(N11952), .A2(N3337), .ZN(N45892));
    NANDX1 U33021 (.A1(n19578), .A2(n33425), .ZN(N45893));
    NOR2X1 U33022 (.A1(n32922), .A2(n21110), .ZN(N45894));
    NANDX1 U33023 (.A1(n22226), .A2(n13794), .ZN(N45895));
    NOR2X1 U33024 (.A1(N11634), .A2(n24497), .ZN(N45896));
    NOR2X1 U33025 (.A1(n42557), .A2(n29861), .ZN(N45897));
    NANDX1 U33026 (.A1(n34849), .A2(n22082), .ZN(N45898));
    NANDX1 U33027 (.A1(n13487), .A2(N1441), .ZN(N45899));
    NANDX1 U33028 (.A1(n36459), .A2(n21708), .ZN(n45900));
    NANDX1 U33029 (.A1(N1855), .A2(N1028), .ZN(N45901));
    INVX1 U33030 (.I(n21319), .ZN(N45902));
    INVX1 U33031 (.I(N10628), .ZN(N45903));
    NOR2X1 U33032 (.A1(N11917), .A2(n33732), .ZN(N45904));
    NANDX1 U33033 (.A1(n34518), .A2(N11369), .ZN(N45905));
    NANDX1 U33034 (.A1(N2952), .A2(n25162), .ZN(N45906));
    INVX1 U33035 (.I(n14585), .ZN(N45907));
    NOR2X1 U33036 (.A1(n13822), .A2(N3350), .ZN(N45908));
    NOR2X1 U33037 (.A1(n32954), .A2(n38198), .ZN(N45909));
    INVX1 U33038 (.I(n34813), .ZN(N45910));
    NANDX1 U33039 (.A1(n38929), .A2(N12200), .ZN(N45911));
    INVX1 U33040 (.I(N6844), .ZN(N45912));
    NANDX1 U33041 (.A1(n15565), .A2(N7871), .ZN(N45913));
    NOR2X1 U33042 (.A1(n36883), .A2(N210), .ZN(N45914));
    NANDX1 U33043 (.A1(N1681), .A2(N12127), .ZN(N45915));
    NOR2X1 U33044 (.A1(n27793), .A2(n36324), .ZN(N45916));
    NOR2X1 U33045 (.A1(n35922), .A2(n39275), .ZN(N45917));
    NOR2X1 U33046 (.A1(n27240), .A2(N10388), .ZN(N45918));
    NOR2X1 U33047 (.A1(n41061), .A2(N3417), .ZN(N45919));
    NOR2X1 U33048 (.A1(n30542), .A2(n41614), .ZN(N45920));
    INVX1 U33049 (.I(N11562), .ZN(N45921));
    NOR2X1 U33050 (.A1(n18116), .A2(n23762), .ZN(N45922));
    NOR2X1 U33051 (.A1(n24959), .A2(n37704), .ZN(N45923));
    NANDX1 U33052 (.A1(n22509), .A2(N5146), .ZN(N45924));
    INVX1 U33053 (.I(N12399), .ZN(N45925));
    INVX1 U33054 (.I(n43231), .ZN(N45926));
    INVX1 U33055 (.I(n28169), .ZN(N45927));
    INVX1 U33056 (.I(N7056), .ZN(N45928));
    NOR2X1 U33057 (.A1(N9680), .A2(N2859), .ZN(N45929));
    NOR2X1 U33058 (.A1(n36919), .A2(N2926), .ZN(N45930));
    NOR2X1 U33059 (.A1(n24187), .A2(N6342), .ZN(N45931));
    INVX1 U33060 (.I(N936), .ZN(N45932));
    NANDX1 U33061 (.A1(n23473), .A2(N12498), .ZN(N45933));
    INVX1 U33062 (.I(n31268), .ZN(N45934));
    NANDX1 U33063 (.A1(n22771), .A2(N2434), .ZN(N45935));
    INVX1 U33064 (.I(n27438), .ZN(N45936));
    NANDX1 U33065 (.A1(n14996), .A2(n25516), .ZN(n45937));
    NANDX1 U33066 (.A1(n41683), .A2(n25274), .ZN(N45938));
    NANDX1 U33067 (.A1(n26379), .A2(n42504), .ZN(N45939));
    INVX1 U33068 (.I(n23924), .ZN(N45940));
    INVX1 U33069 (.I(n40818), .ZN(N45941));
    NANDX1 U33070 (.A1(N2157), .A2(N271), .ZN(N45942));
    NANDX1 U33071 (.A1(n16023), .A2(n39764), .ZN(n45943));
    NANDX1 U33072 (.A1(n16958), .A2(n33926), .ZN(N45944));
    NOR2X1 U33073 (.A1(n29455), .A2(N3482), .ZN(N45945));
    NOR2X1 U33074 (.A1(N11921), .A2(n15932), .ZN(N45946));
    NANDX1 U33075 (.A1(n21771), .A2(n43370), .ZN(N45947));
    NANDX1 U33076 (.A1(n36766), .A2(n15093), .ZN(N45948));
    NOR2X1 U33077 (.A1(n34976), .A2(n40366), .ZN(N45949));
    NOR2X1 U33078 (.A1(N7562), .A2(n39397), .ZN(N45950));
    NOR2X1 U33079 (.A1(n21165), .A2(n37787), .ZN(N45951));
    NOR2X1 U33080 (.A1(n26853), .A2(n39943), .ZN(N45952));
    INVX1 U33081 (.I(n27543), .ZN(N45953));
    NANDX1 U33082 (.A1(N12029), .A2(N8405), .ZN(N45954));
    INVX1 U33083 (.I(n35634), .ZN(N45955));
    NOR2X1 U33084 (.A1(n38265), .A2(n39115), .ZN(N45956));
    NANDX1 U33085 (.A1(N6713), .A2(N1255), .ZN(N45957));
    NANDX1 U33086 (.A1(n28483), .A2(n34304), .ZN(N45958));
    INVX1 U33087 (.I(n21776), .ZN(n45959));
    INVX1 U33088 (.I(n13859), .ZN(N45960));
    NOR2X1 U33089 (.A1(N2817), .A2(n37494), .ZN(N45961));
    NOR2X1 U33090 (.A1(n31893), .A2(n22464), .ZN(N45962));
    INVX1 U33091 (.I(n26207), .ZN(N45963));
    NANDX1 U33092 (.A1(n37897), .A2(N12357), .ZN(N45964));
    NANDX1 U33093 (.A1(N11647), .A2(n14529), .ZN(N45965));
    NANDX1 U33094 (.A1(n20052), .A2(n23338), .ZN(N45966));
    NOR2X1 U33095 (.A1(n32791), .A2(n18130), .ZN(N45967));
    NOR2X1 U33096 (.A1(n27339), .A2(n14523), .ZN(N45968));
    INVX1 U33097 (.I(N6130), .ZN(N45969));
    NOR2X1 U33098 (.A1(n14625), .A2(n37577), .ZN(n45970));
    NANDX1 U33099 (.A1(n20548), .A2(n41116), .ZN(N45971));
    INVX1 U33100 (.I(n13044), .ZN(N45972));
    NANDX1 U33101 (.A1(n36979), .A2(N1464), .ZN(N45973));
    NANDX1 U33102 (.A1(N4551), .A2(n17350), .ZN(N45974));
    INVX1 U33103 (.I(n42447), .ZN(N45975));
    NANDX1 U33104 (.A1(n41615), .A2(N302), .ZN(N45976));
    NANDX1 U33105 (.A1(n43198), .A2(N10033), .ZN(n45977));
    NOR2X1 U33106 (.A1(N3791), .A2(n32503), .ZN(n45978));
    NOR2X1 U33107 (.A1(n26331), .A2(n16369), .ZN(N45979));
    NOR2X1 U33108 (.A1(N6652), .A2(N12179), .ZN(N45980));
    NOR2X1 U33109 (.A1(n21277), .A2(n39435), .ZN(N45981));
    INVX1 U33110 (.I(n41824), .ZN(n45982));
    NANDX1 U33111 (.A1(n42130), .A2(N11396), .ZN(N45983));
    INVX1 U33112 (.I(n35636), .ZN(N45984));
    NOR2X1 U33113 (.A1(n32551), .A2(n40186), .ZN(N45985));
    INVX1 U33114 (.I(n20497), .ZN(N45986));
    NANDX1 U33115 (.A1(n28954), .A2(N8319), .ZN(N45987));
    NANDX1 U33116 (.A1(n42228), .A2(n41197), .ZN(N45988));
    INVX1 U33117 (.I(n35367), .ZN(N45989));
    NOR2X1 U33118 (.A1(n17884), .A2(N3163), .ZN(N45990));
    INVX1 U33119 (.I(n23932), .ZN(N45991));
    INVX1 U33120 (.I(n24177), .ZN(N45992));
    NOR2X1 U33121 (.A1(n23317), .A2(N1981), .ZN(N45993));
    NOR2X1 U33122 (.A1(n18348), .A2(n33484), .ZN(N45994));
    INVX1 U33123 (.I(n17005), .ZN(N45995));
    INVX1 U33124 (.I(N628), .ZN(N45996));
    NOR2X1 U33125 (.A1(n37098), .A2(n22858), .ZN(N45997));
    INVX1 U33126 (.I(N3194), .ZN(n45998));
    NOR2X1 U33127 (.A1(n14082), .A2(n21827), .ZN(N45999));
    NANDX1 U33128 (.A1(n32903), .A2(n20582), .ZN(N46000));
    INVX1 U33129 (.I(n18284), .ZN(n46001));
    NOR2X1 U33130 (.A1(n19952), .A2(n36167), .ZN(N46002));
    NANDX1 U33131 (.A1(n37476), .A2(N6307), .ZN(N46003));
    NANDX1 U33132 (.A1(N7860), .A2(n42416), .ZN(N46004));
    NANDX1 U33133 (.A1(n42992), .A2(n20696), .ZN(N46005));
    NANDX1 U33134 (.A1(n33004), .A2(n36054), .ZN(N46006));
    INVX1 U33135 (.I(n24090), .ZN(N46007));
    NANDX1 U33136 (.A1(n17355), .A2(n17715), .ZN(N46008));
    NOR2X1 U33137 (.A1(N2597), .A2(N10588), .ZN(n46009));
    NOR2X1 U33138 (.A1(n16678), .A2(n32415), .ZN(n46010));
    NANDX1 U33139 (.A1(N6109), .A2(n42676), .ZN(N46011));
    NOR2X1 U33140 (.A1(n14072), .A2(N1360), .ZN(N46012));
    NOR2X1 U33141 (.A1(n39919), .A2(N6678), .ZN(N46013));
    INVX1 U33142 (.I(N2753), .ZN(N46014));
    INVX1 U33143 (.I(n33440), .ZN(N46015));
    INVX1 U33144 (.I(N3464), .ZN(N46016));
    NANDX1 U33145 (.A1(N12072), .A2(n15286), .ZN(N46017));
    NOR2X1 U33146 (.A1(n37805), .A2(n23472), .ZN(N46018));
    INVX1 U33147 (.I(n31013), .ZN(N46019));
    NANDX1 U33148 (.A1(N10502), .A2(N3607), .ZN(N46020));
    NOR2X1 U33149 (.A1(N10770), .A2(n42387), .ZN(N46021));
    INVX1 U33150 (.I(n32864), .ZN(N46022));
    NOR2X1 U33151 (.A1(N2096), .A2(n32067), .ZN(N46023));
    NANDX1 U33152 (.A1(n16168), .A2(n33426), .ZN(N46024));
    NANDX1 U33153 (.A1(N12614), .A2(n29783), .ZN(N46025));
    NANDX1 U33154 (.A1(N5046), .A2(N6619), .ZN(N46026));
    NANDX1 U33155 (.A1(n39893), .A2(N10082), .ZN(N46027));
    INVX1 U33156 (.I(n41644), .ZN(N46028));
    INVX1 U33157 (.I(N9035), .ZN(N46029));
    INVX1 U33158 (.I(n38519), .ZN(N46030));
    INVX1 U33159 (.I(n13197), .ZN(N46031));
    NANDX1 U33160 (.A1(N2004), .A2(N6483), .ZN(N46032));
    NANDX1 U33161 (.A1(N12773), .A2(N5398), .ZN(n46033));
    NANDX1 U33162 (.A1(n35316), .A2(n30653), .ZN(N46034));
    INVX1 U33163 (.I(n23910), .ZN(N46035));
    INVX1 U33164 (.I(n29433), .ZN(N46036));
    NANDX1 U33165 (.A1(n36533), .A2(n31726), .ZN(N46037));
    NANDX1 U33166 (.A1(n20792), .A2(n26451), .ZN(N46038));
    NOR2X1 U33167 (.A1(n28171), .A2(N12551), .ZN(N46039));
    NOR2X1 U33168 (.A1(n14716), .A2(N10723), .ZN(N46040));
    INVX1 U33169 (.I(n13430), .ZN(N46041));
    NOR2X1 U33170 (.A1(N6327), .A2(N4932), .ZN(N46042));
    NOR2X1 U33171 (.A1(n21559), .A2(n40087), .ZN(N46043));
    NOR2X1 U33172 (.A1(n36741), .A2(n42539), .ZN(N46044));
    NANDX1 U33173 (.A1(N4438), .A2(n34382), .ZN(N46045));
    INVX1 U33174 (.I(n17703), .ZN(n46046));
    NOR2X1 U33175 (.A1(n29222), .A2(n36815), .ZN(N46047));
    NANDX1 U33176 (.A1(N11962), .A2(n14748), .ZN(N46048));
    INVX1 U33177 (.I(n32753), .ZN(N46049));
    NOR2X1 U33178 (.A1(n27520), .A2(N7131), .ZN(n46050));
    INVX1 U33179 (.I(n23753), .ZN(N46051));
    NOR2X1 U33180 (.A1(N10679), .A2(n24713), .ZN(N46052));
    NANDX1 U33181 (.A1(n36736), .A2(n20719), .ZN(N46053));
    NOR2X1 U33182 (.A1(n32518), .A2(n42277), .ZN(N46054));
    NOR2X1 U33183 (.A1(n34782), .A2(n25225), .ZN(n46055));
    INVX1 U33184 (.I(n32123), .ZN(N46056));
    INVX1 U33185 (.I(N6156), .ZN(N46057));
    NOR2X1 U33186 (.A1(n37045), .A2(N10654), .ZN(N46058));
    NANDX1 U33187 (.A1(n30388), .A2(n18696), .ZN(N46059));
    NOR2X1 U33188 (.A1(N1663), .A2(N6271), .ZN(N46060));
    INVX1 U33189 (.I(n32541), .ZN(N46061));
    NOR2X1 U33190 (.A1(n33597), .A2(n32497), .ZN(n46062));
    NOR2X1 U33191 (.A1(n34802), .A2(n32855), .ZN(N46063));
    INVX1 U33192 (.I(n16285), .ZN(N46064));
    NOR2X1 U33193 (.A1(n38861), .A2(n25531), .ZN(N46065));
    NOR2X1 U33194 (.A1(n27346), .A2(n41711), .ZN(N46066));
    NOR2X1 U33195 (.A1(N9098), .A2(n13485), .ZN(N46067));
    INVX1 U33196 (.I(n38760), .ZN(N46068));
    NANDX1 U33197 (.A1(N1445), .A2(n22013), .ZN(N46069));
    NANDX1 U33198 (.A1(n36989), .A2(N8928), .ZN(N46070));
    NANDX1 U33199 (.A1(n30702), .A2(N270), .ZN(N46071));
    INVX1 U33200 (.I(n24016), .ZN(N46072));
    NOR2X1 U33201 (.A1(n14616), .A2(N3820), .ZN(N46073));
    NOR2X1 U33202 (.A1(n41197), .A2(n38621), .ZN(N46074));
    NOR2X1 U33203 (.A1(n15867), .A2(N1114), .ZN(N46075));
    INVX1 U33204 (.I(N936), .ZN(n46076));
    INVX1 U33205 (.I(n31856), .ZN(N46077));
    NANDX1 U33206 (.A1(n24883), .A2(n17688), .ZN(N46078));
    NOR2X1 U33207 (.A1(n28047), .A2(n35641), .ZN(N46079));
    NOR2X1 U33208 (.A1(n37367), .A2(n37086), .ZN(N46080));
    NANDX1 U33209 (.A1(n13868), .A2(n20282), .ZN(N46081));
    NOR2X1 U33210 (.A1(n42216), .A2(N7512), .ZN(N46082));
    NOR2X1 U33211 (.A1(n23042), .A2(n21207), .ZN(n46083));
    NOR2X1 U33212 (.A1(n37657), .A2(n14706), .ZN(n46084));
    NANDX1 U33213 (.A1(n25061), .A2(N9854), .ZN(N46085));
    NOR2X1 U33214 (.A1(n40928), .A2(N647), .ZN(N46086));
    NOR2X1 U33215 (.A1(n41863), .A2(n27291), .ZN(N46087));
    NOR2X1 U33216 (.A1(n16351), .A2(n41853), .ZN(n46088));
    NOR2X1 U33217 (.A1(N10256), .A2(n26427), .ZN(N46089));
    NANDX1 U33218 (.A1(n22281), .A2(n20321), .ZN(N46090));
    INVX1 U33219 (.I(N12846), .ZN(N46091));
    INVX1 U33220 (.I(N11887), .ZN(N46092));
    NOR2X1 U33221 (.A1(n22611), .A2(N9078), .ZN(N46093));
    NOR2X1 U33222 (.A1(N2180), .A2(n19964), .ZN(N46094));
    NANDX1 U33223 (.A1(n29516), .A2(n34669), .ZN(N46095));
    INVX1 U33224 (.I(N11105), .ZN(N46096));
    INVX1 U33225 (.I(n30535), .ZN(N46097));
    NOR2X1 U33226 (.A1(n24529), .A2(n17776), .ZN(N46098));
    INVX1 U33227 (.I(N8347), .ZN(N46099));
    INVX1 U33228 (.I(N2660), .ZN(N46100));
    INVX1 U33229 (.I(n32376), .ZN(N46101));
    NANDX1 U33230 (.A1(N12514), .A2(N7536), .ZN(N46102));
    NANDX1 U33231 (.A1(n22514), .A2(n42613), .ZN(N46103));
    NANDX1 U33232 (.A1(N2910), .A2(N708), .ZN(N46104));
    NOR2X1 U33233 (.A1(n15200), .A2(n42937), .ZN(N46105));
    NOR2X1 U33234 (.A1(N7060), .A2(n19429), .ZN(N46106));
    INVX1 U33235 (.I(n26255), .ZN(N46107));
    INVX1 U33236 (.I(N7630), .ZN(N46108));
    NANDX1 U33237 (.A1(n24187), .A2(n27845), .ZN(N46109));
    NANDX1 U33238 (.A1(N5244), .A2(N2148), .ZN(N46110));
    NANDX1 U33239 (.A1(n13590), .A2(N8060), .ZN(N46111));
    INVX1 U33240 (.I(n43149), .ZN(N46112));
    NANDX1 U33241 (.A1(n39673), .A2(N12190), .ZN(N46113));
    INVX1 U33242 (.I(N10756), .ZN(N46114));
    NOR2X1 U33243 (.A1(n36792), .A2(n27836), .ZN(N46115));
    INVX1 U33244 (.I(n27179), .ZN(N46116));
    NOR2X1 U33245 (.A1(n32172), .A2(n26643), .ZN(N46117));
    NANDX1 U33246 (.A1(n39231), .A2(N2599), .ZN(N46118));
    NOR2X1 U33247 (.A1(N11693), .A2(n36056), .ZN(n46119));
    NOR2X1 U33248 (.A1(n38732), .A2(n16770), .ZN(n46120));
    NOR2X1 U33249 (.A1(N10217), .A2(n22013), .ZN(N46121));
    NOR2X1 U33250 (.A1(N1164), .A2(n25283), .ZN(N46122));
    INVX1 U33251 (.I(n38241), .ZN(N46123));
    NANDX1 U33252 (.A1(n37458), .A2(n34441), .ZN(N46124));
    NOR2X1 U33253 (.A1(n31636), .A2(n34876), .ZN(N46125));
    NOR2X1 U33254 (.A1(n14635), .A2(n19240), .ZN(N46126));
    INVX1 U33255 (.I(n31493), .ZN(N46127));
    INVX1 U33256 (.I(n23729), .ZN(N46128));
    NOR2X1 U33257 (.A1(n13888), .A2(N9167), .ZN(N46129));
    NANDX1 U33258 (.A1(n19021), .A2(n20859), .ZN(n46130));
    NANDX1 U33259 (.A1(n31784), .A2(N5798), .ZN(N46131));
    INVX1 U33260 (.I(n18599), .ZN(N46132));
    NOR2X1 U33261 (.A1(n27987), .A2(N7562), .ZN(N46133));
    NANDX1 U33262 (.A1(N9797), .A2(N4584), .ZN(N46134));
    NANDX1 U33263 (.A1(n34755), .A2(n31721), .ZN(N46135));
    INVX1 U33264 (.I(N7790), .ZN(N46136));
    NOR2X1 U33265 (.A1(N6830), .A2(n15528), .ZN(N46137));
    INVX1 U33266 (.I(n15749), .ZN(n46138));
    NANDX1 U33267 (.A1(N1899), .A2(n38450), .ZN(N46139));
    NANDX1 U33268 (.A1(N6242), .A2(n42017), .ZN(N46140));
    NANDX1 U33269 (.A1(n13184), .A2(n17565), .ZN(N46141));
    INVX1 U33270 (.I(N2388), .ZN(N46142));
    NANDX1 U33271 (.A1(N2523), .A2(N8362), .ZN(N46143));
    NOR2X1 U33272 (.A1(N8217), .A2(n36349), .ZN(N46144));
    NANDX1 U33273 (.A1(n15074), .A2(N2673), .ZN(N46145));
    NOR2X1 U33274 (.A1(N6379), .A2(n27108), .ZN(N46146));
    INVX1 U33275 (.I(n21805), .ZN(N46147));
    INVX1 U33276 (.I(N3471), .ZN(N46148));
    NANDX1 U33277 (.A1(N6952), .A2(N7029), .ZN(N46149));
    NOR2X1 U33278 (.A1(N3716), .A2(n42079), .ZN(N46150));
    NOR2X1 U33279 (.A1(n24208), .A2(N4849), .ZN(N46151));
    NANDX1 U33280 (.A1(N74), .A2(N7712), .ZN(N46152));
    NANDX1 U33281 (.A1(N7119), .A2(n43251), .ZN(N46153));
    INVX1 U33282 (.I(n42793), .ZN(N46154));
    INVX1 U33283 (.I(n34219), .ZN(N46155));
    NANDX1 U33284 (.A1(n34169), .A2(N2143), .ZN(N46156));
    NOR2X1 U33285 (.A1(n36841), .A2(N7801), .ZN(N46157));
    NOR2X1 U33286 (.A1(N10156), .A2(N1708), .ZN(N46158));
    INVX1 U33287 (.I(n34733), .ZN(N46159));
    INVX1 U33288 (.I(N4995), .ZN(N46160));
    INVX1 U33289 (.I(n35038), .ZN(N46161));
    NOR2X1 U33290 (.A1(n35080), .A2(n33644), .ZN(N46162));
    NOR2X1 U33291 (.A1(N5495), .A2(n28172), .ZN(N46163));
    NANDX1 U33292 (.A1(N5569), .A2(n35883), .ZN(N46164));
    NOR2X1 U33293 (.A1(N2367), .A2(n35662), .ZN(n46165));
    NOR2X1 U33294 (.A1(N1687), .A2(n33482), .ZN(N46166));
    INVX1 U33295 (.I(n42375), .ZN(N46167));
    NOR2X1 U33296 (.A1(n25557), .A2(N872), .ZN(N46168));
    NOR2X1 U33297 (.A1(n33357), .A2(N9219), .ZN(N46169));
    INVX1 U33298 (.I(n24744), .ZN(N46170));
    NANDX1 U33299 (.A1(n41794), .A2(N9281), .ZN(N46171));
    INVX1 U33300 (.I(n19365), .ZN(N46172));
    NANDX1 U33301 (.A1(n29630), .A2(N652), .ZN(N46173));
    NOR2X1 U33302 (.A1(N462), .A2(N6147), .ZN(N46174));
    NOR2X1 U33303 (.A1(n42349), .A2(N1395), .ZN(N46175));
    NOR2X1 U33304 (.A1(n21801), .A2(n36913), .ZN(N46176));
    NANDX1 U33305 (.A1(n31636), .A2(n28279), .ZN(N46177));
    INVX1 U33306 (.I(N11578), .ZN(N46178));
    INVX1 U33307 (.I(n20167), .ZN(N46179));
    NANDX1 U33308 (.A1(n28052), .A2(n27392), .ZN(N46180));
    INVX1 U33309 (.I(n37270), .ZN(N46181));
    NOR2X1 U33310 (.A1(n41442), .A2(n22849), .ZN(N46182));
    NANDX1 U33311 (.A1(n40403), .A2(N3101), .ZN(N46183));
    NANDX1 U33312 (.A1(n30928), .A2(n22410), .ZN(N46184));
    NOR2X1 U33313 (.A1(N1305), .A2(n22871), .ZN(N46185));
    NOR2X1 U33314 (.A1(n43326), .A2(n21748), .ZN(N46186));
    INVX1 U33315 (.I(n23965), .ZN(N46187));
    NANDX1 U33316 (.A1(n33130), .A2(n40265), .ZN(N46188));
    INVX1 U33317 (.I(n17936), .ZN(n46189));
    INVX1 U33318 (.I(n22649), .ZN(N46190));
    NOR2X1 U33319 (.A1(N2628), .A2(N5990), .ZN(N46191));
    INVX1 U33320 (.I(n30019), .ZN(N46192));
    NOR2X1 U33321 (.A1(N2853), .A2(N10680), .ZN(N46193));
    NANDX1 U33322 (.A1(n15381), .A2(n22813), .ZN(N46194));
    NANDX1 U33323 (.A1(N8161), .A2(n21159), .ZN(N46195));
    INVX1 U33324 (.I(n30571), .ZN(N46196));
    NOR2X1 U33325 (.A1(n29180), .A2(N9969), .ZN(N46197));
    NANDX1 U33326 (.A1(n18713), .A2(n21396), .ZN(N46198));
    INVX1 U33327 (.I(n42677), .ZN(n46199));
    NOR2X1 U33328 (.A1(n13367), .A2(n29149), .ZN(N46200));
    INVX1 U33329 (.I(n20983), .ZN(N46201));
    INVX1 U33330 (.I(N1398), .ZN(N46202));
    NOR2X1 U33331 (.A1(n14237), .A2(N7387), .ZN(N46203));
    NANDX1 U33332 (.A1(N783), .A2(n19755), .ZN(N46204));
    NOR2X1 U33333 (.A1(N1142), .A2(n30092), .ZN(N46205));
    NANDX1 U33334 (.A1(n23955), .A2(n27039), .ZN(N46206));
    NANDX1 U33335 (.A1(n34793), .A2(N11441), .ZN(N46207));
    NANDX1 U33336 (.A1(N1157), .A2(n30300), .ZN(N46208));
    NANDX1 U33337 (.A1(n38969), .A2(n38692), .ZN(N46209));
    INVX1 U33338 (.I(n29526), .ZN(N46210));
    NANDX1 U33339 (.A1(N2934), .A2(n32572), .ZN(N46211));
    NANDX1 U33340 (.A1(n14835), .A2(N10082), .ZN(N46212));
    NANDX1 U33341 (.A1(n16232), .A2(n22388), .ZN(N46213));
    NOR2X1 U33342 (.A1(n13298), .A2(n33428), .ZN(N46214));
    NOR2X1 U33343 (.A1(n33052), .A2(N3848), .ZN(N46215));
    NOR2X1 U33344 (.A1(N9351), .A2(n22800), .ZN(N46216));
    NANDX1 U33345 (.A1(n36389), .A2(N6440), .ZN(N46217));
    NOR2X1 U33346 (.A1(n37510), .A2(n20651), .ZN(N46218));
    NOR2X1 U33347 (.A1(n24337), .A2(n34510), .ZN(N46219));
    NANDX1 U33348 (.A1(n19557), .A2(n15972), .ZN(N46220));
    NANDX1 U33349 (.A1(N3660), .A2(n18905), .ZN(N46221));
    NOR2X1 U33350 (.A1(n16912), .A2(n33739), .ZN(N46222));
    NOR2X1 U33351 (.A1(n41772), .A2(n39650), .ZN(N46223));
    INVX1 U33352 (.I(n37397), .ZN(n46224));
    NOR2X1 U33353 (.A1(n42396), .A2(n23484), .ZN(n46225));
    NANDX1 U33354 (.A1(N2771), .A2(N392), .ZN(N46226));
    NOR2X1 U33355 (.A1(n15250), .A2(N1255), .ZN(N46227));
    INVX1 U33356 (.I(N11370), .ZN(N46228));
    NOR2X1 U33357 (.A1(N7871), .A2(n21700), .ZN(N46229));
    NANDX1 U33358 (.A1(n32208), .A2(N12737), .ZN(N46230));
    INVX1 U33359 (.I(n41444), .ZN(N46231));
    INVX1 U33360 (.I(n18997), .ZN(N46232));
    NANDX1 U33361 (.A1(n37293), .A2(N5817), .ZN(N46233));
    NANDX1 U33362 (.A1(n17239), .A2(n35871), .ZN(N46234));
    NANDX1 U33363 (.A1(N3097), .A2(N1367), .ZN(N46235));
    INVX1 U33364 (.I(n35404), .ZN(N46236));
    NOR2X1 U33365 (.A1(n36441), .A2(n13818), .ZN(N46237));
    INVX1 U33366 (.I(n36832), .ZN(N46238));
    INVX1 U33367 (.I(n41143), .ZN(N46239));
    NANDX1 U33368 (.A1(N5097), .A2(N9040), .ZN(n46240));
    INVX1 U33369 (.I(n12967), .ZN(N46241));
    INVX1 U33370 (.I(n20492), .ZN(N46242));
    INVX1 U33371 (.I(n33155), .ZN(N46243));
    INVX1 U33372 (.I(n22505), .ZN(N46244));
    NANDX1 U33373 (.A1(n17292), .A2(n13816), .ZN(N46245));
    NOR2X1 U33374 (.A1(N12789), .A2(N11717), .ZN(N46246));
    NANDX1 U33375 (.A1(N5187), .A2(N7918), .ZN(N46247));
    NANDX1 U33376 (.A1(n39705), .A2(n20875), .ZN(N46248));
    INVX1 U33377 (.I(n29675), .ZN(N46249));
    NANDX1 U33378 (.A1(n40485), .A2(n22416), .ZN(n46250));
    NANDX1 U33379 (.A1(n31748), .A2(N9766), .ZN(N46251));
    INVX1 U33380 (.I(n36844), .ZN(N46252));
    INVX1 U33381 (.I(n25211), .ZN(N46253));
    NANDX1 U33382 (.A1(N6071), .A2(n35382), .ZN(N46254));
    INVX1 U33383 (.I(n28905), .ZN(N46255));
    NOR2X1 U33384 (.A1(n43056), .A2(n36974), .ZN(N46256));
    NOR2X1 U33385 (.A1(n13399), .A2(n28544), .ZN(N46257));
    NOR2X1 U33386 (.A1(n14796), .A2(n27032), .ZN(N46258));
    INVX1 U33387 (.I(N12393), .ZN(n46259));
    NANDX1 U33388 (.A1(n34215), .A2(n33268), .ZN(N46260));
    NANDX1 U33389 (.A1(n20417), .A2(n36790), .ZN(N46261));
    INVX1 U33390 (.I(n32512), .ZN(N46262));
    INVX1 U33391 (.I(n30250), .ZN(N46263));
    NOR2X1 U33392 (.A1(N4528), .A2(n13301), .ZN(N46264));
    INVX1 U33393 (.I(n19418), .ZN(N46265));
    INVX1 U33394 (.I(N3039), .ZN(n46266));
    NOR2X1 U33395 (.A1(n19550), .A2(n31943), .ZN(N46267));
    NOR2X1 U33396 (.A1(n19133), .A2(n15125), .ZN(N46268));
    NANDX1 U33397 (.A1(n22212), .A2(N196), .ZN(N46269));
    NANDX1 U33398 (.A1(n37007), .A2(n16907), .ZN(N46270));
    NOR2X1 U33399 (.A1(N5927), .A2(n24882), .ZN(N46271));
    NOR2X1 U33400 (.A1(n28874), .A2(n36692), .ZN(N46272));
    NANDX1 U33401 (.A1(n22192), .A2(n24874), .ZN(N46273));
    NANDX1 U33402 (.A1(N2071), .A2(N11652), .ZN(N46274));
    NOR2X1 U33403 (.A1(n39750), .A2(n14632), .ZN(N46275));
    INVX1 U33404 (.I(N5375), .ZN(N46276));
    NANDX1 U33405 (.A1(n29405), .A2(N6381), .ZN(N46277));
    NANDX1 U33406 (.A1(N7555), .A2(n20423), .ZN(N46278));
    INVX1 U33407 (.I(n22679), .ZN(n46279));
    NOR2X1 U33408 (.A1(n20731), .A2(N12554), .ZN(N46280));
    INVX1 U33409 (.I(N3945), .ZN(N46281));
    NOR2X1 U33410 (.A1(N8784), .A2(n43023), .ZN(N46282));
    INVX1 U33411 (.I(N7089), .ZN(N46283));
    NANDX1 U33412 (.A1(n26920), .A2(n15490), .ZN(N46284));
    NANDX1 U33413 (.A1(N8322), .A2(N2610), .ZN(N46285));
    INVX1 U33414 (.I(N9653), .ZN(N46286));
    INVX1 U33415 (.I(n18004), .ZN(n46287));
    INVX1 U33416 (.I(n37733), .ZN(N46288));
    INVX1 U33417 (.I(n27594), .ZN(N46289));
    NANDX1 U33418 (.A1(n19439), .A2(N6980), .ZN(N46290));
    NANDX1 U33419 (.A1(n39861), .A2(N5499), .ZN(N46291));
    NOR2X1 U33420 (.A1(n40541), .A2(n15909), .ZN(N46292));
    NANDX1 U33421 (.A1(n31442), .A2(N9533), .ZN(N46293));
    NANDX1 U33422 (.A1(n40226), .A2(N9084), .ZN(n46294));
    NOR2X1 U33423 (.A1(n36994), .A2(n16868), .ZN(N46295));
    INVX1 U33424 (.I(n42163), .ZN(N46296));
    NOR2X1 U33425 (.A1(n13796), .A2(n34452), .ZN(N46297));
    NOR2X1 U33426 (.A1(n23448), .A2(N12667), .ZN(N46298));
    NANDX1 U33427 (.A1(N4259), .A2(N6927), .ZN(N46299));
    INVX1 U33428 (.I(n21532), .ZN(n46300));
    INVX1 U33429 (.I(n42443), .ZN(n46301));
    NANDX1 U33430 (.A1(n41169), .A2(n28511), .ZN(N46302));
    INVX1 U33431 (.I(n41274), .ZN(N46303));
    INVX1 U33432 (.I(n39599), .ZN(N46304));
    NANDX1 U33433 (.A1(n13549), .A2(N5659), .ZN(N46305));
    INVX1 U33434 (.I(n43454), .ZN(N46306));
    INVX1 U33435 (.I(N173), .ZN(N46307));
    NANDX1 U33436 (.A1(n21289), .A2(N5647), .ZN(n46308));
    NOR2X1 U33437 (.A1(n24659), .A2(n19442), .ZN(N46309));
    NANDX1 U33438 (.A1(N6283), .A2(n32569), .ZN(N46310));
    NANDX1 U33439 (.A1(N5909), .A2(n26508), .ZN(N46311));
    INVX1 U33440 (.I(n28913), .ZN(N46312));
    NANDX1 U33441 (.A1(n25227), .A2(n17563), .ZN(n46313));
    NOR2X1 U33442 (.A1(n22923), .A2(N2602), .ZN(N46314));
    NANDX1 U33443 (.A1(N10405), .A2(n17861), .ZN(N46315));
    NOR2X1 U33444 (.A1(N225), .A2(n21089), .ZN(N46316));
    INVX1 U33445 (.I(n21843), .ZN(N46317));
    INVX1 U33446 (.I(n42334), .ZN(N46318));
    NANDX1 U33447 (.A1(N4253), .A2(n20150), .ZN(N46319));
    NOR2X1 U33448 (.A1(n19278), .A2(n34489), .ZN(N46320));
    INVX1 U33449 (.I(n35602), .ZN(N46321));
    INVX1 U33450 (.I(n15560), .ZN(N46322));
    NOR2X1 U33451 (.A1(N3207), .A2(n31747), .ZN(N46323));
    INVX1 U33452 (.I(n32120), .ZN(N46324));
    NANDX1 U33453 (.A1(n40982), .A2(N6210), .ZN(N46325));
    NOR2X1 U33454 (.A1(n20432), .A2(n41963), .ZN(N46326));
    NANDX1 U33455 (.A1(n20516), .A2(n16351), .ZN(N46327));
    INVX1 U33456 (.I(n20740), .ZN(N46328));
    INVX1 U33457 (.I(n22434), .ZN(N46329));
    INVX1 U33458 (.I(n37870), .ZN(N46330));
    NOR2X1 U33459 (.A1(N10805), .A2(n42122), .ZN(N46331));
    INVX1 U33460 (.I(n17826), .ZN(N46332));
    NANDX1 U33461 (.A1(n22141), .A2(N816), .ZN(N46333));
    NOR2X1 U33462 (.A1(n19439), .A2(N6055), .ZN(n46334));
    NOR2X1 U33463 (.A1(n22645), .A2(n37801), .ZN(n46335));
    NOR2X1 U33464 (.A1(N972), .A2(n20322), .ZN(N46336));
    NANDX1 U33465 (.A1(N7182), .A2(n35920), .ZN(N46337));
    NANDX1 U33466 (.A1(n38824), .A2(N11021), .ZN(N46338));
    INVX1 U33467 (.I(N11703), .ZN(N46339));
    INVX1 U33468 (.I(N11054), .ZN(N46340));
    NOR2X1 U33469 (.A1(n40808), .A2(n43315), .ZN(N46341));
    NANDX1 U33470 (.A1(n18631), .A2(N327), .ZN(N46342));
    NANDX1 U33471 (.A1(N6283), .A2(n18152), .ZN(N46343));
    NANDX1 U33472 (.A1(n18103), .A2(N8648), .ZN(N46344));
    INVX1 U33473 (.I(n37541), .ZN(N46345));
    INVX1 U33474 (.I(N8465), .ZN(N46346));
    NOR2X1 U33475 (.A1(n42183), .A2(n14114), .ZN(N46347));
    NOR2X1 U33476 (.A1(n19032), .A2(n17273), .ZN(N46348));
    NANDX1 U33477 (.A1(N11479), .A2(n30543), .ZN(N46349));
    INVX1 U33478 (.I(N12179), .ZN(N46350));
    NANDX1 U33479 (.A1(N959), .A2(n40873), .ZN(N46351));
    NANDX1 U33480 (.A1(n29460), .A2(n38208), .ZN(N46352));
    INVX1 U33481 (.I(N8886), .ZN(N46353));
    NOR2X1 U33482 (.A1(N11438), .A2(n20114), .ZN(N46354));
    NANDX1 U33483 (.A1(n19270), .A2(n38948), .ZN(N46355));
    INVX1 U33484 (.I(n17597), .ZN(N46356));
    INVX1 U33485 (.I(N858), .ZN(N46357));
    INVX1 U33486 (.I(N12189), .ZN(N46358));
    INVX1 U33487 (.I(n20688), .ZN(N46359));
    INVX1 U33488 (.I(n14615), .ZN(N46360));
    NOR2X1 U33489 (.A1(N103), .A2(N8520), .ZN(N46361));
    INVX1 U33490 (.I(n30645), .ZN(N46362));
    NANDX1 U33491 (.A1(N9583), .A2(n41180), .ZN(n46363));
    INVX1 U33492 (.I(n40135), .ZN(n46364));
    INVX1 U33493 (.I(n28194), .ZN(N46365));
    INVX1 U33494 (.I(n20088), .ZN(N46366));
    NOR2X1 U33495 (.A1(n27596), .A2(n21205), .ZN(N46367));
    NANDX1 U33496 (.A1(n26604), .A2(n30154), .ZN(N46368));
    INVX1 U33497 (.I(N241), .ZN(N46369));
    INVX1 U33498 (.I(N2600), .ZN(N46370));
    INVX1 U33499 (.I(n15936), .ZN(N46371));
    INVX1 U33500 (.I(n41501), .ZN(N46372));
    NANDX1 U33501 (.A1(n30771), .A2(N2323), .ZN(N46373));
    NOR2X1 U33502 (.A1(n20553), .A2(N10842), .ZN(N46374));
    NOR2X1 U33503 (.A1(n40877), .A2(N8617), .ZN(N46375));
    INVX1 U33504 (.I(n28264), .ZN(N46376));
    NANDX1 U33505 (.A1(n38711), .A2(n37240), .ZN(N46377));
    NOR2X1 U33506 (.A1(n19789), .A2(n13855), .ZN(N46378));
    NOR2X1 U33507 (.A1(N3913), .A2(n24740), .ZN(N46379));
    NANDX1 U33508 (.A1(n30516), .A2(N11421), .ZN(N46380));
    NANDX1 U33509 (.A1(n20436), .A2(N5379), .ZN(N46381));
    NOR2X1 U33510 (.A1(N11214), .A2(n21314), .ZN(N46382));
    NOR2X1 U33511 (.A1(N9242), .A2(N4144), .ZN(n46383));
    INVX1 U33512 (.I(N11564), .ZN(N46384));
    NOR2X1 U33513 (.A1(n38216), .A2(N12085), .ZN(N46385));
    INVX1 U33514 (.I(n25300), .ZN(n46386));
    INVX1 U33515 (.I(n14263), .ZN(N46387));
    NOR2X1 U33516 (.A1(n28052), .A2(N9501), .ZN(N46388));
    INVX1 U33517 (.I(N9804), .ZN(N46389));
    INVX1 U33518 (.I(N7394), .ZN(n46390));
    NANDX1 U33519 (.A1(n22882), .A2(n32133), .ZN(N46391));
    NOR2X1 U33520 (.A1(N9925), .A2(N81), .ZN(n46392));
    NANDX1 U33521 (.A1(n20040), .A2(N5459), .ZN(N46393));
    NOR2X1 U33522 (.A1(n31254), .A2(n16452), .ZN(N46394));
    NOR2X1 U33523 (.A1(n30175), .A2(n20596), .ZN(N46395));
    NANDX1 U33524 (.A1(n31419), .A2(n36968), .ZN(N46396));
    INVX1 U33525 (.I(N31), .ZN(N46397));
    INVX1 U33526 (.I(N4566), .ZN(N46398));
    NOR2X1 U33527 (.A1(n23444), .A2(n14657), .ZN(N46399));
    NOR2X1 U33528 (.A1(n22625), .A2(N8195), .ZN(N46400));
    NANDX1 U33529 (.A1(N8442), .A2(n15588), .ZN(N46401));
    NANDX1 U33530 (.A1(n31323), .A2(n37400), .ZN(N46402));
    NANDX1 U33531 (.A1(n30927), .A2(n27161), .ZN(N46403));
    NANDX1 U33532 (.A1(n40646), .A2(n22299), .ZN(N46404));
    INVX1 U33533 (.I(n18107), .ZN(N46405));
    INVX1 U33534 (.I(n33042), .ZN(N46406));
    NANDX1 U33535 (.A1(n15874), .A2(n27884), .ZN(N46407));
    INVX1 U33536 (.I(n42521), .ZN(N46408));
    INVX1 U33537 (.I(n25938), .ZN(N46409));
    NANDX1 U33538 (.A1(N11715), .A2(n36350), .ZN(N46410));
    NOR2X1 U33539 (.A1(n16051), .A2(n21021), .ZN(N46411));
    INVX1 U33540 (.I(n24245), .ZN(N46412));
    NOR2X1 U33541 (.A1(n42099), .A2(n29513), .ZN(N46413));
    NANDX1 U33542 (.A1(n19629), .A2(n23440), .ZN(N46414));
    INVX1 U33543 (.I(n40235), .ZN(N46415));
    NANDX1 U33544 (.A1(N8653), .A2(n27089), .ZN(N46416));
    NANDX1 U33545 (.A1(n21044), .A2(N1723), .ZN(N46417));
    NANDX1 U33546 (.A1(N10613), .A2(n39684), .ZN(n46418));
    INVX1 U33547 (.I(n28177), .ZN(N46419));
    INVX1 U33548 (.I(N8666), .ZN(N46420));
    NANDX1 U33549 (.A1(N4585), .A2(N6576), .ZN(N46421));
    NANDX1 U33550 (.A1(n30614), .A2(n27930), .ZN(N46422));
    NOR2X1 U33551 (.A1(n41314), .A2(n18115), .ZN(N46423));
    NOR2X1 U33552 (.A1(N3016), .A2(N6422), .ZN(N46424));
    NANDX1 U33553 (.A1(N340), .A2(n15730), .ZN(N46425));
    INVX1 U33554 (.I(N9718), .ZN(N46426));
    NOR2X1 U33555 (.A1(N8869), .A2(N8050), .ZN(n46427));
    NANDX1 U33556 (.A1(n27975), .A2(n29093), .ZN(N46428));
    NOR2X1 U33557 (.A1(n32039), .A2(n29385), .ZN(N46429));
    NANDX1 U33558 (.A1(n41656), .A2(n14089), .ZN(N46430));
    NANDX1 U33559 (.A1(N6850), .A2(n28774), .ZN(N46431));
    NOR2X1 U33560 (.A1(n13425), .A2(N11701), .ZN(N46432));
    INVX1 U33561 (.I(n31034), .ZN(N46433));
    NANDX1 U33562 (.A1(n18239), .A2(N5677), .ZN(N46434));
    NOR2X1 U33563 (.A1(n21255), .A2(N1778), .ZN(N46435));
    INVX1 U33564 (.I(N11274), .ZN(N46436));
    INVX1 U33565 (.I(n34582), .ZN(N46437));
    NOR2X1 U33566 (.A1(n29999), .A2(n43451), .ZN(N46438));
    INVX1 U33567 (.I(n15787), .ZN(N46439));
    NOR2X1 U33568 (.A1(N4340), .A2(N3298), .ZN(N46440));
    NANDX1 U33569 (.A1(n23404), .A2(n30492), .ZN(N46441));
    NANDX1 U33570 (.A1(n37493), .A2(n26012), .ZN(N46442));
    NANDX1 U33571 (.A1(N12474), .A2(n26117), .ZN(N46443));
    NANDX1 U33572 (.A1(n24175), .A2(N3042), .ZN(N46444));
    NANDX1 U33573 (.A1(n34852), .A2(n21281), .ZN(N46445));
    NOR2X1 U33574 (.A1(N4639), .A2(n32215), .ZN(N46446));
    INVX1 U33575 (.I(n27160), .ZN(N46447));
    NOR2X1 U33576 (.A1(n39370), .A2(N7949), .ZN(N46448));
    NANDX1 U33577 (.A1(n15576), .A2(N7927), .ZN(N46449));
    NOR2X1 U33578 (.A1(n31363), .A2(n15240), .ZN(N46450));
    INVX1 U33579 (.I(n24340), .ZN(N46451));
    NOR2X1 U33580 (.A1(n26187), .A2(N11359), .ZN(N46452));
    INVX1 U33581 (.I(n20207), .ZN(N46453));
    INVX1 U33582 (.I(n39245), .ZN(N46454));
    NOR2X1 U33583 (.A1(N9694), .A2(n43261), .ZN(N46455));
    NOR2X1 U33584 (.A1(N12736), .A2(n34838), .ZN(N46456));
    NANDX1 U33585 (.A1(n23696), .A2(N11452), .ZN(N46457));
    INVX1 U33586 (.I(N12438), .ZN(n46458));
    NANDX1 U33587 (.A1(n15920), .A2(n35285), .ZN(N46459));
    INVX1 U33588 (.I(n23868), .ZN(N46460));
    NOR2X1 U33589 (.A1(N1315), .A2(n21475), .ZN(N46461));
    NANDX1 U33590 (.A1(n22357), .A2(n36714), .ZN(N46462));
    NOR2X1 U33591 (.A1(N3224), .A2(N4360), .ZN(N46463));
    NANDX1 U33592 (.A1(N4262), .A2(n42692), .ZN(N46464));
    INVX1 U33593 (.I(n31311), .ZN(N46465));
    INVX1 U33594 (.I(n18686), .ZN(N46466));
    NANDX1 U33595 (.A1(n38252), .A2(N11428), .ZN(N46467));
    INVX1 U33596 (.I(n19298), .ZN(N46468));
    INVX1 U33597 (.I(n23643), .ZN(N46469));
    NOR2X1 U33598 (.A1(n27781), .A2(n25760), .ZN(N46470));
    INVX1 U33599 (.I(N228), .ZN(N46471));
    INVX1 U33600 (.I(n39481), .ZN(N46472));
    INVX1 U33601 (.I(N9749), .ZN(N46473));
    NOR2X1 U33602 (.A1(n35250), .A2(N370), .ZN(N46474));
    NOR2X1 U33603 (.A1(n18171), .A2(n37246), .ZN(N46475));
    NOR2X1 U33604 (.A1(N12210), .A2(n13364), .ZN(N46476));
    NANDX1 U33605 (.A1(N11429), .A2(n42841), .ZN(N46477));
    NOR2X1 U33606 (.A1(N6421), .A2(N7734), .ZN(N46478));
    INVX1 U33607 (.I(N1200), .ZN(N46479));
    INVX1 U33608 (.I(n35312), .ZN(N46480));
    INVX1 U33609 (.I(n14710), .ZN(N46481));
    INVX1 U33610 (.I(n40925), .ZN(n46482));
    NANDX1 U33611 (.A1(n41241), .A2(N7723), .ZN(N46483));
    NOR2X1 U33612 (.A1(n15340), .A2(n36883), .ZN(N46484));
    NOR2X1 U33613 (.A1(n14768), .A2(n23885), .ZN(N46485));
    INVX1 U33614 (.I(N4817), .ZN(N46486));
    INVX1 U33615 (.I(n35480), .ZN(N46487));
    NOR2X1 U33616 (.A1(N2352), .A2(N4217), .ZN(n46488));
    NANDX1 U33617 (.A1(N8874), .A2(n15645), .ZN(N46489));
    NOR2X1 U33618 (.A1(n36386), .A2(N11745), .ZN(N46490));
    NANDX1 U33619 (.A1(n28279), .A2(N2625), .ZN(N46491));
    NANDX1 U33620 (.A1(n20118), .A2(N12801), .ZN(N46492));
    INVX1 U33621 (.I(n25280), .ZN(N46493));
    NANDX1 U33622 (.A1(n31303), .A2(N12728), .ZN(N46494));
    NOR2X1 U33623 (.A1(N9908), .A2(n17748), .ZN(N46495));
    INVX1 U33624 (.I(N2288), .ZN(N46496));
    NANDX1 U33625 (.A1(n14630), .A2(n19597), .ZN(N46497));
    NANDX1 U33626 (.A1(N4400), .A2(N11604), .ZN(N46498));
    NANDX1 U33627 (.A1(n39903), .A2(N5500), .ZN(N46499));
    NOR2X1 U33628 (.A1(n38456), .A2(n21144), .ZN(N46500));
    NOR2X1 U33629 (.A1(n31369), .A2(n22569), .ZN(N46501));
    INVX1 U33630 (.I(n16175), .ZN(n46502));
    NANDX1 U33631 (.A1(N11074), .A2(n25973), .ZN(N46503));
    NANDX1 U33632 (.A1(n43359), .A2(n40932), .ZN(n46504));
    NOR2X1 U33633 (.A1(n20869), .A2(N10187), .ZN(N46505));
    NOR2X1 U33634 (.A1(n30776), .A2(n27934), .ZN(N46506));
    INVX1 U33635 (.I(n22743), .ZN(N46507));
    NANDX1 U33636 (.A1(n40635), .A2(n42339), .ZN(N46508));
    NOR2X1 U33637 (.A1(N1562), .A2(N10470), .ZN(N46509));
    INVX1 U33638 (.I(n31144), .ZN(N46510));
    NANDX1 U33639 (.A1(n22390), .A2(n26127), .ZN(N46511));
    INVX1 U33640 (.I(n29985), .ZN(N46512));
    NOR2X1 U33641 (.A1(n39040), .A2(n13163), .ZN(N46513));
    NANDX1 U33642 (.A1(n20760), .A2(n13916), .ZN(N46514));
    INVX1 U33643 (.I(N4961), .ZN(N46515));
    NOR2X1 U33644 (.A1(n43309), .A2(n42886), .ZN(n46516));
    NOR2X1 U33645 (.A1(n43176), .A2(n24355), .ZN(N46517));
    NANDX1 U33646 (.A1(n27637), .A2(N6888), .ZN(N46518));
    NOR2X1 U33647 (.A1(n23973), .A2(n37203), .ZN(N46519));
    INVX1 U33648 (.I(N3848), .ZN(N46520));
    NANDX1 U33649 (.A1(N12770), .A2(N9324), .ZN(N46521));
    NANDX1 U33650 (.A1(n18418), .A2(n21393), .ZN(n46522));
    INVX1 U33651 (.I(n34890), .ZN(N46523));
    NANDX1 U33652 (.A1(N2473), .A2(n20137), .ZN(N46524));
    NOR2X1 U33653 (.A1(n22351), .A2(n40897), .ZN(N46525));
    NANDX1 U33654 (.A1(n14408), .A2(n35537), .ZN(N46526));
    NANDX1 U33655 (.A1(N3925), .A2(n34950), .ZN(N46527));
    NANDX1 U33656 (.A1(N3628), .A2(N5512), .ZN(N46528));
    INVX1 U33657 (.I(n20944), .ZN(N46529));
    INVX1 U33658 (.I(n36620), .ZN(N46530));
    INVX1 U33659 (.I(n39282), .ZN(N46531));
    INVX1 U33660 (.I(N5292), .ZN(N46532));
    NOR2X1 U33661 (.A1(N8218), .A2(N4295), .ZN(N46533));
    INVX1 U33662 (.I(n16316), .ZN(N46534));
    NOR2X1 U33663 (.A1(n39138), .A2(n40885), .ZN(n46535));
    NANDX1 U33664 (.A1(n41610), .A2(n17549), .ZN(N46536));
    INVX1 U33665 (.I(N10168), .ZN(N46537));
    INVX1 U33666 (.I(N4887), .ZN(N46538));
    INVX1 U33667 (.I(n40189), .ZN(N46539));
    NANDX1 U33668 (.A1(n28500), .A2(n21347), .ZN(N46540));
    NOR2X1 U33669 (.A1(n21807), .A2(n26858), .ZN(N46541));
    NOR2X1 U33670 (.A1(n42750), .A2(n28937), .ZN(N46542));
    INVX1 U33671 (.I(n33874), .ZN(N46543));
    INVX1 U33672 (.I(N12231), .ZN(N46544));
    NANDX1 U33673 (.A1(N5527), .A2(n20448), .ZN(N46545));
    NOR2X1 U33674 (.A1(N2422), .A2(n36763), .ZN(N46546));
    NOR2X1 U33675 (.A1(n31239), .A2(n23855), .ZN(N46547));
    INVX1 U33676 (.I(n29377), .ZN(N46548));
    INVX1 U33677 (.I(n41682), .ZN(N46549));
    NANDX1 U33678 (.A1(n35736), .A2(n36248), .ZN(N46550));
    NOR2X1 U33679 (.A1(n32453), .A2(N5165), .ZN(N46551));
    NOR2X1 U33680 (.A1(N7), .A2(N5934), .ZN(N46552));
    NOR2X1 U33681 (.A1(n16544), .A2(n29569), .ZN(N46553));
    NANDX1 U33682 (.A1(N2009), .A2(N2879), .ZN(N46554));
    NOR2X1 U33683 (.A1(n16434), .A2(n15109), .ZN(N46555));
    NANDX1 U33684 (.A1(N11640), .A2(n25236), .ZN(N46556));
    NANDX1 U33685 (.A1(n14062), .A2(N8207), .ZN(N46557));
    NANDX1 U33686 (.A1(n34980), .A2(n32061), .ZN(N46558));
    NANDX1 U33687 (.A1(n20884), .A2(n29992), .ZN(N46559));
    INVX1 U33688 (.I(N6636), .ZN(N46560));
    INVX1 U33689 (.I(n41546), .ZN(N46561));
    INVX1 U33690 (.I(N916), .ZN(N46562));
    INVX1 U33691 (.I(N12316), .ZN(N46563));
    INVX1 U33692 (.I(n42324), .ZN(N46564));
    INVX1 U33693 (.I(N7145), .ZN(N46565));
    INVX1 U33694 (.I(n14952), .ZN(N46566));
    NANDX1 U33695 (.A1(n20978), .A2(N1151), .ZN(N46567));
    INVX1 U33696 (.I(n25766), .ZN(N46568));
    NANDX1 U33697 (.A1(n26906), .A2(N7529), .ZN(N46569));
    INVX1 U33698 (.I(n30647), .ZN(N46570));
    INVX1 U33699 (.I(n40970), .ZN(N46571));
    NOR2X1 U33700 (.A1(N4324), .A2(n14908), .ZN(N46572));
    NANDX1 U33701 (.A1(n23995), .A2(n30526), .ZN(N46573));
    NOR2X1 U33702 (.A1(n35930), .A2(n18280), .ZN(N46574));
    INVX1 U33703 (.I(n26525), .ZN(N46575));
    NOR2X1 U33704 (.A1(n14838), .A2(n17126), .ZN(N46576));
    NANDX1 U33705 (.A1(n23672), .A2(n24271), .ZN(N46577));
    NANDX1 U33706 (.A1(n28304), .A2(n23103), .ZN(N46578));
    INVX1 U33707 (.I(n29454), .ZN(N46579));
    NANDX1 U33708 (.A1(N10777), .A2(N12495), .ZN(N46580));
    NOR2X1 U33709 (.A1(n18306), .A2(N248), .ZN(N46581));
    NOR2X1 U33710 (.A1(n23720), .A2(n30897), .ZN(N46582));
    NOR2X1 U33711 (.A1(n28043), .A2(N2332), .ZN(N46583));
    NANDX1 U33712 (.A1(N8566), .A2(n22538), .ZN(N46584));
    NANDX1 U33713 (.A1(n34175), .A2(n40817), .ZN(N46585));
    NOR2X1 U33714 (.A1(n17228), .A2(n41693), .ZN(N46586));
    INVX1 U33715 (.I(n34353), .ZN(N46587));
    NANDX1 U33716 (.A1(N5688), .A2(n15151), .ZN(N46588));
    INVX1 U33717 (.I(n33991), .ZN(N46589));
    NOR2X1 U33718 (.A1(n23619), .A2(N9652), .ZN(N46590));
    NANDX1 U33719 (.A1(n24075), .A2(N11826), .ZN(N46591));
    INVX1 U33720 (.I(n42380), .ZN(N46592));
    INVX1 U33721 (.I(N12329), .ZN(N46593));
    NOR2X1 U33722 (.A1(n42970), .A2(N12499), .ZN(N46594));
    INVX1 U33723 (.I(n34981), .ZN(n46595));
    NOR2X1 U33724 (.A1(n38595), .A2(n14046), .ZN(N46596));
    NANDX1 U33725 (.A1(n29298), .A2(N1070), .ZN(N46597));
    INVX1 U33726 (.I(N3053), .ZN(N46598));
    NOR2X1 U33727 (.A1(n13030), .A2(n27085), .ZN(N46599));
    NANDX1 U33728 (.A1(n18717), .A2(n42236), .ZN(n46600));
    NANDX1 U33729 (.A1(n42387), .A2(n26697), .ZN(N46601));
    NOR2X1 U33730 (.A1(n41718), .A2(N6054), .ZN(N46602));
    INVX1 U33731 (.I(N10071), .ZN(N46603));
    NOR2X1 U33732 (.A1(N8013), .A2(N11824), .ZN(N46604));
    INVX1 U33733 (.I(n20320), .ZN(N46605));
    NOR2X1 U33734 (.A1(N1080), .A2(n17198), .ZN(N46606));
    NANDX1 U33735 (.A1(n36147), .A2(N12320), .ZN(n46607));
    INVX1 U33736 (.I(N2718), .ZN(N46608));
    INVX1 U33737 (.I(N7624), .ZN(N46609));
    INVX1 U33738 (.I(n24029), .ZN(N46610));
    INVX1 U33739 (.I(n36440), .ZN(N46611));
    NOR2X1 U33740 (.A1(n16664), .A2(N1364), .ZN(N46612));
    NOR2X1 U33741 (.A1(n31869), .A2(n33430), .ZN(N46613));
    NANDX1 U33742 (.A1(n16899), .A2(n31675), .ZN(N46614));
    NOR2X1 U33743 (.A1(n26004), .A2(n31426), .ZN(N46615));
    NANDX1 U33744 (.A1(n34017), .A2(n43249), .ZN(N46616));
    NOR2X1 U33745 (.A1(N544), .A2(N777), .ZN(N46617));
    NOR2X1 U33746 (.A1(n17741), .A2(n36757), .ZN(N46618));
    INVX1 U33747 (.I(n19741), .ZN(N46619));
    NANDX1 U33748 (.A1(n12971), .A2(n40717), .ZN(N46620));
    INVX1 U33749 (.I(n26061), .ZN(N46621));
    NANDX1 U33750 (.A1(n26888), .A2(N8709), .ZN(N46622));
    INVX1 U33751 (.I(N80), .ZN(N46623));
    NOR2X1 U33752 (.A1(n24999), .A2(n21628), .ZN(N46624));
    NANDX1 U33753 (.A1(n37459), .A2(n28206), .ZN(N46625));
    NANDX1 U33754 (.A1(N12500), .A2(N10738), .ZN(N46626));
    NOR2X1 U33755 (.A1(N7267), .A2(n34434), .ZN(N46627));
    INVX1 U33756 (.I(n34086), .ZN(N46628));
    NANDX1 U33757 (.A1(n32721), .A2(n18513), .ZN(N46629));
    NANDX1 U33758 (.A1(n15686), .A2(n28766), .ZN(n46630));
    INVX1 U33759 (.I(n38356), .ZN(N46631));
    NANDX1 U33760 (.A1(n38742), .A2(n25178), .ZN(N46632));
    INVX1 U33761 (.I(n16543), .ZN(N46633));
    NANDX1 U33762 (.A1(n22713), .A2(n35137), .ZN(N46634));
    NANDX1 U33763 (.A1(n22464), .A2(N6343), .ZN(N46635));
    NOR2X1 U33764 (.A1(N12173), .A2(N329), .ZN(N46636));
    NANDX1 U33765 (.A1(n12917), .A2(N12829), .ZN(N46637));
    NOR2X1 U33766 (.A1(N1613), .A2(n20095), .ZN(N46638));
    INVX1 U33767 (.I(n33558), .ZN(N46639));
    NOR2X1 U33768 (.A1(N108), .A2(N12486), .ZN(N46640));
    INVX1 U33769 (.I(n32185), .ZN(N46641));
    INVX1 U33770 (.I(N4194), .ZN(N46642));
    NANDX1 U33771 (.A1(N12735), .A2(n35610), .ZN(N46643));
    INVX1 U33772 (.I(n27592), .ZN(N46644));
    INVX1 U33773 (.I(n31702), .ZN(N46645));
    INVX1 U33774 (.I(N8214), .ZN(N46646));
    INVX1 U33775 (.I(n24217), .ZN(N46647));
    NOR2X1 U33776 (.A1(n29709), .A2(n23556), .ZN(N46648));
    NANDX1 U33777 (.A1(n19717), .A2(N7629), .ZN(N46649));
    NANDX1 U33778 (.A1(n32545), .A2(n35590), .ZN(N46650));
    NANDX1 U33779 (.A1(n42319), .A2(N721), .ZN(N46651));
    INVX1 U33780 (.I(n42707), .ZN(n46652));
    NOR2X1 U33781 (.A1(n39309), .A2(n18135), .ZN(N46653));
    INVX1 U33782 (.I(n13687), .ZN(N46654));
    NANDX1 U33783 (.A1(n32261), .A2(n16101), .ZN(N46655));
    NANDX1 U33784 (.A1(N3947), .A2(N221), .ZN(N46656));
    NANDX1 U33785 (.A1(n35648), .A2(n26085), .ZN(N46657));
    NANDX1 U33786 (.A1(N5222), .A2(N6830), .ZN(N46658));
    NOR2X1 U33787 (.A1(n24610), .A2(n20065), .ZN(N46659));
    NANDX1 U33788 (.A1(N854), .A2(n17373), .ZN(N46660));
    NOR2X1 U33789 (.A1(n23079), .A2(N9491), .ZN(N46661));
    NANDX1 U33790 (.A1(n21925), .A2(n43363), .ZN(N46662));
    INVX1 U33791 (.I(N10839), .ZN(n46663));
    NANDX1 U33792 (.A1(N4530), .A2(n28973), .ZN(N46664));
    NANDX1 U33793 (.A1(N7896), .A2(n30661), .ZN(N46665));
    NANDX1 U33794 (.A1(n23997), .A2(n24485), .ZN(N46666));
    INVX1 U33795 (.I(n24217), .ZN(N46667));
    NANDX1 U33796 (.A1(N10511), .A2(n39981), .ZN(N46668));
    INVX1 U33797 (.I(N5412), .ZN(N46669));
    NOR2X1 U33798 (.A1(N9564), .A2(n30021), .ZN(n46670));
    NOR2X1 U33799 (.A1(N6516), .A2(n20554), .ZN(N46671));
    INVX1 U33800 (.I(n38593), .ZN(N46672));
    NOR2X1 U33801 (.A1(n29625), .A2(n20464), .ZN(N46673));
    NANDX1 U33802 (.A1(n29515), .A2(n29157), .ZN(N46674));
    NOR2X1 U33803 (.A1(N9592), .A2(n33686), .ZN(N46675));
    NOR2X1 U33804 (.A1(N2040), .A2(n31261), .ZN(N46676));
    INVX1 U33805 (.I(n26748), .ZN(N46677));
    NANDX1 U33806 (.A1(n42608), .A2(N11931), .ZN(N46678));
    NANDX1 U33807 (.A1(N2946), .A2(N12121), .ZN(N46679));
    NANDX1 U33808 (.A1(n37767), .A2(n17532), .ZN(N46680));
    INVX1 U33809 (.I(N3858), .ZN(N46681));
    NOR2X1 U33810 (.A1(n17969), .A2(N10374), .ZN(N46682));
    INVX1 U33811 (.I(N4952), .ZN(N46683));
    NOR2X1 U33812 (.A1(N4153), .A2(n24256), .ZN(N46684));
    INVX1 U33813 (.I(n15917), .ZN(N46685));
    NOR2X1 U33814 (.A1(N1321), .A2(n28199), .ZN(N46686));
    INVX1 U33815 (.I(n24686), .ZN(N46687));
    NOR2X1 U33816 (.A1(N11610), .A2(N12475), .ZN(N46688));
    NOR2X1 U33817 (.A1(n38357), .A2(n13939), .ZN(N46689));
    NANDX1 U33818 (.A1(n39967), .A2(n39620), .ZN(N46690));
    INVX1 U33819 (.I(N8615), .ZN(N46691));
    INVX1 U33820 (.I(n30160), .ZN(N46692));
    INVX1 U33821 (.I(n12903), .ZN(N46693));
    INVX1 U33822 (.I(N9585), .ZN(N46694));
    NOR2X1 U33823 (.A1(n34071), .A2(n23898), .ZN(N46695));
    NANDX1 U33824 (.A1(n29244), .A2(n28050), .ZN(N46696));
    INVX1 U33825 (.I(N1409), .ZN(N46697));
    NANDX1 U33826 (.A1(N6264), .A2(n35881), .ZN(n46698));
    INVX1 U33827 (.I(n15834), .ZN(N46699));
    INVX1 U33828 (.I(n34034), .ZN(N46700));
    NANDX1 U33829 (.A1(n19249), .A2(n24346), .ZN(N46701));
    NANDX1 U33830 (.A1(n33187), .A2(N3474), .ZN(N46702));
    INVX1 U33831 (.I(n19014), .ZN(N46703));
    INVX1 U33832 (.I(n17116), .ZN(N46704));
    INVX1 U33833 (.I(n26027), .ZN(N46705));
    INVX1 U33834 (.I(n29613), .ZN(n46706));
    NOR2X1 U33835 (.A1(n32206), .A2(n17012), .ZN(N46707));
    NANDX1 U33836 (.A1(N2311), .A2(n32194), .ZN(N46708));
    NOR2X1 U33837 (.A1(n20040), .A2(n28159), .ZN(N46709));
    NANDX1 U33838 (.A1(N10213), .A2(n34423), .ZN(N46710));
    NANDX1 U33839 (.A1(n18265), .A2(N6784), .ZN(n46711));
    NOR2X1 U33840 (.A1(n41978), .A2(n23906), .ZN(N46712));
    NANDX1 U33841 (.A1(N12531), .A2(N2760), .ZN(N46713));
    INVX1 U33842 (.I(n16005), .ZN(N46714));
    NOR2X1 U33843 (.A1(n13380), .A2(N1552), .ZN(N46715));
    NANDX1 U33844 (.A1(n30090), .A2(n17258), .ZN(N46716));
    NOR2X1 U33845 (.A1(N5910), .A2(n23510), .ZN(N46717));
    NANDX1 U33846 (.A1(N12601), .A2(N10039), .ZN(N46718));
    INVX1 U33847 (.I(N1322), .ZN(N46719));
    NOR2X1 U33848 (.A1(n31121), .A2(n29480), .ZN(N46720));
    NANDX1 U33849 (.A1(n31014), .A2(N10110), .ZN(N46721));
    NANDX1 U33850 (.A1(n38958), .A2(N6573), .ZN(N46722));
    NANDX1 U33851 (.A1(n27143), .A2(n30478), .ZN(N46723));
    INVX1 U33852 (.I(n39673), .ZN(n46724));
    NOR2X1 U33853 (.A1(N6044), .A2(N1885), .ZN(N46725));
    NANDX1 U33854 (.A1(N9103), .A2(N3436), .ZN(N46726));
    INVX1 U33855 (.I(n39192), .ZN(N46727));
    INVX1 U33856 (.I(n18479), .ZN(N46728));
    NANDX1 U33857 (.A1(n33883), .A2(n27250), .ZN(N46729));
    INVX1 U33858 (.I(n33601), .ZN(N46730));
    NOR2X1 U33859 (.A1(n38382), .A2(n38773), .ZN(N46731));
    NANDX1 U33860 (.A1(n14070), .A2(N7333), .ZN(N46732));
    INVX1 U33861 (.I(n24179), .ZN(N46733));
    NOR2X1 U33862 (.A1(n42157), .A2(n30752), .ZN(N46734));
    NANDX1 U33863 (.A1(n25827), .A2(n17757), .ZN(N46735));
    NOR2X1 U33864 (.A1(N11708), .A2(n40674), .ZN(N46736));
    NOR2X1 U33865 (.A1(N3272), .A2(n21060), .ZN(N46737));
    NOR2X1 U33866 (.A1(N6708), .A2(n42333), .ZN(N46738));
    NANDX1 U33867 (.A1(n17081), .A2(n17340), .ZN(n46739));
    NOR2X1 U33868 (.A1(n40643), .A2(N1117), .ZN(N46740));
    NANDX1 U33869 (.A1(n20451), .A2(n39447), .ZN(N46741));
    NANDX1 U33870 (.A1(n15751), .A2(N11633), .ZN(N46742));
    INVX1 U33871 (.I(N12764), .ZN(N46743));
    NOR2X1 U33872 (.A1(n14657), .A2(N10758), .ZN(N46744));
    INVX1 U33873 (.I(N1936), .ZN(N46745));
    INVX1 U33874 (.I(n18704), .ZN(N46746));
    NOR2X1 U33875 (.A1(n22155), .A2(n20091), .ZN(N46747));
    NANDX1 U33876 (.A1(n24255), .A2(n23362), .ZN(N46748));
    NANDX1 U33877 (.A1(N2306), .A2(n19749), .ZN(N46749));
    NANDX1 U33878 (.A1(n42380), .A2(n26509), .ZN(N46750));
    NANDX1 U33879 (.A1(n30290), .A2(n13359), .ZN(N46751));
    INVX1 U33880 (.I(n22109), .ZN(N46752));
    INVX1 U33881 (.I(N9962), .ZN(N46753));
    NOR2X1 U33882 (.A1(n39240), .A2(N11275), .ZN(N46754));
    INVX1 U33883 (.I(N8531), .ZN(n46755));
    INVX1 U33884 (.I(N3651), .ZN(N46756));
    NOR2X1 U33885 (.A1(N8663), .A2(N5586), .ZN(N46757));
    INVX1 U33886 (.I(n17046), .ZN(N46758));
    NANDX1 U33887 (.A1(n36581), .A2(n37136), .ZN(N46759));
    NOR2X1 U33888 (.A1(n17363), .A2(N6706), .ZN(N46760));
    INVX1 U33889 (.I(N9348), .ZN(N46761));
    INVX1 U33890 (.I(n13735), .ZN(N46762));
    NANDX1 U33891 (.A1(n42643), .A2(n36927), .ZN(N46763));
    INVX1 U33892 (.I(N12529), .ZN(N46764));
    NOR2X1 U33893 (.A1(N6861), .A2(n36018), .ZN(N46765));
    NOR2X1 U33894 (.A1(N5378), .A2(n31786), .ZN(N46766));
    INVX1 U33895 (.I(n37845), .ZN(N46767));
    NANDX1 U33896 (.A1(n34144), .A2(n31175), .ZN(N46768));
    NANDX1 U33897 (.A1(n42806), .A2(n36761), .ZN(N46769));
    NOR2X1 U33898 (.A1(n16380), .A2(n41398), .ZN(n46770));
    INVX1 U33899 (.I(n43195), .ZN(n46771));
    INVX1 U33900 (.I(n20388), .ZN(N46772));
    NOR2X1 U33901 (.A1(N6698), .A2(n29736), .ZN(N46773));
    NANDX1 U33902 (.A1(n20432), .A2(n27670), .ZN(N46774));
    NANDX1 U33903 (.A1(N3566), .A2(N12422), .ZN(N46775));
    INVX1 U33904 (.I(N11008), .ZN(N46776));
    INVX1 U33905 (.I(n16486), .ZN(N46777));
    NOR2X1 U33906 (.A1(n14340), .A2(N4799), .ZN(N46778));
    INVX1 U33907 (.I(n41864), .ZN(N46779));
    NANDX1 U33908 (.A1(n27119), .A2(n29567), .ZN(N46780));
    INVX1 U33909 (.I(n16132), .ZN(N46781));
    INVX1 U33910 (.I(n40203), .ZN(N46782));
    NOR2X1 U33911 (.A1(N140), .A2(n43228), .ZN(N46783));
    INVX1 U33912 (.I(n32107), .ZN(N46784));
    NOR2X1 U33913 (.A1(n18021), .A2(n38804), .ZN(N46785));
    NANDX1 U33914 (.A1(n40582), .A2(N5443), .ZN(N46786));
    NANDX1 U33915 (.A1(N8521), .A2(n42161), .ZN(N46787));
    INVX1 U33916 (.I(n22141), .ZN(N46788));
    NANDX1 U33917 (.A1(n34819), .A2(n38626), .ZN(n46789));
    NANDX1 U33918 (.A1(n38839), .A2(n33104), .ZN(N46790));
    NANDX1 U33919 (.A1(n26910), .A2(n14105), .ZN(N46791));
    INVX1 U33920 (.I(N2684), .ZN(N46792));
    INVX1 U33921 (.I(n43370), .ZN(N46793));
    NANDX1 U33922 (.A1(n20480), .A2(n22089), .ZN(N46794));
    INVX1 U33923 (.I(N9915), .ZN(N46795));
    INVX1 U33924 (.I(n37143), .ZN(N46796));
    NANDX1 U33925 (.A1(N8230), .A2(n22154), .ZN(N46797));
    INVX1 U33926 (.I(n38492), .ZN(N46798));
    NOR2X1 U33927 (.A1(n18938), .A2(n36692), .ZN(N46799));
    NOR2X1 U33928 (.A1(n34475), .A2(n15360), .ZN(N46800));
    INVX1 U33929 (.I(n25821), .ZN(N46801));
    NANDX1 U33930 (.A1(n32805), .A2(N10867), .ZN(N46802));
    INVX1 U33931 (.I(n32925), .ZN(N46803));
    NOR2X1 U33932 (.A1(n37081), .A2(n16691), .ZN(N46804));
    INVX1 U33933 (.I(n17358), .ZN(N46805));
    INVX1 U33934 (.I(N12206), .ZN(N46806));
    NOR2X1 U33935 (.A1(n18036), .A2(N6922), .ZN(N46807));
    INVX1 U33936 (.I(N8245), .ZN(N46808));
    INVX1 U33937 (.I(N3377), .ZN(N46809));
    NOR2X1 U33938 (.A1(n22746), .A2(N8880), .ZN(N46810));
    NOR2X1 U33939 (.A1(n40022), .A2(n17497), .ZN(n46811));
    NOR2X1 U33940 (.A1(N12514), .A2(N8499), .ZN(N46812));
    NOR2X1 U33941 (.A1(n27853), .A2(n34320), .ZN(N46813));
    INVX1 U33942 (.I(n17185), .ZN(N46814));
    NANDX1 U33943 (.A1(n22601), .A2(N6637), .ZN(N46815));
    INVX1 U33944 (.I(n16209), .ZN(N46816));
    NOR2X1 U33945 (.A1(n26158), .A2(n33566), .ZN(N46817));
    NANDX1 U33946 (.A1(n28043), .A2(n17611), .ZN(N46818));
    NOR2X1 U33947 (.A1(n34964), .A2(N1251), .ZN(N46819));
    INVX1 U33948 (.I(n35556), .ZN(N46820));
    NANDX1 U33949 (.A1(n20749), .A2(N4510), .ZN(N46821));
    NOR2X1 U33950 (.A1(n21922), .A2(n34211), .ZN(N46822));
    NOR2X1 U33951 (.A1(N5994), .A2(N3253), .ZN(N46823));
    NANDX1 U33952 (.A1(N5426), .A2(n20785), .ZN(N46824));
    INVX1 U33953 (.I(n38203), .ZN(N46825));
    INVX1 U33954 (.I(N1102), .ZN(N46826));
    NOR2X1 U33955 (.A1(n23966), .A2(n30271), .ZN(N46827));
    INVX1 U33956 (.I(n36973), .ZN(N46828));
    NANDX1 U33957 (.A1(n13312), .A2(n35607), .ZN(N46829));
    NOR2X1 U33958 (.A1(n20603), .A2(N8804), .ZN(N46830));
    NOR2X1 U33959 (.A1(n21853), .A2(n23398), .ZN(n46831));
    NANDX1 U33960 (.A1(n16159), .A2(N674), .ZN(N46832));
    NOR2X1 U33961 (.A1(n19345), .A2(N12275), .ZN(N46833));
    NANDX1 U33962 (.A1(n29707), .A2(n18269), .ZN(N46834));
    INVX1 U33963 (.I(n15415), .ZN(N46835));
    NOR2X1 U33964 (.A1(n35729), .A2(n14803), .ZN(N46836));
    NOR2X1 U33965 (.A1(n19906), .A2(n15904), .ZN(N46837));
    NANDX1 U33966 (.A1(N400), .A2(n35854), .ZN(N46838));
    NOR2X1 U33967 (.A1(n27052), .A2(n38490), .ZN(N46839));
    NOR2X1 U33968 (.A1(n19186), .A2(n15375), .ZN(N46840));
    INVX1 U33969 (.I(n27989), .ZN(N46841));
    INVX1 U33970 (.I(N7154), .ZN(n46842));
    INVX1 U33971 (.I(N10517), .ZN(N46843));
    NANDX1 U33972 (.A1(n41740), .A2(n41790), .ZN(N46844));
    NANDX1 U33973 (.A1(N10543), .A2(n20330), .ZN(N46845));
    INVX1 U33974 (.I(n18491), .ZN(N46846));
    INVX1 U33975 (.I(n13345), .ZN(N46847));
    NOR2X1 U33976 (.A1(n17211), .A2(n28147), .ZN(N46848));
    INVX1 U33977 (.I(n26796), .ZN(n46849));
    INVX1 U33978 (.I(N1289), .ZN(N46850));
    NANDX1 U33979 (.A1(n15791), .A2(N6469), .ZN(N46851));
    NOR2X1 U33980 (.A1(N488), .A2(n14640), .ZN(N46852));
    NOR2X1 U33981 (.A1(n15863), .A2(N10261), .ZN(N46853));
    INVX1 U33982 (.I(n32766), .ZN(N46854));
    NANDX1 U33983 (.A1(n34902), .A2(n32962), .ZN(N46855));
    INVX1 U33984 (.I(n33169), .ZN(N46856));
    NANDX1 U33985 (.A1(n21461), .A2(N239), .ZN(N46857));
    NANDX1 U33986 (.A1(n29710), .A2(N8409), .ZN(n46858));
    NOR2X1 U33987 (.A1(n32734), .A2(n40273), .ZN(N46859));
    NOR2X1 U33988 (.A1(N7088), .A2(n16128), .ZN(N46860));
    NOR2X1 U33989 (.A1(n40817), .A2(n17416), .ZN(n46861));
    NOR2X1 U33990 (.A1(n13136), .A2(n13564), .ZN(N46862));
    NOR2X1 U33991 (.A1(n13623), .A2(n28203), .ZN(N46863));
    NOR2X1 U33992 (.A1(n19165), .A2(n28143), .ZN(N46864));
    INVX1 U33993 (.I(n41611), .ZN(N46865));
    NOR2X1 U33994 (.A1(n14575), .A2(n20780), .ZN(N46866));
    NANDX1 U33995 (.A1(n37423), .A2(n41739), .ZN(N46867));
    NANDX1 U33996 (.A1(n27342), .A2(n29236), .ZN(N46868));
    NOR2X1 U33997 (.A1(n35750), .A2(n41686), .ZN(N46869));
    NANDX1 U33998 (.A1(n22230), .A2(n17554), .ZN(N46870));
    INVX1 U33999 (.I(n38357), .ZN(N46871));
    NOR2X1 U34000 (.A1(N5112), .A2(N1981), .ZN(N46872));
    NOR2X1 U34001 (.A1(N7927), .A2(n15544), .ZN(N46873));
    NOR2X1 U34002 (.A1(n21549), .A2(N275), .ZN(N46874));
    NOR2X1 U34003 (.A1(n30394), .A2(n28417), .ZN(N46875));
    NOR2X1 U34004 (.A1(n18212), .A2(N9861), .ZN(N46876));
    NANDX1 U34005 (.A1(n38991), .A2(N1069), .ZN(N46877));
    NOR2X1 U34006 (.A1(n26938), .A2(N3417), .ZN(N46878));
    INVX1 U34007 (.I(N12701), .ZN(N46879));
    NANDX1 U34008 (.A1(n32761), .A2(N594), .ZN(N46880));
    NOR2X1 U34009 (.A1(N11518), .A2(N7827), .ZN(N46881));
    INVX1 U34010 (.I(N6403), .ZN(N46882));
    NANDX1 U34011 (.A1(N5559), .A2(n41535), .ZN(N46883));
    NANDX1 U34012 (.A1(n13485), .A2(n13606), .ZN(N46884));
    INVX1 U34013 (.I(n24713), .ZN(N46885));
    NANDX1 U34014 (.A1(n42712), .A2(N11634), .ZN(N46886));
    NOR2X1 U34015 (.A1(n14177), .A2(n19525), .ZN(N46887));
    NANDX1 U34016 (.A1(N216), .A2(N4724), .ZN(N46888));
    NANDX1 U34017 (.A1(n13357), .A2(n31661), .ZN(N46889));
    NOR2X1 U34018 (.A1(N10368), .A2(n34041), .ZN(N46890));
    NANDX1 U34019 (.A1(n43128), .A2(n34634), .ZN(N46891));
    NANDX1 U34020 (.A1(N11173), .A2(n32140), .ZN(N46892));
    NOR2X1 U34021 (.A1(N7255), .A2(n16710), .ZN(N46893));
    NANDX1 U34022 (.A1(N5317), .A2(n30715), .ZN(N46894));
    NOR2X1 U34023 (.A1(n18923), .A2(n17522), .ZN(N46895));
    INVX1 U34024 (.I(n22482), .ZN(N46896));
    INVX1 U34025 (.I(n35238), .ZN(N46897));
    NOR2X1 U34026 (.A1(n20617), .A2(N11290), .ZN(N46898));
    INVX1 U34027 (.I(N10512), .ZN(N46899));
    INVX1 U34028 (.I(n41934), .ZN(N46900));
    NOR2X1 U34029 (.A1(N4201), .A2(n24142), .ZN(n46901));
    NANDX1 U34030 (.A1(n27921), .A2(n31504), .ZN(N46902));
    INVX1 U34031 (.I(N8762), .ZN(N46903));
    NANDX1 U34032 (.A1(n24423), .A2(n40901), .ZN(N46904));
    NANDX1 U34033 (.A1(n31678), .A2(n14139), .ZN(N46905));
    INVX1 U34034 (.I(n26674), .ZN(N46906));
    NANDX1 U34035 (.A1(n26653), .A2(N2124), .ZN(N46907));
    INVX1 U34036 (.I(n17104), .ZN(N46908));
    NOR2X1 U34037 (.A1(n25343), .A2(n42021), .ZN(N46909));
    NANDX1 U34038 (.A1(n35640), .A2(N9839), .ZN(N46910));
    NOR2X1 U34039 (.A1(N2679), .A2(n15531), .ZN(N46911));
    INVX1 U34040 (.I(n26547), .ZN(N46912));
    INVX1 U34041 (.I(n13752), .ZN(N46913));
    NANDX1 U34042 (.A1(n37332), .A2(n34935), .ZN(N46914));
    NOR2X1 U34043 (.A1(N2622), .A2(N12688), .ZN(N46915));
    NANDX1 U34044 (.A1(N50), .A2(n34402), .ZN(N46916));
    NANDX1 U34045 (.A1(N3868), .A2(n41523), .ZN(N46917));
    NOR2X1 U34046 (.A1(n38401), .A2(n24703), .ZN(N46918));
    NOR2X1 U34047 (.A1(N3511), .A2(n31486), .ZN(N46919));
    NANDX1 U34048 (.A1(n18533), .A2(n19715), .ZN(N46920));
    INVX1 U34049 (.I(N380), .ZN(N46921));
    NANDX1 U34050 (.A1(n28256), .A2(N3059), .ZN(N46922));
    NOR2X1 U34051 (.A1(N7546), .A2(n19285), .ZN(N46923));
    NOR2X1 U34052 (.A1(N10977), .A2(n26275), .ZN(N46924));
    INVX1 U34053 (.I(N2439), .ZN(N46925));
    INVX1 U34054 (.I(n30335), .ZN(N46926));
    INVX1 U34055 (.I(n37384), .ZN(n46927));
    INVX1 U34056 (.I(n39207), .ZN(N46928));
    NANDX1 U34057 (.A1(n23932), .A2(n37257), .ZN(N46929));
    NANDX1 U34058 (.A1(N8540), .A2(N8167), .ZN(n46930));
    NANDX1 U34059 (.A1(N1730), .A2(n29332), .ZN(N46931));
    INVX1 U34060 (.I(n20262), .ZN(N46932));
    INVX1 U34061 (.I(n35552), .ZN(N46933));
    INVX1 U34062 (.I(n24806), .ZN(N46934));
    NANDX1 U34063 (.A1(n13380), .A2(n16097), .ZN(N46935));
    INVX1 U34064 (.I(n32664), .ZN(N46936));
    NOR2X1 U34065 (.A1(n18217), .A2(N5146), .ZN(N46937));
    NOR2X1 U34066 (.A1(N10335), .A2(n41340), .ZN(n46938));
    NOR2X1 U34067 (.A1(n15140), .A2(n35251), .ZN(N46939));
    NANDX1 U34068 (.A1(N10874), .A2(N8238), .ZN(N46940));
    NOR2X1 U34069 (.A1(n37810), .A2(n30445), .ZN(N46941));
    INVX1 U34070 (.I(n35656), .ZN(N46942));
    NANDX1 U34071 (.A1(n31844), .A2(N11195), .ZN(n46943));
    NANDX1 U34072 (.A1(n41785), .A2(N6449), .ZN(n46944));
    NOR2X1 U34073 (.A1(N8634), .A2(n20934), .ZN(N46945));
    NANDX1 U34074 (.A1(N11693), .A2(n37030), .ZN(N46946));
    NANDX1 U34075 (.A1(N885), .A2(N36), .ZN(N46947));
    INVX1 U34076 (.I(N6030), .ZN(N46948));
    INVX1 U34077 (.I(N12100), .ZN(N46949));
    NOR2X1 U34078 (.A1(N11807), .A2(n27239), .ZN(N46950));
    NANDX1 U34079 (.A1(N9451), .A2(n38112), .ZN(N46951));
    NOR2X1 U34080 (.A1(n31026), .A2(n22129), .ZN(N46952));
    NANDX1 U34081 (.A1(N7348), .A2(N3992), .ZN(N46953));
    NOR2X1 U34082 (.A1(n28871), .A2(n15187), .ZN(N46954));
    NANDX1 U34083 (.A1(n27183), .A2(n21635), .ZN(N46955));
    NANDX1 U34084 (.A1(n25497), .A2(n42568), .ZN(N46956));
    INVX1 U34085 (.I(n37189), .ZN(N46957));
    NOR2X1 U34086 (.A1(N5568), .A2(n38073), .ZN(N46958));
    INVX1 U34087 (.I(N7334), .ZN(N46959));
    NOR2X1 U34088 (.A1(n39426), .A2(n19433), .ZN(N46960));
    NOR2X1 U34089 (.A1(n40912), .A2(n36352), .ZN(N46961));
    INVX1 U34090 (.I(n40042), .ZN(N46962));
    INVX1 U34091 (.I(n18818), .ZN(N46963));
    NANDX1 U34092 (.A1(n42800), .A2(n32534), .ZN(N46964));
    NANDX1 U34093 (.A1(N3319), .A2(n42661), .ZN(N46965));
    NANDX1 U34094 (.A1(N8185), .A2(N4171), .ZN(N46966));
    INVX1 U34095 (.I(n29819), .ZN(N46967));
    INVX1 U34096 (.I(N8907), .ZN(N46968));
    INVX1 U34097 (.I(n40938), .ZN(N46969));
    NANDX1 U34098 (.A1(n34080), .A2(N3033), .ZN(N46970));
    NANDX1 U34099 (.A1(n39280), .A2(N10366), .ZN(N46971));
    NANDX1 U34100 (.A1(n24913), .A2(n19479), .ZN(N46972));
    INVX1 U34101 (.I(n22353), .ZN(N46973));
    NOR2X1 U34102 (.A1(n19478), .A2(n18922), .ZN(n46974));
    INVX1 U34103 (.I(n38295), .ZN(N46975));
    NANDX1 U34104 (.A1(n22035), .A2(n17037), .ZN(N46976));
    INVX1 U34105 (.I(n25354), .ZN(N46977));
    INVX1 U34106 (.I(n17046), .ZN(N46978));
    INVX1 U34107 (.I(N10076), .ZN(N46979));
    INVX1 U34108 (.I(N9565), .ZN(N46980));
    NOR2X1 U34109 (.A1(n42514), .A2(n17839), .ZN(N46981));
    INVX1 U34110 (.I(n34816), .ZN(N46982));
    NOR2X1 U34111 (.A1(n39812), .A2(N11399), .ZN(N46983));
    NANDX1 U34112 (.A1(n39858), .A2(n21764), .ZN(N46984));
    NANDX1 U34113 (.A1(N5544), .A2(n38848), .ZN(N46985));
    INVX1 U34114 (.I(n17901), .ZN(n46986));
    INVX1 U34115 (.I(n39479), .ZN(N46987));
    NOR2X1 U34116 (.A1(n42827), .A2(n21883), .ZN(N46988));
    INVX1 U34117 (.I(n16391), .ZN(N46989));
    NOR2X1 U34118 (.A1(n34204), .A2(n22296), .ZN(N46990));
    NOR2X1 U34119 (.A1(n13949), .A2(n32371), .ZN(N46991));
    INVX1 U34120 (.I(n13193), .ZN(N46992));
    NOR2X1 U34121 (.A1(n14489), .A2(n20711), .ZN(N46993));
    NOR2X1 U34122 (.A1(n38985), .A2(n18836), .ZN(N46994));
    INVX1 U34123 (.I(N6911), .ZN(N46995));
    INVX1 U34124 (.I(n37076), .ZN(n46996));
    NOR2X1 U34125 (.A1(N653), .A2(n32299), .ZN(N46997));
    INVX1 U34126 (.I(n21209), .ZN(N46998));
    NANDX1 U34127 (.A1(N7942), .A2(N6895), .ZN(N46999));
    NANDX1 U34128 (.A1(n40448), .A2(n28777), .ZN(n47000));
    NOR2X1 U34129 (.A1(n13367), .A2(N3893), .ZN(N47001));
    NOR2X1 U34130 (.A1(n25342), .A2(n29205), .ZN(N47002));
    NOR2X1 U34131 (.A1(n14240), .A2(n34333), .ZN(N47003));
    NANDX1 U34132 (.A1(n32132), .A2(N5349), .ZN(N47004));
    NOR2X1 U34133 (.A1(n33011), .A2(n34013), .ZN(N47005));
    NOR2X1 U34134 (.A1(n30229), .A2(n30604), .ZN(N47006));
    INVX1 U34135 (.I(n13513), .ZN(N47007));
    INVX1 U34136 (.I(n21630), .ZN(N47008));
    NANDX1 U34137 (.A1(n31727), .A2(n42839), .ZN(N47009));
    NANDX1 U34138 (.A1(n39668), .A2(N6261), .ZN(N47010));
    NOR2X1 U34139 (.A1(n36643), .A2(n24718), .ZN(N47011));
    NOR2X1 U34140 (.A1(n39689), .A2(n18290), .ZN(N47012));
    NANDX1 U34141 (.A1(n21558), .A2(n37174), .ZN(N47013));
    NANDX1 U34142 (.A1(n25477), .A2(n28034), .ZN(N47014));
    NOR2X1 U34143 (.A1(N3816), .A2(n23063), .ZN(N47015));
    NOR2X1 U34144 (.A1(n36826), .A2(n13603), .ZN(N47016));
    NOR2X1 U34145 (.A1(n13263), .A2(n33886), .ZN(N47017));
    INVX1 U34146 (.I(n26775), .ZN(N47018));
    NANDX1 U34147 (.A1(N1538), .A2(n18793), .ZN(N47019));
    NOR2X1 U34148 (.A1(n34056), .A2(N7218), .ZN(N47020));
    NANDX1 U34149 (.A1(n29996), .A2(n22337), .ZN(N47021));
    INVX1 U34150 (.I(N11241), .ZN(n47022));
    INVX1 U34151 (.I(n25719), .ZN(N47023));
    NANDX1 U34152 (.A1(n29842), .A2(N3805), .ZN(N47024));
    NOR2X1 U34153 (.A1(n16588), .A2(n29281), .ZN(N47025));
    NOR2X1 U34154 (.A1(N2957), .A2(n33097), .ZN(N47026));
    NANDX1 U34155 (.A1(N9661), .A2(n16130), .ZN(N47027));
    NOR2X1 U34156 (.A1(N1743), .A2(n29392), .ZN(N47028));
    NANDX1 U34157 (.A1(n14803), .A2(N12694), .ZN(N47029));
    NANDX1 U34158 (.A1(n16340), .A2(n21167), .ZN(N47030));
    NANDX1 U34159 (.A1(n40075), .A2(n18064), .ZN(N47031));
    INVX1 U34160 (.I(n26598), .ZN(N47032));
    INVX1 U34161 (.I(n18836), .ZN(n47033));
    NOR2X1 U34162 (.A1(n26456), .A2(N1082), .ZN(N47034));
    INVX1 U34163 (.I(N2506), .ZN(N47035));
    NOR2X1 U34164 (.A1(n16167), .A2(N8773), .ZN(N47036));
    NOR2X1 U34165 (.A1(N3320), .A2(N11729), .ZN(N47037));
    INVX1 U34166 (.I(N3214), .ZN(N47038));
    INVX1 U34167 (.I(n19280), .ZN(N47039));
    NOR2X1 U34168 (.A1(N12812), .A2(n38352), .ZN(N47040));
    NANDX1 U34169 (.A1(n17294), .A2(n40725), .ZN(N47041));
    NOR2X1 U34170 (.A1(n33633), .A2(n18419), .ZN(N47042));
    INVX1 U34171 (.I(n19915), .ZN(N47043));
    INVX1 U34172 (.I(N8429), .ZN(N47044));
    NOR2X1 U34173 (.A1(n23091), .A2(n27264), .ZN(N47045));
    NANDX1 U34174 (.A1(n39226), .A2(n18026), .ZN(N47046));
    NANDX1 U34175 (.A1(n31411), .A2(N12591), .ZN(N47047));
    NOR2X1 U34176 (.A1(n40183), .A2(n26117), .ZN(N47048));
    INVX1 U34177 (.I(n41592), .ZN(N47049));
    NANDX1 U34178 (.A1(n35873), .A2(N9189), .ZN(N47050));
    NOR2X1 U34179 (.A1(N9112), .A2(N11680), .ZN(N47051));
    INVX1 U34180 (.I(n19413), .ZN(N47052));
    INVX1 U34181 (.I(n20038), .ZN(N47053));
    INVX1 U34182 (.I(N8814), .ZN(N47054));
    NANDX1 U34183 (.A1(n38298), .A2(n28729), .ZN(N47055));
    NOR2X1 U34184 (.A1(N3255), .A2(n21449), .ZN(N47056));
    NANDX1 U34185 (.A1(n30518), .A2(N8535), .ZN(n47057));
    INVX1 U34186 (.I(n38223), .ZN(N47058));
    INVX1 U34187 (.I(N7289), .ZN(N47059));
    NOR2X1 U34188 (.A1(n17896), .A2(n37151), .ZN(N47060));
    NOR2X1 U34189 (.A1(n40235), .A2(n35270), .ZN(N47061));
    NANDX1 U34190 (.A1(n22316), .A2(n34138), .ZN(N47062));
    INVX1 U34191 (.I(n31427), .ZN(N47063));
    NANDX1 U34192 (.A1(N5832), .A2(n40519), .ZN(N47064));
    NOR2X1 U34193 (.A1(n25869), .A2(n16249), .ZN(N47065));
    NANDX1 U34194 (.A1(N10533), .A2(N754), .ZN(N47066));
    NOR2X1 U34195 (.A1(N11039), .A2(N4008), .ZN(N47067));
    NOR2X1 U34196 (.A1(n34635), .A2(n24206), .ZN(N47068));
    NANDX1 U34197 (.A1(N10513), .A2(n18956), .ZN(N47069));
    NOR2X1 U34198 (.A1(N7481), .A2(n26297), .ZN(N47070));
    INVX1 U34199 (.I(N1159), .ZN(N47071));
    NANDX1 U34200 (.A1(N6984), .A2(n26109), .ZN(N47072));
    INVX1 U34201 (.I(n29299), .ZN(N47073));
    NOR2X1 U34202 (.A1(n41413), .A2(N6933), .ZN(N47074));
    NANDX1 U34203 (.A1(N3772), .A2(N3979), .ZN(N47075));
    INVX1 U34204 (.I(n19320), .ZN(N47076));
    NANDX1 U34205 (.A1(n28649), .A2(n19533), .ZN(N47077));
    INVX1 U34206 (.I(N12756), .ZN(N47078));
    INVX1 U34207 (.I(N4348), .ZN(N47079));
    NOR2X1 U34208 (.A1(n21734), .A2(n28553), .ZN(N47080));
    NANDX1 U34209 (.A1(n21926), .A2(n37188), .ZN(N47081));
    INVX1 U34210 (.I(n29406), .ZN(N47082));
    NOR2X1 U34211 (.A1(n34947), .A2(n20244), .ZN(N47083));
    INVX1 U34212 (.I(n41930), .ZN(N47084));
    INVX1 U34213 (.I(n20229), .ZN(n47085));
    INVX1 U34214 (.I(n42486), .ZN(N47086));
    NANDX1 U34215 (.A1(n24368), .A2(n40964), .ZN(N47087));
    INVX1 U34216 (.I(n28346), .ZN(N47088));
    INVX1 U34217 (.I(N10299), .ZN(N47089));
    NOR2X1 U34218 (.A1(n24977), .A2(n29831), .ZN(N47090));
    NOR2X1 U34219 (.A1(n37732), .A2(n16930), .ZN(N47091));
    INVX1 U34220 (.I(N12571), .ZN(N47092));
    NANDX1 U34221 (.A1(n17698), .A2(N1500), .ZN(N47093));
    NOR2X1 U34222 (.A1(N1094), .A2(n26225), .ZN(N47094));
    INVX1 U34223 (.I(N10786), .ZN(N47095));
    NOR2X1 U34224 (.A1(N2652), .A2(n16120), .ZN(N47096));
    INVX1 U34225 (.I(n28364), .ZN(N47097));
    NOR2X1 U34226 (.A1(n23271), .A2(n27377), .ZN(N47098));
    NANDX1 U34227 (.A1(n37318), .A2(n24868), .ZN(N47099));
    NANDX1 U34228 (.A1(N11871), .A2(n21196), .ZN(N47100));
    NOR2X1 U34229 (.A1(n39802), .A2(N2700), .ZN(N47101));
    NOR2X1 U34230 (.A1(n24601), .A2(n30112), .ZN(N47102));
    INVX1 U34231 (.I(n13746), .ZN(N47103));
    NANDX1 U34232 (.A1(N2671), .A2(n31444), .ZN(N47104));
    INVX1 U34233 (.I(n42618), .ZN(N47105));
    NANDX1 U34234 (.A1(n39446), .A2(n25026), .ZN(N47106));
    NOR2X1 U34235 (.A1(N3352), .A2(n17357), .ZN(N47107));
    INVX1 U34236 (.I(n42340), .ZN(N47108));
    NANDX1 U34237 (.A1(n31676), .A2(n22138), .ZN(N47109));
    NANDX1 U34238 (.A1(N11759), .A2(N5664), .ZN(N47110));
    NANDX1 U34239 (.A1(n26293), .A2(n17534), .ZN(N47111));
    NOR2X1 U34240 (.A1(N7653), .A2(N3544), .ZN(N47112));
    INVX1 U34241 (.I(N8524), .ZN(N47113));
    INVX1 U34242 (.I(N914), .ZN(n47114));
    NANDX1 U34243 (.A1(n31569), .A2(n33275), .ZN(N47115));
    INVX1 U34244 (.I(n19540), .ZN(N47116));
    NANDX1 U34245 (.A1(N7499), .A2(n41756), .ZN(n47117));
    NOR2X1 U34246 (.A1(n32524), .A2(n20965), .ZN(N47118));
    NOR2X1 U34247 (.A1(N6409), .A2(n26613), .ZN(N47119));
    NANDX1 U34248 (.A1(N8656), .A2(n14816), .ZN(N47120));
    NOR2X1 U34249 (.A1(n38280), .A2(n16254), .ZN(N47121));
    NOR2X1 U34250 (.A1(n38979), .A2(n42546), .ZN(N47122));
    NANDX1 U34251 (.A1(n17401), .A2(N6727), .ZN(N47123));
    NOR2X1 U34252 (.A1(n31675), .A2(N4930), .ZN(N47124));
    INVX1 U34253 (.I(n32588), .ZN(N47125));
    INVX1 U34254 (.I(n35372), .ZN(n47126));
    NOR2X1 U34255 (.A1(n39607), .A2(N1119), .ZN(N47127));
    NANDX1 U34256 (.A1(N3634), .A2(n32555), .ZN(N47128));
    INVX1 U34257 (.I(n25837), .ZN(N47129));
    INVX1 U34258 (.I(n37077), .ZN(N47130));
    NANDX1 U34259 (.A1(n36660), .A2(n38292), .ZN(N47131));
    INVX1 U34260 (.I(n41155), .ZN(n47132));
    INVX1 U34261 (.I(n25388), .ZN(N47133));
    NOR2X1 U34262 (.A1(n26547), .A2(N10574), .ZN(N47134));
    NANDX1 U34263 (.A1(N8983), .A2(n17654), .ZN(N47135));
    INVX1 U34264 (.I(n28115), .ZN(N47136));
    NANDX1 U34265 (.A1(N4026), .A2(n31917), .ZN(N47137));
    NOR2X1 U34266 (.A1(n24959), .A2(n23816), .ZN(N47138));
    NOR2X1 U34267 (.A1(n21093), .A2(n24935), .ZN(N47139));
    NANDX1 U34268 (.A1(n14406), .A2(n14017), .ZN(n47140));
    NANDX1 U34269 (.A1(n40243), .A2(n24063), .ZN(N47141));
    INVX1 U34270 (.I(n18695), .ZN(N47142));
    NANDX1 U34271 (.A1(n24648), .A2(N5803), .ZN(N47143));
    INVX1 U34272 (.I(n22179), .ZN(n47144));
    NANDX1 U34273 (.A1(N8229), .A2(N5253), .ZN(N47145));
    NOR2X1 U34274 (.A1(N10918), .A2(N3915), .ZN(N47146));
    NANDX1 U34275 (.A1(N10014), .A2(n32029), .ZN(N47147));
    NOR2X1 U34276 (.A1(n14039), .A2(n20474), .ZN(N47148));
    NOR2X1 U34277 (.A1(n38997), .A2(N817), .ZN(N47149));
    NOR2X1 U34278 (.A1(N6297), .A2(n15431), .ZN(N47150));
    INVX1 U34279 (.I(N10383), .ZN(N47151));
    NANDX1 U34280 (.A1(N9932), .A2(n40305), .ZN(N47152));
    NOR2X1 U34281 (.A1(n29440), .A2(n15527), .ZN(N47153));
    INVX1 U34282 (.I(N295), .ZN(n47154));
    INVX1 U34283 (.I(n34091), .ZN(N47155));
    INVX1 U34284 (.I(n31879), .ZN(N47156));
    NANDX1 U34285 (.A1(n27725), .A2(N9530), .ZN(N47157));
    NOR2X1 U34286 (.A1(n21319), .A2(N4834), .ZN(N47158));
    INVX1 U34287 (.I(N9876), .ZN(N47159));
    NOR2X1 U34288 (.A1(n23496), .A2(n30349), .ZN(N47160));
    NANDX1 U34289 (.A1(N8700), .A2(n20845), .ZN(N47161));
    NANDX1 U34290 (.A1(n14996), .A2(n25956), .ZN(N47162));
    INVX1 U34291 (.I(n25378), .ZN(N47163));
    INVX1 U34292 (.I(n16153), .ZN(N47164));
    NANDX1 U34293 (.A1(n24159), .A2(N2120), .ZN(N47165));
    NOR2X1 U34294 (.A1(n20486), .A2(n35566), .ZN(N47166));
    NOR2X1 U34295 (.A1(N784), .A2(n14566), .ZN(N47167));
    INVX1 U34296 (.I(n32783), .ZN(N47168));
    NOR2X1 U34297 (.A1(n36361), .A2(n32227), .ZN(n47169));
    NANDX1 U34298 (.A1(n30874), .A2(n41684), .ZN(N47170));
    INVX1 U34299 (.I(n16227), .ZN(N47171));
    INVX1 U34300 (.I(n39719), .ZN(N47172));
    NOR2X1 U34301 (.A1(n20086), .A2(N6772), .ZN(N47173));
    NANDX1 U34302 (.A1(n35081), .A2(n32727), .ZN(N47174));
    NANDX1 U34303 (.A1(N6667), .A2(n24016), .ZN(N47175));
    NOR2X1 U34304 (.A1(n28876), .A2(N4703), .ZN(N47176));
    NANDX1 U34305 (.A1(N2500), .A2(n14868), .ZN(N47177));
    NOR2X1 U34306 (.A1(n40925), .A2(n15651), .ZN(N47178));
    INVX1 U34307 (.I(n24285), .ZN(N47179));
    INVX1 U34308 (.I(n41744), .ZN(N47180));
    NOR2X1 U34309 (.A1(n26867), .A2(N8088), .ZN(N47181));
    NANDX1 U34310 (.A1(n14758), .A2(n17458), .ZN(N47182));
    NANDX1 U34311 (.A1(n26144), .A2(N3385), .ZN(n47183));
    NANDX1 U34312 (.A1(n35909), .A2(N10156), .ZN(N47184));
    INVX1 U34313 (.I(n17198), .ZN(N47185));
    NANDX1 U34314 (.A1(n35774), .A2(n23864), .ZN(N47186));
    NANDX1 U34315 (.A1(N3620), .A2(n42419), .ZN(N47187));
    NANDX1 U34316 (.A1(n17056), .A2(N1447), .ZN(N47188));
    NANDX1 U34317 (.A1(n22586), .A2(n42371), .ZN(N47189));
    NOR2X1 U34318 (.A1(n32360), .A2(N12863), .ZN(N47190));
    NOR2X1 U34319 (.A1(n30632), .A2(N9396), .ZN(N47191));
    INVX1 U34320 (.I(n28399), .ZN(N47192));
    NOR2X1 U34321 (.A1(n43309), .A2(N2384), .ZN(N47193));
    INVX1 U34322 (.I(n15661), .ZN(n47194));
    INVX1 U34323 (.I(N3874), .ZN(n47195));
    INVX1 U34324 (.I(N5603), .ZN(N47196));
    INVX1 U34325 (.I(n25294), .ZN(N47197));
    NANDX1 U34326 (.A1(n38975), .A2(n38837), .ZN(N47198));
    INVX1 U34327 (.I(n42594), .ZN(N47199));
    NANDX1 U34328 (.A1(n27795), .A2(n16178), .ZN(N47200));
    INVX1 U34329 (.I(n39829), .ZN(N47201));
    INVX1 U34330 (.I(n27808), .ZN(N47202));
    NANDX1 U34331 (.A1(N7010), .A2(n30351), .ZN(N47203));
    INVX1 U34332 (.I(n37641), .ZN(N47204));
    NANDX1 U34333 (.A1(N484), .A2(n22567), .ZN(N47205));
    NANDX1 U34334 (.A1(n33473), .A2(n14631), .ZN(N47206));
    NOR2X1 U34335 (.A1(N5661), .A2(N10078), .ZN(N47207));
    NOR2X1 U34336 (.A1(n13757), .A2(N5361), .ZN(N47208));
    NOR2X1 U34337 (.A1(n28731), .A2(n33204), .ZN(N47209));
    INVX1 U34338 (.I(n24095), .ZN(N47210));
    INVX1 U34339 (.I(n40774), .ZN(N47211));
    NANDX1 U34340 (.A1(n37835), .A2(N3159), .ZN(N47212));
    NOR2X1 U34341 (.A1(n34191), .A2(n31601), .ZN(N47213));
    NANDX1 U34342 (.A1(n27271), .A2(n38611), .ZN(N47214));
    NOR2X1 U34343 (.A1(n42675), .A2(n22459), .ZN(N47215));
    NANDX1 U34344 (.A1(n32839), .A2(n34706), .ZN(N47216));
    NOR2X1 U34345 (.A1(N12519), .A2(N5864), .ZN(N47217));
    NOR2X1 U34346 (.A1(n18179), .A2(N5621), .ZN(n47218));
    NOR2X1 U34347 (.A1(n21615), .A2(N10981), .ZN(N47219));
    NOR2X1 U34348 (.A1(n40025), .A2(n33865), .ZN(N47220));
    NOR2X1 U34349 (.A1(N10328), .A2(N432), .ZN(N47221));
    NOR2X1 U34350 (.A1(n18413), .A2(n38266), .ZN(N47222));
    INVX1 U34351 (.I(N11936), .ZN(N47223));
    NOR2X1 U34352 (.A1(n13954), .A2(n22946), .ZN(N47224));
    INVX1 U34353 (.I(n42244), .ZN(N47225));
    NANDX1 U34354 (.A1(n34817), .A2(n21230), .ZN(N47226));
    NOR2X1 U34355 (.A1(n13863), .A2(N2143), .ZN(N47227));
    NOR2X1 U34356 (.A1(n26381), .A2(n41158), .ZN(N47228));
    NOR2X1 U34357 (.A1(N1087), .A2(N3307), .ZN(N47229));
    NANDX1 U34358 (.A1(N12381), .A2(N3967), .ZN(N47230));
    NOR2X1 U34359 (.A1(N8934), .A2(n27511), .ZN(N47231));
    NOR2X1 U34360 (.A1(n19261), .A2(n27943), .ZN(N47232));
    NANDX1 U34361 (.A1(n27353), .A2(n22736), .ZN(n47233));
    INVX1 U34362 (.I(n39288), .ZN(N47234));
    NOR2X1 U34363 (.A1(N10040), .A2(N8441), .ZN(N47235));
    NOR2X1 U34364 (.A1(n41963), .A2(n18954), .ZN(N47236));
    INVX1 U34365 (.I(N9400), .ZN(N47237));
    NANDX1 U34366 (.A1(n28427), .A2(N11543), .ZN(N47238));
    INVX1 U34367 (.I(N11335), .ZN(N47239));
    INVX1 U34368 (.I(N7085), .ZN(N47240));
    NOR2X1 U34369 (.A1(N2214), .A2(n34739), .ZN(N47241));
    NANDX1 U34370 (.A1(n39333), .A2(n12954), .ZN(N47242));
    NANDX1 U34371 (.A1(n23371), .A2(n37174), .ZN(N47243));
    INVX1 U34372 (.I(N7841), .ZN(N47244));
    NANDX1 U34373 (.A1(n39067), .A2(n20257), .ZN(n47245));
    NANDX1 U34374 (.A1(n24563), .A2(n41016), .ZN(N47246));
    NOR2X1 U34375 (.A1(n33003), .A2(n31084), .ZN(N47247));
    NOR2X1 U34376 (.A1(n41637), .A2(n35329), .ZN(N47248));
    INVX1 U34377 (.I(N11472), .ZN(N47249));
    INVX1 U34378 (.I(N12352), .ZN(N47250));
    NOR2X1 U34379 (.A1(n21298), .A2(N11259), .ZN(N47251));
    INVX1 U34380 (.I(n13078), .ZN(N47252));
    NANDX1 U34381 (.A1(n36591), .A2(N6919), .ZN(N47253));
    INVX1 U34382 (.I(N6073), .ZN(N47254));
    INVX1 U34383 (.I(n22383), .ZN(N47255));
    INVX1 U34384 (.I(n21407), .ZN(N47256));
    NOR2X1 U34385 (.A1(n30040), .A2(N6682), .ZN(N47257));
    NANDX1 U34386 (.A1(n12921), .A2(n31244), .ZN(N47258));
    NOR2X1 U34387 (.A1(N5840), .A2(N10454), .ZN(N47259));
    INVX1 U34388 (.I(n30402), .ZN(N47260));
    INVX1 U34389 (.I(n40002), .ZN(N47261));
    NANDX1 U34390 (.A1(N9770), .A2(N6493), .ZN(N47262));
    NOR2X1 U34391 (.A1(n25178), .A2(n17470), .ZN(N47263));
    NANDX1 U34392 (.A1(n27030), .A2(n30547), .ZN(N47264));
    NOR2X1 U34393 (.A1(n20148), .A2(n27146), .ZN(n47265));
    INVX1 U34394 (.I(n15900), .ZN(N47266));
    INVX1 U34395 (.I(n38087), .ZN(N47267));
    NANDX1 U34396 (.A1(N4453), .A2(N4198), .ZN(N47268));
    INVX1 U34397 (.I(N11134), .ZN(N47269));
    NOR2X1 U34398 (.A1(n27673), .A2(n42377), .ZN(N47270));
    NOR2X1 U34399 (.A1(n23192), .A2(n42510), .ZN(N47271));
    INVX1 U34400 (.I(N10121), .ZN(N47272));
    NANDX1 U34401 (.A1(n31662), .A2(n31011), .ZN(N47273));
    NANDX1 U34402 (.A1(n27834), .A2(N10460), .ZN(N47274));
    NOR2X1 U34403 (.A1(N1831), .A2(n34320), .ZN(N47275));
    NOR2X1 U34404 (.A1(n22057), .A2(n17859), .ZN(N47276));
    NOR2X1 U34405 (.A1(N5730), .A2(N411), .ZN(N47277));
    INVX1 U34406 (.I(n32248), .ZN(N47278));
    NOR2X1 U34407 (.A1(n26278), .A2(n36700), .ZN(N47279));
    INVX1 U34408 (.I(n41030), .ZN(N47280));
    INVX1 U34409 (.I(n22938), .ZN(N47281));
    NOR2X1 U34410 (.A1(N3265), .A2(n20244), .ZN(N47282));
    INVX1 U34411 (.I(n35454), .ZN(N47283));
    INVX1 U34412 (.I(n37902), .ZN(N47284));
    INVX1 U34413 (.I(N92), .ZN(N47285));
    NANDX1 U34414 (.A1(N6741), .A2(n27925), .ZN(N47286));
    NOR2X1 U34415 (.A1(n28702), .A2(n19435), .ZN(N47287));
    NOR2X1 U34416 (.A1(n23900), .A2(n41492), .ZN(N47288));
    NANDX1 U34417 (.A1(n39246), .A2(n36901), .ZN(N47289));
    NOR2X1 U34418 (.A1(n27019), .A2(n25676), .ZN(N47290));
    NANDX1 U34419 (.A1(n42976), .A2(n18903), .ZN(N47291));
    NOR2X1 U34420 (.A1(n40534), .A2(n23263), .ZN(N47292));
    INVX1 U34421 (.I(N11971), .ZN(N47293));
    NOR2X1 U34422 (.A1(n30841), .A2(n39752), .ZN(N47294));
    NOR2X1 U34423 (.A1(n42743), .A2(n34182), .ZN(N47295));
    INVX1 U34424 (.I(n42835), .ZN(N47296));
    NOR2X1 U34425 (.A1(n37398), .A2(n16967), .ZN(N47297));
    NANDX1 U34426 (.A1(n22627), .A2(n36402), .ZN(N47298));
    NOR2X1 U34427 (.A1(n36207), .A2(n24101), .ZN(N47299));
    INVX1 U34428 (.I(n31980), .ZN(N47300));
    INVX1 U34429 (.I(n34256), .ZN(N47301));
    INVX1 U34430 (.I(n43205), .ZN(N47302));
    NANDX1 U34431 (.A1(n15029), .A2(n18635), .ZN(N47303));
    NANDX1 U34432 (.A1(N1770), .A2(n31578), .ZN(N47304));
    NANDX1 U34433 (.A1(N3421), .A2(N4312), .ZN(N47305));
    NANDX1 U34434 (.A1(n43172), .A2(N2180), .ZN(N47306));
    INVX1 U34435 (.I(n23561), .ZN(N47307));
    INVX1 U34436 (.I(N6952), .ZN(N47308));
    NOR2X1 U34437 (.A1(n37082), .A2(n13599), .ZN(N47309));
    NOR2X1 U34438 (.A1(N5916), .A2(N6528), .ZN(N47310));
    NANDX1 U34439 (.A1(n42122), .A2(n20308), .ZN(N47311));
    NOR2X1 U34440 (.A1(n30629), .A2(n37836), .ZN(N47312));
    NOR2X1 U34441 (.A1(n35834), .A2(n37568), .ZN(N47313));
    NANDX1 U34442 (.A1(n40543), .A2(N2411), .ZN(N47314));
    NOR2X1 U34443 (.A1(n42312), .A2(n33988), .ZN(N47315));
    NANDX1 U34444 (.A1(n35412), .A2(n27979), .ZN(N47316));
    INVX1 U34445 (.I(n35112), .ZN(N47317));
    NOR2X1 U34446 (.A1(N9700), .A2(n15200), .ZN(N47318));
    INVX1 U34447 (.I(N6332), .ZN(N47319));
    NANDX1 U34448 (.A1(N2812), .A2(n19930), .ZN(N47320));
    INVX1 U34449 (.I(n41879), .ZN(N47321));
    NANDX1 U34450 (.A1(n15749), .A2(n40529), .ZN(N47322));
    NOR2X1 U34451 (.A1(N8230), .A2(n17365), .ZN(N47323));
    NANDX1 U34452 (.A1(n14326), .A2(n42879), .ZN(N47324));
    NANDX1 U34453 (.A1(N9964), .A2(n29629), .ZN(N47325));
    NANDX1 U34454 (.A1(n15956), .A2(n18148), .ZN(N47326));
    NANDX1 U34455 (.A1(N9747), .A2(N10088), .ZN(N47327));
    INVX1 U34456 (.I(N11857), .ZN(N47328));
    INVX1 U34457 (.I(n34684), .ZN(N47329));
    NANDX1 U34458 (.A1(N6606), .A2(N10734), .ZN(N47330));
    NANDX1 U34459 (.A1(n30555), .A2(N3225), .ZN(N47331));
    INVX1 U34460 (.I(n30550), .ZN(N47332));
    NANDX1 U34461 (.A1(n43312), .A2(n35978), .ZN(n47333));
    NANDX1 U34462 (.A1(n25963), .A2(n33887), .ZN(n47334));
    NANDX1 U34463 (.A1(N2978), .A2(N4740), .ZN(N47335));
    NOR2X1 U34464 (.A1(N7240), .A2(N4383), .ZN(N47336));
    INVX1 U34465 (.I(n13912), .ZN(N47337));
    NANDX1 U34466 (.A1(n42594), .A2(n33931), .ZN(N47338));
    NOR2X1 U34467 (.A1(N9209), .A2(N5304), .ZN(N47339));
    INVX1 U34468 (.I(N615), .ZN(N47340));
    INVX1 U34469 (.I(n32536), .ZN(N47341));
    NOR2X1 U34470 (.A1(n40401), .A2(N6630), .ZN(N47342));
    NOR2X1 U34471 (.A1(N154), .A2(n33806), .ZN(N47343));
    NOR2X1 U34472 (.A1(N1785), .A2(n23325), .ZN(N47344));
    INVX1 U34473 (.I(n33624), .ZN(N47345));
    NOR2X1 U34474 (.A1(n30604), .A2(n29035), .ZN(N47346));
    INVX1 U34475 (.I(n25024), .ZN(N47347));
    NOR2X1 U34476 (.A1(n38864), .A2(n29406), .ZN(N47348));
    INVX1 U34477 (.I(N9303), .ZN(N47349));
    NANDX1 U34478 (.A1(n16459), .A2(n32913), .ZN(N47350));
    INVX1 U34479 (.I(n15347), .ZN(N47351));
    NOR2X1 U34480 (.A1(n37015), .A2(n15961), .ZN(N47352));
    INVX1 U34481 (.I(n15758), .ZN(N47353));
    NANDX1 U34482 (.A1(n21340), .A2(n22387), .ZN(N47354));
    NANDX1 U34483 (.A1(N11173), .A2(N2400), .ZN(N47355));
    INVX1 U34484 (.I(N2637), .ZN(N47356));
    NANDX1 U34485 (.A1(n41243), .A2(n25940), .ZN(N47357));
    NANDX1 U34486 (.A1(n28375), .A2(N1182), .ZN(N47358));
    NANDX1 U34487 (.A1(n43078), .A2(n14714), .ZN(N47359));
    NANDX1 U34488 (.A1(n29011), .A2(n32052), .ZN(N47360));
    NOR2X1 U34489 (.A1(n14642), .A2(N5038), .ZN(N47361));
    NOR2X1 U34490 (.A1(n20037), .A2(n20385), .ZN(N47362));
    NOR2X1 U34491 (.A1(N3259), .A2(n26025), .ZN(N47363));
    INVX1 U34492 (.I(n19016), .ZN(N47364));
    NOR2X1 U34493 (.A1(n23358), .A2(n41402), .ZN(N47365));
    INVX1 U34494 (.I(n34530), .ZN(N47366));
    NOR2X1 U34495 (.A1(n36781), .A2(n26846), .ZN(N47367));
    INVX1 U34496 (.I(n34551), .ZN(N47368));
    NOR2X1 U34497 (.A1(n36953), .A2(N9133), .ZN(N47369));
    INVX1 U34498 (.I(N2852), .ZN(N47370));
    NOR2X1 U34499 (.A1(n14888), .A2(N7614), .ZN(N47371));
    NOR2X1 U34500 (.A1(N3467), .A2(n21678), .ZN(N47372));
    NOR2X1 U34501 (.A1(N8504), .A2(n14862), .ZN(N47373));
    NANDX1 U34502 (.A1(n18568), .A2(N2789), .ZN(N47374));
    NOR2X1 U34503 (.A1(n34273), .A2(N4807), .ZN(n47375));
    NOR2X1 U34504 (.A1(n29685), .A2(n28164), .ZN(N47376));
    INVX1 U34505 (.I(N11620), .ZN(n47377));
    INVX1 U34506 (.I(n41358), .ZN(N47378));
    INVX1 U34507 (.I(n35746), .ZN(N47379));
    INVX1 U34508 (.I(n29158), .ZN(N47380));
    NOR2X1 U34509 (.A1(n40251), .A2(n27971), .ZN(N47381));
    NANDX1 U34510 (.A1(n43102), .A2(n26388), .ZN(N47382));
    INVX1 U34511 (.I(N7243), .ZN(N47383));
    NANDX1 U34512 (.A1(n20113), .A2(n18600), .ZN(N47384));
    NOR2X1 U34513 (.A1(n18296), .A2(n33461), .ZN(N47385));
    NANDX1 U34514 (.A1(n26544), .A2(n25929), .ZN(N47386));
    NOR2X1 U34515 (.A1(n17344), .A2(n30736), .ZN(N47387));
    NANDX1 U34516 (.A1(n36708), .A2(n15427), .ZN(N47388));
    NOR2X1 U34517 (.A1(n38007), .A2(n14008), .ZN(N47389));
    NOR2X1 U34518 (.A1(n32614), .A2(N6281), .ZN(N47390));
    NOR2X1 U34519 (.A1(N7980), .A2(n41019), .ZN(N47391));
    NANDX1 U34520 (.A1(n25630), .A2(n32458), .ZN(N47392));
    NANDX1 U34521 (.A1(N8545), .A2(N5632), .ZN(N47393));
    INVX1 U34522 (.I(n41721), .ZN(N47394));
    INVX1 U34523 (.I(n18480), .ZN(N47395));
    NOR2X1 U34524 (.A1(n33719), .A2(n41620), .ZN(N47396));
    INVX1 U34525 (.I(N6470), .ZN(N47397));
    NOR2X1 U34526 (.A1(N6054), .A2(n13493), .ZN(N47398));
    NANDX1 U34527 (.A1(N3547), .A2(n39881), .ZN(N47399));
    INVX1 U34528 (.I(N8915), .ZN(N47400));
    NANDX1 U34529 (.A1(n20133), .A2(N12169), .ZN(N47401));
    NOR2X1 U34530 (.A1(n26414), .A2(n18720), .ZN(N47402));
    NOR2X1 U34531 (.A1(n13640), .A2(n22050), .ZN(N47403));
    NOR2X1 U34532 (.A1(N2625), .A2(n14688), .ZN(N47404));
    NOR2X1 U34533 (.A1(n41408), .A2(n14569), .ZN(N47405));
    NANDX1 U34534 (.A1(n13359), .A2(n22728), .ZN(N47406));
    NANDX1 U34535 (.A1(n36757), .A2(N10556), .ZN(N47407));
    INVX1 U34536 (.I(n43227), .ZN(N47408));
    NOR2X1 U34537 (.A1(n23467), .A2(N2927), .ZN(N47409));
    INVX1 U34538 (.I(n16693), .ZN(N47410));
    NANDX1 U34539 (.A1(n31456), .A2(n15288), .ZN(N47411));
    INVX1 U34540 (.I(N8117), .ZN(N47412));
    NANDX1 U34541 (.A1(N3514), .A2(n24210), .ZN(N47413));
    NANDX1 U34542 (.A1(n24729), .A2(n37849), .ZN(N47414));
    NOR2X1 U34543 (.A1(n28101), .A2(n30153), .ZN(N47415));
    NOR2X1 U34544 (.A1(n29697), .A2(n17768), .ZN(N47416));
    INVX1 U34545 (.I(n19222), .ZN(N47417));
    NANDX1 U34546 (.A1(N2303), .A2(n18127), .ZN(N47418));
    NANDX1 U34547 (.A1(N2538), .A2(n35540), .ZN(n47419));
    NANDX1 U34548 (.A1(n26849), .A2(N5215), .ZN(N47420));
    NOR2X1 U34549 (.A1(N8707), .A2(n21907), .ZN(N47421));
    INVX1 U34550 (.I(n40163), .ZN(N47422));
    NANDX1 U34551 (.A1(n29214), .A2(N4807), .ZN(N47423));
    NOR2X1 U34552 (.A1(n32727), .A2(n29016), .ZN(N47424));
    NOR2X1 U34553 (.A1(n13983), .A2(n13072), .ZN(N47425));
    NANDX1 U34554 (.A1(n42083), .A2(n32904), .ZN(N47426));
    INVX1 U34555 (.I(n17988), .ZN(N47427));
    NANDX1 U34556 (.A1(n28557), .A2(n37209), .ZN(N47428));
    NOR2X1 U34557 (.A1(n20540), .A2(N1543), .ZN(N47429));
    NANDX1 U34558 (.A1(n23077), .A2(n26763), .ZN(N47430));
    INVX1 U34559 (.I(N6454), .ZN(n47431));
    NANDX1 U34560 (.A1(N8595), .A2(N4840), .ZN(N47432));
    NOR2X1 U34561 (.A1(N4059), .A2(N1530), .ZN(N47433));
    NOR2X1 U34562 (.A1(n33273), .A2(N6336), .ZN(N47434));
    NANDX1 U34563 (.A1(n22527), .A2(n25031), .ZN(N47435));
    INVX1 U34564 (.I(n36510), .ZN(N47436));
    NOR2X1 U34565 (.A1(n29963), .A2(n24800), .ZN(N47437));
    NANDX1 U34566 (.A1(n25152), .A2(n32467), .ZN(N47438));
    NOR2X1 U34567 (.A1(n43389), .A2(n15883), .ZN(N47439));
    NOR2X1 U34568 (.A1(n20456), .A2(n17426), .ZN(N47440));
    NANDX1 U34569 (.A1(n33212), .A2(n33868), .ZN(N47441));
    NANDX1 U34570 (.A1(n39665), .A2(N12052), .ZN(N47442));
    NANDX1 U34571 (.A1(N1033), .A2(N1822), .ZN(N47443));
    NANDX1 U34572 (.A1(n35714), .A2(n18466), .ZN(N47444));
    INVX1 U34573 (.I(n31730), .ZN(N47445));
    NOR2X1 U34574 (.A1(n24366), .A2(n13288), .ZN(N47446));
    INVX1 U34575 (.I(N7083), .ZN(N47447));
    INVX1 U34576 (.I(N1276), .ZN(N47448));
    NANDX1 U34577 (.A1(n14810), .A2(n26428), .ZN(N47449));
    INVX1 U34578 (.I(n39221), .ZN(N47450));
    INVX1 U34579 (.I(n26439), .ZN(n47451));
    NANDX1 U34580 (.A1(n36479), .A2(n33544), .ZN(N47452));
    NOR2X1 U34581 (.A1(n26218), .A2(n23939), .ZN(N47453));
    NANDX1 U34582 (.A1(N12091), .A2(n35990), .ZN(n47454));
    NOR2X1 U34583 (.A1(N2803), .A2(n37812), .ZN(N47455));
    NANDX1 U34584 (.A1(n38516), .A2(N12805), .ZN(N47456));
    NOR2X1 U34585 (.A1(n26773), .A2(n38131), .ZN(N47457));
    INVX1 U34586 (.I(n29741), .ZN(N47458));
    INVX1 U34587 (.I(n33982), .ZN(N47459));
    NANDX1 U34588 (.A1(N10720), .A2(N1752), .ZN(N47460));
    NOR2X1 U34589 (.A1(n37147), .A2(N12308), .ZN(N47461));
    NANDX1 U34590 (.A1(N9698), .A2(n28426), .ZN(N47462));
    NANDX1 U34591 (.A1(N2704), .A2(n18498), .ZN(N47463));
    INVX1 U34592 (.I(n18602), .ZN(N47464));
    INVX1 U34593 (.I(n37706), .ZN(N47465));
    NOR2X1 U34594 (.A1(n24634), .A2(N3531), .ZN(N47466));
    NANDX1 U34595 (.A1(N8653), .A2(n14547), .ZN(N47467));
    NOR2X1 U34596 (.A1(N11137), .A2(n27402), .ZN(N47468));
    NOR2X1 U34597 (.A1(N5796), .A2(N10829), .ZN(N47469));
    INVX1 U34598 (.I(n15240), .ZN(N47470));
    NOR2X1 U34599 (.A1(n37955), .A2(n15639), .ZN(n47471));
    INVX1 U34600 (.I(n15989), .ZN(N47472));
    INVX1 U34601 (.I(n38229), .ZN(N47473));
    NANDX1 U34602 (.A1(N8691), .A2(n23182), .ZN(N47474));
    NOR2X1 U34603 (.A1(N11395), .A2(n31359), .ZN(n47475));
    INVX1 U34604 (.I(n29996), .ZN(N47476));
    INVX1 U34605 (.I(N11376), .ZN(N47477));
    NANDX1 U34606 (.A1(N1164), .A2(n14907), .ZN(N47478));
    INVX1 U34607 (.I(n42968), .ZN(N47479));
    NOR2X1 U34608 (.A1(n15132), .A2(N10632), .ZN(N47480));
    NANDX1 U34609 (.A1(N6329), .A2(N6107), .ZN(N47481));
    NOR2X1 U34610 (.A1(n27266), .A2(N11026), .ZN(N47482));
    NANDX1 U34611 (.A1(N11428), .A2(n26665), .ZN(N47483));
    NOR2X1 U34612 (.A1(n17097), .A2(n25658), .ZN(N47484));
    NANDX1 U34613 (.A1(n40020), .A2(n34348), .ZN(N47485));
    NANDX1 U34614 (.A1(N10455), .A2(N2270), .ZN(N47486));
    NANDX1 U34615 (.A1(n27597), .A2(n21945), .ZN(N47487));
    NOR2X1 U34616 (.A1(n38973), .A2(n28839), .ZN(N47488));
    NOR2X1 U34617 (.A1(N87), .A2(n25754), .ZN(N47489));
    NOR2X1 U34618 (.A1(N8899), .A2(n30566), .ZN(N47490));
    NANDX1 U34619 (.A1(N1641), .A2(n36894), .ZN(N47491));
    NANDX1 U34620 (.A1(n38363), .A2(N10368), .ZN(N47492));
    NOR2X1 U34621 (.A1(N12311), .A2(N11475), .ZN(N47493));
    NANDX1 U34622 (.A1(N12180), .A2(n28571), .ZN(N47494));
    NANDX1 U34623 (.A1(n17125), .A2(n14798), .ZN(n47495));
    NOR2X1 U34624 (.A1(n34931), .A2(n25252), .ZN(N47496));
    INVX1 U34625 (.I(n40624), .ZN(N47497));
    NOR2X1 U34626 (.A1(N3624), .A2(n22847), .ZN(N47498));
    INVX1 U34627 (.I(n32462), .ZN(n47499));
    NANDX1 U34628 (.A1(n38115), .A2(N4424), .ZN(N47500));
    NANDX1 U34629 (.A1(n36693), .A2(n34989), .ZN(N47501));
    NANDX1 U34630 (.A1(n38333), .A2(n18090), .ZN(N47502));
    NOR2X1 U34631 (.A1(n22903), .A2(n18137), .ZN(N47503));
    NANDX1 U34632 (.A1(n24893), .A2(n29612), .ZN(N47504));
    NANDX1 U34633 (.A1(n37072), .A2(n14710), .ZN(N47505));
    NOR2X1 U34634 (.A1(N10724), .A2(n29508), .ZN(N47506));
    NOR2X1 U34635 (.A1(n35335), .A2(N11287), .ZN(N47507));
    INVX1 U34636 (.I(n32486), .ZN(N47508));
    NOR2X1 U34637 (.A1(n20979), .A2(N11861), .ZN(n47509));
    NOR2X1 U34638 (.A1(n43120), .A2(N7773), .ZN(N47510));
    NANDX1 U34639 (.A1(n37223), .A2(n19719), .ZN(N47511));
    NOR2X1 U34640 (.A1(n18419), .A2(n14857), .ZN(N47512));
    INVX1 U34641 (.I(n36509), .ZN(N47513));
    NOR2X1 U34642 (.A1(n23037), .A2(N11173), .ZN(n47514));
    NANDX1 U34643 (.A1(N4457), .A2(n40784), .ZN(N47515));
    NOR2X1 U34644 (.A1(n31209), .A2(N1702), .ZN(n47516));
    INVX1 U34645 (.I(n31612), .ZN(N47517));
    NOR2X1 U34646 (.A1(n25829), .A2(n23474), .ZN(N47518));
    NOR2X1 U34647 (.A1(n43184), .A2(N12488), .ZN(N47519));
    INVX1 U34648 (.I(n20690), .ZN(N47520));
    NANDX1 U34649 (.A1(n37096), .A2(N10018), .ZN(N47521));
    NOR2X1 U34650 (.A1(n15997), .A2(N3768), .ZN(N47522));
    INVX1 U34651 (.I(n31590), .ZN(N47523));
    NANDX1 U34652 (.A1(n12902), .A2(n31723), .ZN(N47524));
    NANDX1 U34653 (.A1(N1875), .A2(N11287), .ZN(N47525));
    NANDX1 U34654 (.A1(n41914), .A2(N5424), .ZN(N47526));
    NANDX1 U34655 (.A1(N8950), .A2(n36632), .ZN(N47527));
    NANDX1 U34656 (.A1(n42574), .A2(n24771), .ZN(N47528));
    INVX1 U34657 (.I(n24931), .ZN(N47529));
    INVX1 U34658 (.I(n37190), .ZN(N47530));
    INVX1 U34659 (.I(N6940), .ZN(N47531));
    INVX1 U34660 (.I(n35012), .ZN(N47532));
    INVX1 U34661 (.I(N9219), .ZN(N47533));
    NOR2X1 U34662 (.A1(N9614), .A2(n14895), .ZN(N47534));
    INVX1 U34663 (.I(N7660), .ZN(n47535));
    NANDX1 U34664 (.A1(N6870), .A2(n20561), .ZN(N47536));
    NANDX1 U34665 (.A1(N1452), .A2(n22436), .ZN(N47537));
    NOR2X1 U34666 (.A1(n40359), .A2(n20877), .ZN(N47538));
    NOR2X1 U34667 (.A1(n22785), .A2(n29826), .ZN(N47539));
    NOR2X1 U34668 (.A1(N6912), .A2(n18608), .ZN(N47540));
    NOR2X1 U34669 (.A1(N11927), .A2(n33218), .ZN(N47541));
    NOR2X1 U34670 (.A1(N5644), .A2(N4067), .ZN(N47542));
    NANDX1 U34671 (.A1(n21239), .A2(n28758), .ZN(N47543));
    NOR2X1 U34672 (.A1(n20137), .A2(n19994), .ZN(N47544));
    INVX1 U34673 (.I(n35031), .ZN(N47545));
    INVX1 U34674 (.I(n13931), .ZN(n47546));
    NOR2X1 U34675 (.A1(N1227), .A2(n34491), .ZN(N47547));
    NANDX1 U34676 (.A1(N2679), .A2(n13454), .ZN(N47548));
    INVX1 U34677 (.I(n32717), .ZN(N47549));
    NANDX1 U34678 (.A1(n23566), .A2(N12029), .ZN(N47550));
    NANDX1 U34679 (.A1(n26888), .A2(n18940), .ZN(N47551));
    INVX1 U34680 (.I(N1189), .ZN(N47552));
    NANDX1 U34681 (.A1(n41548), .A2(n13413), .ZN(N47553));
    INVX1 U34682 (.I(n35294), .ZN(N47554));
    NANDX1 U34683 (.A1(n37107), .A2(n20580), .ZN(N47555));
    INVX1 U34684 (.I(n13771), .ZN(N47556));
    NOR2X1 U34685 (.A1(n25185), .A2(n38481), .ZN(N47557));
    INVX1 U34686 (.I(n28795), .ZN(N47558));
    INVX1 U34687 (.I(n36157), .ZN(N47559));
    NOR2X1 U34688 (.A1(n33585), .A2(n28515), .ZN(N47560));
    INVX1 U34689 (.I(N3515), .ZN(N47561));
    NOR2X1 U34690 (.A1(n36637), .A2(n16761), .ZN(N47562));
    INVX1 U34691 (.I(n26360), .ZN(N47563));
    NANDX1 U34692 (.A1(n38406), .A2(n34690), .ZN(N47564));
    NANDX1 U34693 (.A1(n15479), .A2(n22445), .ZN(N47565));
    INVX1 U34694 (.I(n31347), .ZN(N47566));
    NOR2X1 U34695 (.A1(n16393), .A2(n24982), .ZN(N47567));
    NANDX1 U34696 (.A1(n35306), .A2(n28432), .ZN(N47568));
    NOR2X1 U34697 (.A1(N6699), .A2(n13121), .ZN(N47569));
    NOR2X1 U34698 (.A1(n35493), .A2(n15210), .ZN(N47570));
    NOR2X1 U34699 (.A1(N1514), .A2(N5322), .ZN(N47571));
    INVX1 U34700 (.I(n14141), .ZN(N47572));
    INVX1 U34701 (.I(n31399), .ZN(N47573));
    INVX1 U34702 (.I(n15277), .ZN(N47574));
    INVX1 U34703 (.I(n23344), .ZN(N47575));
    INVX1 U34704 (.I(n35478), .ZN(N47576));
    INVX1 U34705 (.I(N6496), .ZN(N47577));
    NANDX1 U34706 (.A1(n26685), .A2(N632), .ZN(N47578));
    NOR2X1 U34707 (.A1(n30630), .A2(N6704), .ZN(N47579));
    NOR2X1 U34708 (.A1(N11683), .A2(n42009), .ZN(N47580));
    INVX1 U34709 (.I(n22988), .ZN(N47581));
    INVX1 U34710 (.I(n30931), .ZN(N47582));
    NANDX1 U34711 (.A1(n30408), .A2(N2669), .ZN(N47583));
    NOR2X1 U34712 (.A1(n31921), .A2(N7990), .ZN(N47584));
    INVX1 U34713 (.I(n35741), .ZN(N47585));
    INVX1 U34714 (.I(N12444), .ZN(N47586));
    INVX1 U34715 (.I(N11462), .ZN(N47587));
    NANDX1 U34716 (.A1(N12596), .A2(n26914), .ZN(N47588));
    NANDX1 U34717 (.A1(n16836), .A2(n23089), .ZN(N47589));
    NOR2X1 U34718 (.A1(n33200), .A2(n13400), .ZN(N47590));
    NOR2X1 U34719 (.A1(n20358), .A2(n20103), .ZN(N47591));
    NANDX1 U34720 (.A1(n21720), .A2(N8319), .ZN(N47592));
    NOR2X1 U34721 (.A1(n34387), .A2(N3234), .ZN(N47593));
    INVX1 U34722 (.I(N6344), .ZN(N47594));
    NANDX1 U34723 (.A1(n14191), .A2(n17220), .ZN(N47595));
    INVX1 U34724 (.I(N11861), .ZN(N47596));
    NANDX1 U34725 (.A1(N4038), .A2(N8046), .ZN(N47597));
    NOR2X1 U34726 (.A1(n36762), .A2(n19508), .ZN(N47598));
    NANDX1 U34727 (.A1(N5886), .A2(n36101), .ZN(N47599));
    INVX1 U34728 (.I(N12401), .ZN(N47600));
    NANDX1 U34729 (.A1(N10109), .A2(N2129), .ZN(N47601));
    INVX1 U34730 (.I(n26983), .ZN(N47602));
    NANDX1 U34731 (.A1(n28578), .A2(n33237), .ZN(N47603));
    INVX1 U34732 (.I(n26576), .ZN(N47604));
    NOR2X1 U34733 (.A1(n24799), .A2(n29809), .ZN(N47605));
    NOR2X1 U34734 (.A1(n31142), .A2(n19977), .ZN(N47606));
    INVX1 U34735 (.I(n38042), .ZN(N47607));
    NANDX1 U34736 (.A1(n30762), .A2(n36306), .ZN(N47608));
    NANDX1 U34737 (.A1(n38807), .A2(n36693), .ZN(N47609));
    NOR2X1 U34738 (.A1(n14842), .A2(N3123), .ZN(N47610));
    NANDX1 U34739 (.A1(n40622), .A2(n14547), .ZN(n47611));
    NANDX1 U34740 (.A1(N2546), .A2(n14335), .ZN(N47612));
    NANDX1 U34741 (.A1(N11021), .A2(n30997), .ZN(N47613));
    NOR2X1 U34742 (.A1(n29278), .A2(N10441), .ZN(N47614));
    NOR2X1 U34743 (.A1(N12382), .A2(n24269), .ZN(N47615));
    NOR2X1 U34744 (.A1(n42190), .A2(n39300), .ZN(N47616));
    INVX1 U34745 (.I(N8375), .ZN(N47617));
    NANDX1 U34746 (.A1(n40651), .A2(n19480), .ZN(N47618));
    NANDX1 U34747 (.A1(n33484), .A2(N1470), .ZN(N47619));
    NOR2X1 U34748 (.A1(n16384), .A2(N9901), .ZN(N47620));
    NOR2X1 U34749 (.A1(n19507), .A2(n13898), .ZN(n47621));
    INVX1 U34750 (.I(n23733), .ZN(N47622));
    NANDX1 U34751 (.A1(n34721), .A2(n27747), .ZN(N47623));
    NOR2X1 U34752 (.A1(N2269), .A2(n15271), .ZN(N47624));
    NANDX1 U34753 (.A1(n31547), .A2(n25712), .ZN(N47625));
    NANDX1 U34754 (.A1(n33608), .A2(n39660), .ZN(N47626));
    NANDX1 U34755 (.A1(n22005), .A2(n35487), .ZN(N47627));
    NANDX1 U34756 (.A1(n30379), .A2(N6743), .ZN(N47628));
    NANDX1 U34757 (.A1(n39538), .A2(N8760), .ZN(n47629));
    NANDX1 U34758 (.A1(n41007), .A2(n39264), .ZN(N47630));
    NOR2X1 U34759 (.A1(n40588), .A2(n41137), .ZN(N47631));
    INVX1 U34760 (.I(N693), .ZN(N47632));
    INVX1 U34761 (.I(N5789), .ZN(N47633));
    NANDX1 U34762 (.A1(n21087), .A2(n33535), .ZN(N47634));
    NANDX1 U34763 (.A1(n13036), .A2(n38485), .ZN(n47635));
    INVX1 U34764 (.I(n34262), .ZN(N47636));
    NANDX1 U34765 (.A1(n38822), .A2(n24397), .ZN(n47637));
    INVX1 U34766 (.I(n15829), .ZN(n47638));
    INVX1 U34767 (.I(n31758), .ZN(N47639));
    INVX1 U34768 (.I(n22988), .ZN(n47640));
    NOR2X1 U34769 (.A1(N5392), .A2(n19053), .ZN(N47641));
    NOR2X1 U34770 (.A1(N5351), .A2(N6268), .ZN(N47642));
    NOR2X1 U34771 (.A1(n21693), .A2(N3383), .ZN(N47643));
    NOR2X1 U34772 (.A1(N3749), .A2(n37227), .ZN(N47644));
    NANDX1 U34773 (.A1(n42689), .A2(N4101), .ZN(n47645));
    NOR2X1 U34774 (.A1(n22431), .A2(n42626), .ZN(N47646));
    NANDX1 U34775 (.A1(n17443), .A2(n32436), .ZN(N47647));
    INVX1 U34776 (.I(n27847), .ZN(N47648));
    NANDX1 U34777 (.A1(n24788), .A2(n24118), .ZN(N47649));
    INVX1 U34778 (.I(n27717), .ZN(N47650));
    NANDX1 U34779 (.A1(n18417), .A2(N7232), .ZN(N47651));
    INVX1 U34780 (.I(n23809), .ZN(N47652));
    INVX1 U34781 (.I(n34051), .ZN(N47653));
    NOR2X1 U34782 (.A1(n32551), .A2(n23309), .ZN(N47654));
    INVX1 U34783 (.I(n25613), .ZN(N47655));
    NANDX1 U34784 (.A1(N807), .A2(N9047), .ZN(N47656));
    NOR2X1 U34785 (.A1(N23), .A2(n13147), .ZN(N47657));
    NOR2X1 U34786 (.A1(n22453), .A2(N12300), .ZN(N47658));
    NANDX1 U34787 (.A1(n29575), .A2(n34415), .ZN(N47659));
    NOR2X1 U34788 (.A1(N3629), .A2(N8407), .ZN(N47660));
    INVX1 U34789 (.I(n27746), .ZN(n47661));
    NOR2X1 U34790 (.A1(n21946), .A2(n40149), .ZN(N47662));
    NANDX1 U34791 (.A1(n18857), .A2(n37259), .ZN(n47663));
    INVX1 U34792 (.I(n34820), .ZN(N47664));
    NOR2X1 U34793 (.A1(N5498), .A2(n13579), .ZN(N47665));
    INVX1 U34794 (.I(N2556), .ZN(N47666));
    NOR2X1 U34795 (.A1(n40737), .A2(n36514), .ZN(N47667));
    NANDX1 U34796 (.A1(n26449), .A2(n26216), .ZN(N47668));
    NOR2X1 U34797 (.A1(N8728), .A2(n38348), .ZN(n47669));
    NANDX1 U34798 (.A1(n21250), .A2(n24450), .ZN(N47670));
    NANDX1 U34799 (.A1(n34164), .A2(n28079), .ZN(N47671));
    INVX1 U34800 (.I(n18073), .ZN(N47672));
    NOR2X1 U34801 (.A1(n29979), .A2(n40018), .ZN(n47673));
    INVX1 U34802 (.I(n36302), .ZN(N47674));
    NOR2X1 U34803 (.A1(n35967), .A2(N12641), .ZN(N47675));
    NANDX1 U34804 (.A1(n20331), .A2(N7818), .ZN(N47676));
    INVX1 U34805 (.I(n17684), .ZN(N47677));
    NANDX1 U34806 (.A1(n38878), .A2(N4628), .ZN(N47678));
    NANDX1 U34807 (.A1(n33323), .A2(n20756), .ZN(N47679));
    NANDX1 U34808 (.A1(n40914), .A2(n29484), .ZN(N47680));
    NOR2X1 U34809 (.A1(n40165), .A2(N7261), .ZN(N47681));
    NANDX1 U34810 (.A1(n40679), .A2(n31104), .ZN(N47682));
    INVX1 U34811 (.I(n39279), .ZN(N47683));
    NOR2X1 U34812 (.A1(n14951), .A2(n25785), .ZN(N47684));
    INVX1 U34813 (.I(N3339), .ZN(N47685));
    INVX1 U34814 (.I(n40482), .ZN(N47686));
    INVX1 U34815 (.I(N10615), .ZN(N47687));
    NANDX1 U34816 (.A1(n16163), .A2(n18433), .ZN(N47688));
    NOR2X1 U34817 (.A1(n23527), .A2(N8165), .ZN(N47689));
    INVX1 U34818 (.I(n28154), .ZN(N47690));
    NOR2X1 U34819 (.A1(N11532), .A2(N5438), .ZN(N47691));
    NANDX1 U34820 (.A1(n42126), .A2(n24601), .ZN(N47692));
    NOR2X1 U34821 (.A1(n38818), .A2(n31861), .ZN(N47693));
    INVX1 U34822 (.I(n25704), .ZN(N47694));
    NANDX1 U34823 (.A1(N1551), .A2(n21510), .ZN(N47695));
    NANDX1 U34824 (.A1(N6181), .A2(n36975), .ZN(N47696));
    NOR2X1 U34825 (.A1(N9519), .A2(n34949), .ZN(N47697));
    NOR2X1 U34826 (.A1(n38503), .A2(N2091), .ZN(N47698));
    NANDX1 U34827 (.A1(N11194), .A2(N10203), .ZN(N47699));
    NANDX1 U34828 (.A1(n24400), .A2(n18368), .ZN(N47700));
    NOR2X1 U34829 (.A1(N9081), .A2(N9306), .ZN(N47701));
    NANDX1 U34830 (.A1(N4198), .A2(n19552), .ZN(N47702));
    NANDX1 U34831 (.A1(n28798), .A2(n23342), .ZN(N47703));
    NOR2X1 U34832 (.A1(N6867), .A2(n22293), .ZN(N47704));
    INVX1 U34833 (.I(n16039), .ZN(N47705));
    NANDX1 U34834 (.A1(N2881), .A2(N10274), .ZN(N47706));
    INVX1 U34835 (.I(n29535), .ZN(N47707));
    INVX1 U34836 (.I(n18902), .ZN(N47708));
    NANDX1 U34837 (.A1(n23084), .A2(n13933), .ZN(N47709));
    NOR2X1 U34838 (.A1(n32847), .A2(n14806), .ZN(N47710));
    NANDX1 U34839 (.A1(n25415), .A2(n39205), .ZN(N47711));
    INVX1 U34840 (.I(n39665), .ZN(N47712));
    INVX1 U34841 (.I(n30016), .ZN(N47713));
    INVX1 U34842 (.I(n42163), .ZN(N47714));
    NOR2X1 U34843 (.A1(n36088), .A2(n27488), .ZN(n47715));
    NOR2X1 U34844 (.A1(N2075), .A2(n34354), .ZN(N47716));
    NANDX1 U34845 (.A1(n26918), .A2(n40072), .ZN(n47717));
    NOR2X1 U34846 (.A1(n19479), .A2(N6874), .ZN(N47718));
    NOR2X1 U34847 (.A1(N5541), .A2(N3311), .ZN(N47719));
    NOR2X1 U34848 (.A1(n16232), .A2(n16074), .ZN(N47720));
    NANDX1 U34849 (.A1(n29013), .A2(n38601), .ZN(N47721));
    NOR2X1 U34850 (.A1(n41676), .A2(n20543), .ZN(N47722));
    NANDX1 U34851 (.A1(n18915), .A2(N6415), .ZN(N47723));
    NANDX1 U34852 (.A1(n38610), .A2(n18068), .ZN(N47724));
    NOR2X1 U34853 (.A1(n34385), .A2(N363), .ZN(N47725));
    NANDX1 U34854 (.A1(n43182), .A2(n35590), .ZN(N47726));
    NOR2X1 U34855 (.A1(n30799), .A2(n19035), .ZN(n47727));
    NOR2X1 U34856 (.A1(n21618), .A2(n38513), .ZN(N47728));
    INVX1 U34857 (.I(n21821), .ZN(N47729));
    INVX1 U34858 (.I(n33140), .ZN(N47730));
    NOR2X1 U34859 (.A1(N6493), .A2(n38894), .ZN(N47731));
    INVX1 U34860 (.I(n25185), .ZN(N47732));
    NANDX1 U34861 (.A1(n26730), .A2(n13068), .ZN(N47733));
    NANDX1 U34862 (.A1(n39343), .A2(n21662), .ZN(N47734));
    NANDX1 U34863 (.A1(n36128), .A2(n16800), .ZN(N47735));
    NOR2X1 U34864 (.A1(n31604), .A2(n40864), .ZN(N47736));
    INVX1 U34865 (.I(N775), .ZN(N47737));
    NOR2X1 U34866 (.A1(N7414), .A2(n37451), .ZN(N47738));
    NANDX1 U34867 (.A1(n16128), .A2(n16935), .ZN(N47739));
    NANDX1 U34868 (.A1(N849), .A2(N3292), .ZN(n47740));
    INVX1 U34869 (.I(n34582), .ZN(N47741));
    NANDX1 U34870 (.A1(n37829), .A2(n30754), .ZN(N47742));
    NANDX1 U34871 (.A1(n37357), .A2(N12466), .ZN(N47743));
    NOR2X1 U34872 (.A1(n20614), .A2(n25533), .ZN(N47744));
    NANDX1 U34873 (.A1(N6164), .A2(n36875), .ZN(N47745));
    INVX1 U34874 (.I(n42291), .ZN(N47746));
    NANDX1 U34875 (.A1(n14333), .A2(n20102), .ZN(N47747));
    NANDX1 U34876 (.A1(n19309), .A2(N10556), .ZN(N47748));
    NOR2X1 U34877 (.A1(n26722), .A2(N4535), .ZN(N47749));
    INVX1 U34878 (.I(n32529), .ZN(N47750));
    INVX1 U34879 (.I(n20188), .ZN(N47751));
    NOR2X1 U34880 (.A1(N4121), .A2(n27412), .ZN(n47752));
    INVX1 U34881 (.I(n30232), .ZN(N47753));
    NANDX1 U34882 (.A1(N1447), .A2(n41444), .ZN(N47754));
    NOR2X1 U34883 (.A1(n13912), .A2(n43205), .ZN(N47755));
    NOR2X1 U34884 (.A1(n29125), .A2(N2265), .ZN(N47756));
    NANDX1 U34885 (.A1(n22527), .A2(N1664), .ZN(N47757));
    NOR2X1 U34886 (.A1(n22408), .A2(N5676), .ZN(n47758));
    NOR2X1 U34887 (.A1(N9360), .A2(n24984), .ZN(N47759));
    NOR2X1 U34888 (.A1(n36885), .A2(N8233), .ZN(N47760));
    NANDX1 U34889 (.A1(n28197), .A2(n30441), .ZN(N47761));
    NOR2X1 U34890 (.A1(N4912), .A2(n20346), .ZN(N47762));
    NOR2X1 U34891 (.A1(n32324), .A2(n24191), .ZN(N47763));
    INVX1 U34892 (.I(N299), .ZN(N47764));
    NOR2X1 U34893 (.A1(n24836), .A2(N5631), .ZN(N47765));
    NOR2X1 U34894 (.A1(n24568), .A2(n21255), .ZN(N47766));
    INVX1 U34895 (.I(n16513), .ZN(N47767));
    NOR2X1 U34896 (.A1(n27087), .A2(n18176), .ZN(N47768));
    NANDX1 U34897 (.A1(n39174), .A2(n23851), .ZN(N47769));
    NANDX1 U34898 (.A1(N5062), .A2(n38514), .ZN(N47770));
    INVX1 U34899 (.I(n31626), .ZN(n47771));
    NOR2X1 U34900 (.A1(N6568), .A2(n16350), .ZN(N47772));
    NANDX1 U34901 (.A1(N9402), .A2(n21262), .ZN(N47773));
    NANDX1 U34902 (.A1(n16355), .A2(n43265), .ZN(N47774));
    NOR2X1 U34903 (.A1(n43220), .A2(n33243), .ZN(N47775));
    NANDX1 U34904 (.A1(n14263), .A2(n28553), .ZN(N47776));
    NANDX1 U34905 (.A1(n38831), .A2(N6336), .ZN(N47777));
    NOR2X1 U34906 (.A1(N1551), .A2(n39058), .ZN(N47778));
    NOR2X1 U34907 (.A1(N9406), .A2(n15762), .ZN(N47779));
    NANDX1 U34908 (.A1(n22936), .A2(N12533), .ZN(N47780));
    NANDX1 U34909 (.A1(n17977), .A2(n27416), .ZN(N47781));
    INVX1 U34910 (.I(N10930), .ZN(N47782));
    INVX1 U34911 (.I(n21164), .ZN(N47783));
    NANDX1 U34912 (.A1(n22744), .A2(n42425), .ZN(N47784));
    NANDX1 U34913 (.A1(n39099), .A2(n31897), .ZN(N47785));
    INVX1 U34914 (.I(n28526), .ZN(N47786));
    NOR2X1 U34915 (.A1(n14069), .A2(n42788), .ZN(N47787));
    INVX1 U34916 (.I(n29279), .ZN(N47788));
    NANDX1 U34917 (.A1(n35915), .A2(N5578), .ZN(N47789));
    NANDX1 U34918 (.A1(n31500), .A2(n31796), .ZN(N47790));
    INVX1 U34919 (.I(n36941), .ZN(N47791));
    NOR2X1 U34920 (.A1(N7924), .A2(N6001), .ZN(N47792));
    INVX1 U34921 (.I(n25900), .ZN(N47793));
    INVX1 U34922 (.I(n42036), .ZN(N47794));
    NANDX1 U34923 (.A1(N3287), .A2(n19727), .ZN(N47795));
    NANDX1 U34924 (.A1(n15710), .A2(N8359), .ZN(N47796));
    NOR2X1 U34925 (.A1(N11336), .A2(n40255), .ZN(N47797));
    NOR2X1 U34926 (.A1(n29541), .A2(N8130), .ZN(N47798));
    NANDX1 U34927 (.A1(n18537), .A2(N4557), .ZN(N47799));
    NOR2X1 U34928 (.A1(N2890), .A2(n30151), .ZN(N47800));
    INVX1 U34929 (.I(n21946), .ZN(N47801));
    NOR2X1 U34930 (.A1(n22210), .A2(n40086), .ZN(N47802));
    INVX1 U34931 (.I(n32452), .ZN(N47803));
    NOR2X1 U34932 (.A1(N7326), .A2(n26202), .ZN(N47804));
    INVX1 U34933 (.I(n30422), .ZN(N47805));
    INVX1 U34934 (.I(N3154), .ZN(N47806));
    NOR2X1 U34935 (.A1(n34172), .A2(N10193), .ZN(N47807));
    NANDX1 U34936 (.A1(n42530), .A2(n20861), .ZN(N47808));
    NANDX1 U34937 (.A1(n39313), .A2(n26463), .ZN(n47809));
    NANDX1 U34938 (.A1(n37122), .A2(n35813), .ZN(N47810));
    NANDX1 U34939 (.A1(n41678), .A2(n30969), .ZN(N47811));
    NANDX1 U34940 (.A1(n28356), .A2(n21383), .ZN(N47812));
    INVX1 U34941 (.I(n36213), .ZN(N47813));
    INVX1 U34942 (.I(n35205), .ZN(N47814));
    NANDX1 U34943 (.A1(n32571), .A2(n29422), .ZN(N47815));
    INVX1 U34944 (.I(N4980), .ZN(N47816));
    INVX1 U34945 (.I(n21492), .ZN(N47817));
    NANDX1 U34946 (.A1(n42372), .A2(n34559), .ZN(N47818));
    INVX1 U34947 (.I(n42244), .ZN(N47819));
    NANDX1 U34948 (.A1(N9181), .A2(n19632), .ZN(N47820));
    INVX1 U34949 (.I(n38173), .ZN(N47821));
    INVX1 U34950 (.I(n22044), .ZN(N47822));
    NOR2X1 U34951 (.A1(n28114), .A2(N2649), .ZN(N47823));
    NANDX1 U34952 (.A1(N5290), .A2(n19295), .ZN(N47824));
    INVX1 U34953 (.I(n26673), .ZN(N47825));
    INVX1 U34954 (.I(n30482), .ZN(N47826));
    NOR2X1 U34955 (.A1(N6146), .A2(n24547), .ZN(N47827));
    INVX1 U34956 (.I(n35568), .ZN(N47828));
    NANDX1 U34957 (.A1(n33382), .A2(n31314), .ZN(N47829));
    INVX1 U34958 (.I(N9334), .ZN(N47830));
    INVX1 U34959 (.I(N7556), .ZN(N47831));
    NOR2X1 U34960 (.A1(n28984), .A2(n27419), .ZN(N47832));
    NANDX1 U34961 (.A1(N5143), .A2(n33602), .ZN(N47833));
    NANDX1 U34962 (.A1(n40916), .A2(N1853), .ZN(N47834));
    NOR2X1 U34963 (.A1(n15237), .A2(n37653), .ZN(N47835));
    INVX1 U34964 (.I(n20526), .ZN(N47836));
    NOR2X1 U34965 (.A1(n38176), .A2(N3726), .ZN(N47837));
    NOR2X1 U34966 (.A1(n25185), .A2(N9878), .ZN(n47838));
    INVX1 U34967 (.I(n39412), .ZN(N47839));
    NOR2X1 U34968 (.A1(N5489), .A2(N1237), .ZN(N47840));
    NOR2X1 U34969 (.A1(n36802), .A2(n28025), .ZN(N47841));
    NOR2X1 U34970 (.A1(n13222), .A2(n35580), .ZN(N47842));
    NANDX1 U34971 (.A1(n42205), .A2(N9206), .ZN(N47843));
    NOR2X1 U34972 (.A1(n37027), .A2(n32487), .ZN(n47844));
    NOR2X1 U34973 (.A1(n24150), .A2(n34340), .ZN(N47845));
    NANDX1 U34974 (.A1(n39386), .A2(n18200), .ZN(N47846));
    NANDX1 U34975 (.A1(n16439), .A2(n31675), .ZN(N47847));
    INVX1 U34976 (.I(N9845), .ZN(N47848));
    INVX1 U34977 (.I(n27442), .ZN(N47849));
    NOR2X1 U34978 (.A1(n29483), .A2(n13061), .ZN(N47850));
    NOR2X1 U34979 (.A1(n34971), .A2(n14297), .ZN(N47851));
    NOR2X1 U34980 (.A1(n17980), .A2(n42321), .ZN(N47852));
    NANDX1 U34981 (.A1(n31201), .A2(n24109), .ZN(N47853));
    NANDX1 U34982 (.A1(n19613), .A2(n33314), .ZN(N47854));
    NANDX1 U34983 (.A1(n13167), .A2(N12009), .ZN(N47855));
    INVX1 U34984 (.I(n26996), .ZN(N47856));
    INVX1 U34985 (.I(n18346), .ZN(N47857));
    INVX1 U34986 (.I(N10755), .ZN(N47858));
    NANDX1 U34987 (.A1(n29028), .A2(n42429), .ZN(N47859));
    NOR2X1 U34988 (.A1(n38872), .A2(N4727), .ZN(N47860));
    INVX1 U34989 (.I(N4801), .ZN(N47861));
    INVX1 U34990 (.I(n35505), .ZN(N47862));
    NANDX1 U34991 (.A1(n15388), .A2(N6329), .ZN(N47863));
    NANDX1 U34992 (.A1(n23047), .A2(n38330), .ZN(N47864));
    NANDX1 U34993 (.A1(N10776), .A2(N8646), .ZN(N47865));
    NOR2X1 U34994 (.A1(n30388), .A2(n31639), .ZN(N47866));
    INVX1 U34995 (.I(n33235), .ZN(N47867));
    NOR2X1 U34996 (.A1(n31623), .A2(N6438), .ZN(N47868));
    NOR2X1 U34997 (.A1(n39648), .A2(n29347), .ZN(N47869));
    NANDX1 U34998 (.A1(n32395), .A2(n14902), .ZN(N47870));
    NANDX1 U34999 (.A1(n27399), .A2(n43453), .ZN(N47871));
    NOR2X1 U35000 (.A1(n39523), .A2(N4781), .ZN(N47872));
    INVX1 U35001 (.I(n21236), .ZN(n47873));
    INVX1 U35002 (.I(n25803), .ZN(N47874));
    NOR2X1 U35003 (.A1(n22041), .A2(N5377), .ZN(N47875));
    NANDX1 U35004 (.A1(n13268), .A2(N5832), .ZN(N47876));
    INVX1 U35005 (.I(n23808), .ZN(N47877));
    NOR2X1 U35006 (.A1(n42065), .A2(n21373), .ZN(N47878));
    NANDX1 U35007 (.A1(n31919), .A2(N9523), .ZN(n47879));
    INVX1 U35008 (.I(n24649), .ZN(N47880));
    NANDX1 U35009 (.A1(n41125), .A2(n17813), .ZN(N47881));
    NOR2X1 U35010 (.A1(N2234), .A2(N9933), .ZN(N47882));
    NOR2X1 U35011 (.A1(N2214), .A2(n39932), .ZN(N47883));
    INVX1 U35012 (.I(n40146), .ZN(N47884));
    NANDX1 U35013 (.A1(N8344), .A2(N10462), .ZN(N47885));
    NANDX1 U35014 (.A1(n25588), .A2(n32503), .ZN(N47886));
    NANDX1 U35015 (.A1(n27368), .A2(n35450), .ZN(N47887));
    NOR2X1 U35016 (.A1(n37794), .A2(n15786), .ZN(N47888));
    NANDX1 U35017 (.A1(n26066), .A2(n26838), .ZN(N47889));
    NOR2X1 U35018 (.A1(n14512), .A2(n36360), .ZN(N47890));
    INVX1 U35019 (.I(n28840), .ZN(N47891));
    NANDX1 U35020 (.A1(n20444), .A2(N3180), .ZN(N47892));
    NANDX1 U35021 (.A1(N12357), .A2(n13113), .ZN(N47893));
    INVX1 U35022 (.I(N4251), .ZN(N47894));
    NANDX1 U35023 (.A1(n37676), .A2(N924), .ZN(N47895));
    NOR2X1 U35024 (.A1(n35699), .A2(N1066), .ZN(N47896));
    NANDX1 U35025 (.A1(n17814), .A2(n23248), .ZN(N47897));
    INVX1 U35026 (.I(n34862), .ZN(N47898));
    NOR2X1 U35027 (.A1(N2834), .A2(n29183), .ZN(N47899));
    INVX1 U35028 (.I(N8505), .ZN(N47900));
    INVX1 U35029 (.I(N4055), .ZN(N47901));
    NANDX1 U35030 (.A1(n15967), .A2(n40414), .ZN(n47902));
    NOR2X1 U35031 (.A1(N1335), .A2(n18359), .ZN(N47903));
    NANDX1 U35032 (.A1(N4514), .A2(n24075), .ZN(N47904));
    NANDX1 U35033 (.A1(N7306), .A2(n20850), .ZN(N47905));
    NOR2X1 U35034 (.A1(N6557), .A2(N4733), .ZN(N47906));
    NOR2X1 U35035 (.A1(N12682), .A2(n40431), .ZN(N47907));
    INVX1 U35036 (.I(N8011), .ZN(N47908));
    INVX1 U35037 (.I(n19841), .ZN(N47909));
    INVX1 U35038 (.I(n39314), .ZN(N47910));
    NANDX1 U35039 (.A1(N2946), .A2(n14704), .ZN(N47911));
    NOR2X1 U35040 (.A1(N11451), .A2(n16159), .ZN(N47912));
    NOR2X1 U35041 (.A1(n20647), .A2(n32125), .ZN(N47913));
    NOR2X1 U35042 (.A1(N9162), .A2(n23139), .ZN(N47914));
    INVX1 U35043 (.I(N7800), .ZN(N47915));
    NOR2X1 U35044 (.A1(n24751), .A2(N8475), .ZN(N47916));
    NANDX1 U35045 (.A1(N2128), .A2(n13399), .ZN(N47917));
    NOR2X1 U35046 (.A1(n40012), .A2(N8927), .ZN(N47918));
    NOR2X1 U35047 (.A1(n36971), .A2(N5520), .ZN(N47919));
    NOR2X1 U35048 (.A1(n41423), .A2(n15040), .ZN(N47920));
    NOR2X1 U35049 (.A1(n26944), .A2(n39785), .ZN(n47921));
    NOR2X1 U35050 (.A1(n41647), .A2(n41747), .ZN(N47922));
    NOR2X1 U35051 (.A1(n14333), .A2(N4291), .ZN(N47923));
    NOR2X1 U35052 (.A1(n36137), .A2(n40401), .ZN(n47924));
    NANDX1 U35053 (.A1(N5484), .A2(n41077), .ZN(N47925));
    INVX1 U35054 (.I(n22816), .ZN(N47926));
    NANDX1 U35055 (.A1(n17404), .A2(n37133), .ZN(N47927));
    INVX1 U35056 (.I(n30802), .ZN(N47928));
    NOR2X1 U35057 (.A1(N10703), .A2(n29409), .ZN(N47929));
    NOR2X1 U35058 (.A1(N4201), .A2(n24608), .ZN(N47930));
    NOR2X1 U35059 (.A1(n35303), .A2(n39648), .ZN(N47931));
    NOR2X1 U35060 (.A1(n18774), .A2(n35960), .ZN(N47932));
    NANDX1 U35061 (.A1(N6628), .A2(n34234), .ZN(N47933));
    NOR2X1 U35062 (.A1(N10640), .A2(n28204), .ZN(N47934));
    NOR2X1 U35063 (.A1(N3304), .A2(n25133), .ZN(N47935));
    INVX1 U35064 (.I(n41939), .ZN(N47936));
    INVX1 U35065 (.I(n18890), .ZN(N47937));
    NANDX1 U35066 (.A1(N1620), .A2(n25973), .ZN(N47938));
    NOR2X1 U35067 (.A1(n15783), .A2(N2983), .ZN(N47939));
    NANDX1 U35068 (.A1(n16165), .A2(n32391), .ZN(N47940));
    NANDX1 U35069 (.A1(n20365), .A2(n13526), .ZN(N47941));
    INVX1 U35070 (.I(N1875), .ZN(N47942));
    INVX1 U35071 (.I(n33981), .ZN(N47943));
    NOR2X1 U35072 (.A1(n25020), .A2(n27923), .ZN(N47944));
    NOR2X1 U35073 (.A1(N5461), .A2(n24146), .ZN(N47945));
    NOR2X1 U35074 (.A1(n33665), .A2(N12337), .ZN(N47946));
    NOR2X1 U35075 (.A1(n15325), .A2(n22297), .ZN(n47947));
    NOR2X1 U35076 (.A1(n27741), .A2(n30867), .ZN(N47948));
    NANDX1 U35077 (.A1(n19041), .A2(n13367), .ZN(N47949));
    INVX1 U35078 (.I(n24503), .ZN(N47950));
    NANDX1 U35079 (.A1(N12504), .A2(n40667), .ZN(N47951));
    INVX1 U35080 (.I(n28150), .ZN(N47952));
    NANDX1 U35081 (.A1(n41625), .A2(n25869), .ZN(N47953));
    NANDX1 U35082 (.A1(n41005), .A2(N6057), .ZN(N47954));
    INVX1 U35083 (.I(N12233), .ZN(N47955));
    INVX1 U35084 (.I(n26074), .ZN(n47956));
    NANDX1 U35085 (.A1(N4332), .A2(n43347), .ZN(N47957));
    NANDX1 U35086 (.A1(n16668), .A2(n20451), .ZN(N47958));
    NOR2X1 U35087 (.A1(n38965), .A2(n29174), .ZN(N47959));
    NANDX1 U35088 (.A1(n16039), .A2(N5387), .ZN(N47960));
    INVX1 U35089 (.I(n29405), .ZN(N47961));
    NOR2X1 U35090 (.A1(n30380), .A2(n35434), .ZN(N47962));
    NANDX1 U35091 (.A1(n27574), .A2(n30380), .ZN(N47963));
    INVX1 U35092 (.I(n34812), .ZN(N47964));
    NANDX1 U35093 (.A1(n21782), .A2(N452), .ZN(N47965));
    NANDX1 U35094 (.A1(n17518), .A2(N9571), .ZN(N47966));
    NANDX1 U35095 (.A1(N8025), .A2(n35644), .ZN(N47967));
    NOR2X1 U35096 (.A1(N12356), .A2(n35518), .ZN(N47968));
    NOR2X1 U35097 (.A1(n29024), .A2(N2176), .ZN(N47969));
    NANDX1 U35098 (.A1(n14196), .A2(n21030), .ZN(N47970));
    INVX1 U35099 (.I(n30234), .ZN(N47971));
    INVX1 U35100 (.I(n38516), .ZN(N47972));
    NANDX1 U35101 (.A1(n25148), .A2(n25423), .ZN(N47973));
    NANDX1 U35102 (.A1(n36384), .A2(n42676), .ZN(N47974));
    INVX1 U35103 (.I(n32297), .ZN(N47975));
    NOR2X1 U35104 (.A1(n36078), .A2(N286), .ZN(N47976));
    NOR2X1 U35105 (.A1(n41502), .A2(n17803), .ZN(N47977));
    NOR2X1 U35106 (.A1(n15686), .A2(n25827), .ZN(N47978));
    INVX1 U35107 (.I(N7563), .ZN(N47979));
    NOR2X1 U35108 (.A1(n40764), .A2(n40476), .ZN(N47980));
    NANDX1 U35109 (.A1(n32620), .A2(n32485), .ZN(N47981));
    NANDX1 U35110 (.A1(N10177), .A2(n21652), .ZN(N47982));
    NANDX1 U35111 (.A1(n26272), .A2(N6375), .ZN(N47983));
    NOR2X1 U35112 (.A1(n41099), .A2(n31798), .ZN(N47984));
    NOR2X1 U35113 (.A1(n23690), .A2(n31001), .ZN(N47985));
    NOR2X1 U35114 (.A1(N12514), .A2(N11224), .ZN(N47986));
    NANDX1 U35115 (.A1(N12799), .A2(n25049), .ZN(N47987));
    NANDX1 U35116 (.A1(n20282), .A2(n15293), .ZN(N47988));
    INVX1 U35117 (.I(n35788), .ZN(N47989));
    NANDX1 U35118 (.A1(N8490), .A2(n20178), .ZN(N47990));
    INVX1 U35119 (.I(n38645), .ZN(N47991));
    INVX1 U35120 (.I(n40130), .ZN(N47992));
    INVX1 U35121 (.I(n40559), .ZN(N47993));
    NOR2X1 U35122 (.A1(n38989), .A2(N1136), .ZN(N47994));
    NANDX1 U35123 (.A1(N1891), .A2(N711), .ZN(N47995));
    INVX1 U35124 (.I(n23368), .ZN(N47996));
    INVX1 U35125 (.I(n33781), .ZN(N47997));
    NANDX1 U35126 (.A1(N3019), .A2(N2822), .ZN(N47998));
    NANDX1 U35127 (.A1(N551), .A2(N5301), .ZN(N47999));
    NANDX1 U35128 (.A1(n39585), .A2(n25582), .ZN(N48000));
    NOR2X1 U35129 (.A1(N7361), .A2(N7577), .ZN(N48001));
    NOR2X1 U35130 (.A1(n15850), .A2(n27755), .ZN(N48002));
    INVX1 U35131 (.I(N703), .ZN(N48003));
    INVX1 U35132 (.I(N12734), .ZN(N48004));
    NANDX1 U35133 (.A1(N4640), .A2(N9247), .ZN(N48005));
    NANDX1 U35134 (.A1(n38927), .A2(n32031), .ZN(N48006));
    NOR2X1 U35135 (.A1(n29317), .A2(n42121), .ZN(N48007));
    NANDX1 U35136 (.A1(n17088), .A2(n22109), .ZN(N48008));
    NOR2X1 U35137 (.A1(N9786), .A2(n24931), .ZN(N48009));
    NANDX1 U35138 (.A1(N10337), .A2(n19911), .ZN(N48010));
    INVX1 U35139 (.I(n39601), .ZN(N48011));
    NANDX1 U35140 (.A1(N1632), .A2(n36641), .ZN(N48012));
    NOR2X1 U35141 (.A1(N10198), .A2(n42171), .ZN(N48013));
    INVX1 U35142 (.I(n15954), .ZN(N48014));
    INVX1 U35143 (.I(n24263), .ZN(N48015));
    NOR2X1 U35144 (.A1(n27760), .A2(n18582), .ZN(N48016));
    INVX1 U35145 (.I(n30995), .ZN(N48017));
    NANDX1 U35146 (.A1(n16171), .A2(N2968), .ZN(N48018));
    NOR2X1 U35147 (.A1(N4499), .A2(n21141), .ZN(N48019));
    INVX1 U35148 (.I(n26608), .ZN(N48020));
    INVX1 U35149 (.I(N6114), .ZN(N48021));
    NANDX1 U35150 (.A1(n26966), .A2(N6130), .ZN(N48022));
    INVX1 U35151 (.I(n40570), .ZN(N48023));
    INVX1 U35152 (.I(n42507), .ZN(N48024));
    NANDX1 U35153 (.A1(n38899), .A2(n41782), .ZN(N48025));
    NOR2X1 U35154 (.A1(n37597), .A2(n15020), .ZN(N48026));
    INVX1 U35155 (.I(n36997), .ZN(N48027));
    NANDX1 U35156 (.A1(n32925), .A2(N10964), .ZN(n48028));
    INVX1 U35157 (.I(n17065), .ZN(N48029));
    NOR2X1 U35158 (.A1(n40938), .A2(n22915), .ZN(N48030));
    NOR2X1 U35159 (.A1(n20178), .A2(n27413), .ZN(N48031));
    NANDX1 U35160 (.A1(N6186), .A2(N10548), .ZN(N48032));
    NOR2X1 U35161 (.A1(N12299), .A2(N8293), .ZN(N48033));
    NOR2X1 U35162 (.A1(n18428), .A2(n15628), .ZN(N48034));
    NOR2X1 U35163 (.A1(N10365), .A2(n14662), .ZN(N48035));
    NANDX1 U35164 (.A1(n38943), .A2(N2652), .ZN(N48036));
    INVX1 U35165 (.I(n33067), .ZN(N48037));
    INVX1 U35166 (.I(n24005), .ZN(N48038));
    INVX1 U35167 (.I(n36312), .ZN(n48039));
    NOR2X1 U35168 (.A1(n16914), .A2(n30062), .ZN(N48040));
    NANDX1 U35169 (.A1(n15399), .A2(n17207), .ZN(N48041));
    INVX1 U35170 (.I(n39684), .ZN(N48042));
    NOR2X1 U35171 (.A1(n16735), .A2(N8485), .ZN(N48043));
    NOR2X1 U35172 (.A1(n16963), .A2(n17175), .ZN(N48044));
    NANDX1 U35173 (.A1(n14935), .A2(N9359), .ZN(N48045));
    NANDX1 U35174 (.A1(n30563), .A2(n31792), .ZN(N48046));
    NOR2X1 U35175 (.A1(N1752), .A2(N9481), .ZN(N48047));
    NOR2X1 U35176 (.A1(n37555), .A2(n18927), .ZN(n48048));
    NOR2X1 U35177 (.A1(N1433), .A2(n32611), .ZN(N48049));
    INVX1 U35178 (.I(n37744), .ZN(N48050));
    INVX1 U35179 (.I(n18156), .ZN(N48051));
    NANDX1 U35180 (.A1(n35307), .A2(n23235), .ZN(N48052));
    NOR2X1 U35181 (.A1(n14309), .A2(n19446), .ZN(N48053));
    NOR2X1 U35182 (.A1(n31044), .A2(n17610), .ZN(N48054));
    NOR2X1 U35183 (.A1(n37686), .A2(n24464), .ZN(N48055));
    NANDX1 U35184 (.A1(N9148), .A2(n23503), .ZN(N48056));
    NOR2X1 U35185 (.A1(n39710), .A2(N11822), .ZN(n48057));
    NOR2X1 U35186 (.A1(n31142), .A2(N10983), .ZN(N48058));
    NANDX1 U35187 (.A1(n25224), .A2(n29909), .ZN(N48059));
    NANDX1 U35188 (.A1(n16337), .A2(N8728), .ZN(n48060));
    NOR2X1 U35189 (.A1(N288), .A2(n34154), .ZN(N48061));
    INVX1 U35190 (.I(n14301), .ZN(N48062));
    INVX1 U35191 (.I(n19092), .ZN(N48063));
    INVX1 U35192 (.I(n29977), .ZN(N48064));
    INVX1 U35193 (.I(n39691), .ZN(N48065));
    NOR2X1 U35194 (.A1(n35506), .A2(n33959), .ZN(N48066));
    NOR2X1 U35195 (.A1(n16498), .A2(n30302), .ZN(N48067));
    NANDX1 U35196 (.A1(n40000), .A2(n26507), .ZN(N48068));
    INVX1 U35197 (.I(n41501), .ZN(N48069));
    INVX1 U35198 (.I(n17327), .ZN(N48070));
    NANDX1 U35199 (.A1(N1595), .A2(n32231), .ZN(N48071));
    NANDX1 U35200 (.A1(n31847), .A2(N5095), .ZN(N48072));
    NANDX1 U35201 (.A1(n19869), .A2(N5382), .ZN(N48073));
    NOR2X1 U35202 (.A1(N5406), .A2(N9362), .ZN(N48074));
    NOR2X1 U35203 (.A1(n14178), .A2(n34241), .ZN(N48075));
    NOR2X1 U35204 (.A1(n42394), .A2(n20139), .ZN(N48076));
    NOR2X1 U35205 (.A1(n24108), .A2(N10625), .ZN(N48077));
    NOR2X1 U35206 (.A1(n30285), .A2(n30606), .ZN(N48078));
    NANDX1 U35207 (.A1(n26812), .A2(n13640), .ZN(N48079));
    NOR2X1 U35208 (.A1(n14520), .A2(n36258), .ZN(N48080));
    NANDX1 U35209 (.A1(n23531), .A2(n27532), .ZN(N48081));
    NOR2X1 U35210 (.A1(N8658), .A2(n15906), .ZN(N48082));
    NANDX1 U35211 (.A1(n35664), .A2(n25454), .ZN(N48083));
    NOR2X1 U35212 (.A1(N9879), .A2(n30859), .ZN(N48084));
    NOR2X1 U35213 (.A1(n43235), .A2(N1564), .ZN(N48085));
    NANDX1 U35214 (.A1(N9303), .A2(n33638), .ZN(n48086));
    NOR2X1 U35215 (.A1(n15750), .A2(n14273), .ZN(N48087));
    INVX1 U35216 (.I(n33958), .ZN(N48088));
    INVX1 U35217 (.I(N8289), .ZN(N48089));
    NOR2X1 U35218 (.A1(n17576), .A2(N11608), .ZN(N48090));
    NOR2X1 U35219 (.A1(n32095), .A2(N4393), .ZN(N48091));
    INVX1 U35220 (.I(N1833), .ZN(N48092));
    NOR2X1 U35221 (.A1(n25718), .A2(N10490), .ZN(N48093));
    INVX1 U35222 (.I(n31238), .ZN(N48094));
    NANDX1 U35223 (.A1(n19490), .A2(n42139), .ZN(N48095));
    NANDX1 U35224 (.A1(n40029), .A2(n41762), .ZN(N48096));
    NOR2X1 U35225 (.A1(n41592), .A2(n42474), .ZN(N48097));
    NANDX1 U35226 (.A1(n21437), .A2(N9532), .ZN(N48098));
    NOR2X1 U35227 (.A1(n25389), .A2(n30686), .ZN(N48099));
    NANDX1 U35228 (.A1(n26473), .A2(n28654), .ZN(N48100));
    NANDX1 U35229 (.A1(n33728), .A2(n40262), .ZN(n48101));
    INVX1 U35230 (.I(N12031), .ZN(N48102));
    INVX1 U35231 (.I(N3494), .ZN(N48103));
    NOR2X1 U35232 (.A1(n22786), .A2(n29211), .ZN(N48104));
    NOR2X1 U35233 (.A1(n16822), .A2(N6656), .ZN(N48105));
    NANDX1 U35234 (.A1(n25992), .A2(N5323), .ZN(N48106));
    NOR2X1 U35235 (.A1(N12228), .A2(N3612), .ZN(N48107));
    NOR2X1 U35236 (.A1(N27), .A2(n35765), .ZN(N48108));
    NANDX1 U35237 (.A1(n21464), .A2(n34976), .ZN(N48109));
    NOR2X1 U35238 (.A1(N3380), .A2(n22190), .ZN(N48110));
    INVX1 U35239 (.I(n19533), .ZN(N48111));
    NOR2X1 U35240 (.A1(n33298), .A2(N9788), .ZN(n48112));
    NOR2X1 U35241 (.A1(N11501), .A2(n21818), .ZN(N48113));
    NANDX1 U35242 (.A1(N4674), .A2(n25361), .ZN(n48114));
    INVX1 U35243 (.I(n23565), .ZN(N48115));
    NOR2X1 U35244 (.A1(n13988), .A2(n30220), .ZN(N48116));
    INVX1 U35245 (.I(n39979), .ZN(N48117));
    NANDX1 U35246 (.A1(n21265), .A2(n41886), .ZN(N48118));
    NANDX1 U35247 (.A1(n21577), .A2(n41913), .ZN(N48119));
    INVX1 U35248 (.I(N12553), .ZN(N48120));
    INVX1 U35249 (.I(N2310), .ZN(N48121));
    INVX1 U35250 (.I(n12963), .ZN(N48122));
    INVX1 U35251 (.I(n24867), .ZN(N48123));
    NANDX1 U35252 (.A1(N11229), .A2(N4372), .ZN(N48124));
    NANDX1 U35253 (.A1(N5069), .A2(N5552), .ZN(N48125));
    INVX1 U35254 (.I(N90), .ZN(N48126));
    INVX1 U35255 (.I(n25348), .ZN(N48127));
    NOR2X1 U35256 (.A1(n33790), .A2(n21268), .ZN(n48128));
    NANDX1 U35257 (.A1(n20537), .A2(n23581), .ZN(N48129));
    INVX1 U35258 (.I(N2287), .ZN(N48130));
    NOR2X1 U35259 (.A1(n39315), .A2(n20800), .ZN(N48131));
    INVX1 U35260 (.I(n37755), .ZN(N48132));
    INVX1 U35261 (.I(n14861), .ZN(N48133));
    NOR2X1 U35262 (.A1(n13274), .A2(n35121), .ZN(n48134));
    NOR2X1 U35263 (.A1(n27452), .A2(n16515), .ZN(N48135));
    NANDX1 U35264 (.A1(n38681), .A2(N10567), .ZN(n48136));
    INVX1 U35265 (.I(N277), .ZN(N48137));
    INVX1 U35266 (.I(N6841), .ZN(N48138));
    NANDX1 U35267 (.A1(n26343), .A2(n32188), .ZN(N48139));
    NANDX1 U35268 (.A1(N6340), .A2(n43136), .ZN(N48140));
    INVX1 U35269 (.I(n26877), .ZN(N48141));
    NANDX1 U35270 (.A1(N6292), .A2(n18843), .ZN(N48142));
    NANDX1 U35271 (.A1(N2135), .A2(n29322), .ZN(N48143));
    NOR2X1 U35272 (.A1(n29569), .A2(n40286), .ZN(n48144));
    NOR2X1 U35273 (.A1(n33435), .A2(N10088), .ZN(N48145));
    NANDX1 U35274 (.A1(n39943), .A2(n37539), .ZN(n48146));
    NOR2X1 U35275 (.A1(n25153), .A2(n22427), .ZN(N48147));
    NOR2X1 U35276 (.A1(n32006), .A2(n22703), .ZN(N48148));
    INVX1 U35277 (.I(n38846), .ZN(N48149));
    INVX1 U35278 (.I(N7902), .ZN(N48150));
    NOR2X1 U35279 (.A1(n33200), .A2(n14241), .ZN(n48151));
    INVX1 U35280 (.I(n31743), .ZN(N48152));
    INVX1 U35281 (.I(n29827), .ZN(N48153));
    INVX1 U35282 (.I(n39319), .ZN(N48154));
    INVX1 U35283 (.I(n19528), .ZN(N48155));
    NOR2X1 U35284 (.A1(n40086), .A2(N5625), .ZN(N48156));
    NANDX1 U35285 (.A1(n17758), .A2(n28739), .ZN(N48157));
    NANDX1 U35286 (.A1(n30550), .A2(n25209), .ZN(N48158));
    NANDX1 U35287 (.A1(N6065), .A2(n40041), .ZN(N48159));
    NOR2X1 U35288 (.A1(n25298), .A2(n28574), .ZN(N48160));
    NANDX1 U35289 (.A1(n17177), .A2(n13627), .ZN(N48161));
    NOR2X1 U35290 (.A1(n25078), .A2(n30868), .ZN(N48162));
    INVX1 U35291 (.I(n28998), .ZN(n48163));
    INVX1 U35292 (.I(N10409), .ZN(N48164));
    INVX1 U35293 (.I(n34126), .ZN(N48165));
    NANDX1 U35294 (.A1(N1849), .A2(n24455), .ZN(n48166));
    INVX1 U35295 (.I(n16697), .ZN(N48167));
    INVX1 U35296 (.I(N9482), .ZN(N48168));
    INVX1 U35297 (.I(n38825), .ZN(N48169));
    NOR2X1 U35298 (.A1(N6634), .A2(n25903), .ZN(N48170));
    NANDX1 U35299 (.A1(N12128), .A2(n21647), .ZN(N48171));
    INVX1 U35300 (.I(n40049), .ZN(N48172));
    INVX1 U35301 (.I(n24458), .ZN(N48173));
    NANDX1 U35302 (.A1(N10329), .A2(n38085), .ZN(N48174));
    INVX1 U35303 (.I(n25086), .ZN(N48175));
    NANDX1 U35304 (.A1(N4486), .A2(N10611), .ZN(N48176));
    NANDX1 U35305 (.A1(N4575), .A2(n16613), .ZN(N48177));
    NOR2X1 U35306 (.A1(n42697), .A2(n18462), .ZN(N48178));
    INVX1 U35307 (.I(N3082), .ZN(N48179));
    NOR2X1 U35308 (.A1(N1841), .A2(N12564), .ZN(N48180));
    NOR2X1 U35309 (.A1(n40666), .A2(n40463), .ZN(N48181));
    NANDX1 U35310 (.A1(N12776), .A2(N6627), .ZN(N48182));
    INVX1 U35311 (.I(n24102), .ZN(N48183));
    INVX1 U35312 (.I(n14740), .ZN(N48184));
    INVX1 U35313 (.I(n26968), .ZN(N48185));
    NANDX1 U35314 (.A1(n27582), .A2(n21580), .ZN(n48186));
    NOR2X1 U35315 (.A1(N9195), .A2(n36739), .ZN(N48187));
    INVX1 U35316 (.I(n19806), .ZN(N48188));
    INVX1 U35317 (.I(n22386), .ZN(N48189));
    NOR2X1 U35318 (.A1(n22835), .A2(N11290), .ZN(N48190));
    INVX1 U35319 (.I(n13928), .ZN(N48191));
    NOR2X1 U35320 (.A1(n25924), .A2(N5449), .ZN(N48192));
    NANDX1 U35321 (.A1(N2494), .A2(n35794), .ZN(N48193));
    NOR2X1 U35322 (.A1(N8529), .A2(N5097), .ZN(N48194));
    NOR2X1 U35323 (.A1(n37012), .A2(n18878), .ZN(N48195));
    INVX1 U35324 (.I(N8279), .ZN(N48196));
    INVX1 U35325 (.I(N6237), .ZN(N48197));
    NANDX1 U35326 (.A1(n20241), .A2(n17496), .ZN(N48198));
    INVX1 U35327 (.I(n29436), .ZN(N48199));
    NANDX1 U35328 (.A1(n16603), .A2(N5769), .ZN(N48200));
    NOR2X1 U35329 (.A1(n28669), .A2(n31866), .ZN(N48201));
    NOR2X1 U35330 (.A1(n39958), .A2(n22633), .ZN(N48202));
    NANDX1 U35331 (.A1(N537), .A2(N5084), .ZN(N48203));
    NOR2X1 U35332 (.A1(N6831), .A2(n40730), .ZN(N48204));
    NANDX1 U35333 (.A1(n20436), .A2(N5786), .ZN(N48205));
    NOR2X1 U35334 (.A1(n30346), .A2(n32477), .ZN(N48206));
    NOR2X1 U35335 (.A1(n42767), .A2(n40755), .ZN(N48207));
    INVX1 U35336 (.I(n38683), .ZN(N48208));
    NANDX1 U35337 (.A1(n20459), .A2(N12706), .ZN(n48209));
    NANDX1 U35338 (.A1(N6422), .A2(n13148), .ZN(N48210));
    INVX1 U35339 (.I(N1870), .ZN(N48211));
    INVX1 U35340 (.I(n37130), .ZN(N48212));
    NANDX1 U35341 (.A1(n29163), .A2(n23295), .ZN(N48213));
    INVX1 U35342 (.I(n25299), .ZN(N48214));
    INVX1 U35343 (.I(N7659), .ZN(n48215));
    NOR2X1 U35344 (.A1(n20342), .A2(n38068), .ZN(N48216));
    INVX1 U35345 (.I(n40777), .ZN(N48217));
    NOR2X1 U35346 (.A1(N9469), .A2(n17331), .ZN(n48218));
    INVX1 U35347 (.I(n17027), .ZN(N48219));
    INVX1 U35348 (.I(n19820), .ZN(N48220));
    INVX1 U35349 (.I(N11835), .ZN(N48221));
    INVX1 U35350 (.I(n37703), .ZN(N48222));
    INVX1 U35351 (.I(n27578), .ZN(N48223));
    INVX1 U35352 (.I(n27368), .ZN(N48224));
    NOR2X1 U35353 (.A1(n35673), .A2(N10209), .ZN(N48225));
    INVX1 U35354 (.I(n15615), .ZN(N48226));
    NOR2X1 U35355 (.A1(n22031), .A2(n18190), .ZN(N48227));
    NOR2X1 U35356 (.A1(N2390), .A2(n15528), .ZN(N48228));
    NANDX1 U35357 (.A1(n22731), .A2(N10123), .ZN(N48229));
    NOR2X1 U35358 (.A1(N9716), .A2(N183), .ZN(N48230));
    NOR2X1 U35359 (.A1(n16726), .A2(n22720), .ZN(N48231));
    NOR2X1 U35360 (.A1(n33350), .A2(n32220), .ZN(n48232));
    INVX1 U35361 (.I(n34864), .ZN(N48233));
    NOR2X1 U35362 (.A1(n32403), .A2(n38763), .ZN(N48234));
    NANDX1 U35363 (.A1(n22734), .A2(N12338), .ZN(N48235));
    NOR2X1 U35364 (.A1(n14934), .A2(N12227), .ZN(N48236));
    NOR2X1 U35365 (.A1(n30548), .A2(n41277), .ZN(N48237));
    NANDX1 U35366 (.A1(n38417), .A2(N8682), .ZN(N48238));
    NANDX1 U35367 (.A1(N10472), .A2(n36120), .ZN(n48239));
    NANDX1 U35368 (.A1(N10274), .A2(n40874), .ZN(N48240));
    NOR2X1 U35369 (.A1(N10457), .A2(N11623), .ZN(N48241));
    INVX1 U35370 (.I(n22856), .ZN(N48242));
    NOR2X1 U35371 (.A1(N1421), .A2(N11603), .ZN(N48243));
    INVX1 U35372 (.I(n25964), .ZN(N48244));
    NOR2X1 U35373 (.A1(n39013), .A2(N10934), .ZN(N48245));
    NANDX1 U35374 (.A1(n18274), .A2(n23272), .ZN(N48246));
    INVX1 U35375 (.I(n22887), .ZN(n48247));
    INVX1 U35376 (.I(N6564), .ZN(N48248));
    NANDX1 U35377 (.A1(n22982), .A2(n40980), .ZN(N48249));
    INVX1 U35378 (.I(n31663), .ZN(N48250));
    NOR2X1 U35379 (.A1(n38211), .A2(n24311), .ZN(N48251));
    NANDX1 U35380 (.A1(N5012), .A2(N11392), .ZN(N48252));
    INVX1 U35381 (.I(N5148), .ZN(N48253));
    NOR2X1 U35382 (.A1(n36096), .A2(n28004), .ZN(N48254));
    NOR2X1 U35383 (.A1(n27196), .A2(n29286), .ZN(N48255));
    NOR2X1 U35384 (.A1(N9687), .A2(N11563), .ZN(N48256));
    NOR2X1 U35385 (.A1(n20621), .A2(n25243), .ZN(N48257));
    NANDX1 U35386 (.A1(n33572), .A2(N9101), .ZN(N48258));
    NANDX1 U35387 (.A1(n15277), .A2(N5344), .ZN(N48259));
    NOR2X1 U35388 (.A1(n38258), .A2(N2851), .ZN(N48260));
    INVX1 U35389 (.I(n16129), .ZN(n48261));
    INVX1 U35390 (.I(N3090), .ZN(N48262));
    INVX1 U35391 (.I(n35937), .ZN(N48263));
    INVX1 U35392 (.I(n41510), .ZN(N48264));
    INVX1 U35393 (.I(N2929), .ZN(N48265));
    NOR2X1 U35394 (.A1(n42793), .A2(n30932), .ZN(n48266));
    NANDX1 U35395 (.A1(n26517), .A2(N6426), .ZN(N48267));
    NOR2X1 U35396 (.A1(n25883), .A2(N7668), .ZN(N48268));
    NOR2X1 U35397 (.A1(n36183), .A2(n32910), .ZN(N48269));
    NANDX1 U35398 (.A1(n15962), .A2(n31690), .ZN(N48270));
    NOR2X1 U35399 (.A1(n31238), .A2(n37033), .ZN(N48271));
    NOR2X1 U35400 (.A1(n15704), .A2(n29564), .ZN(N48272));
    NANDX1 U35401 (.A1(n31832), .A2(N2614), .ZN(N48273));
    INVX1 U35402 (.I(n18478), .ZN(N48274));
    NOR2X1 U35403 (.A1(n17811), .A2(n16515), .ZN(N48275));
    NOR2X1 U35404 (.A1(n20740), .A2(n27245), .ZN(n48276));
    NOR2X1 U35405 (.A1(n41351), .A2(n29428), .ZN(N48277));
    INVX1 U35406 (.I(n37456), .ZN(N48278));
    INVX1 U35407 (.I(n22534), .ZN(N48279));
    NANDX1 U35408 (.A1(n21329), .A2(N4925), .ZN(N48280));
    NOR2X1 U35409 (.A1(N4221), .A2(n20886), .ZN(N48281));
    NOR2X1 U35410 (.A1(n32197), .A2(N8652), .ZN(N48282));
    INVX1 U35411 (.I(n30465), .ZN(N48283));
    NOR2X1 U35412 (.A1(n35581), .A2(N3933), .ZN(N48284));
    INVX1 U35413 (.I(n27874), .ZN(n48285));
    NANDX1 U35414 (.A1(n20871), .A2(N2311), .ZN(N48286));
    INVX1 U35415 (.I(n37385), .ZN(N48287));
    NOR2X1 U35416 (.A1(n41872), .A2(N10837), .ZN(N48288));
    NANDX1 U35417 (.A1(n29431), .A2(n40264), .ZN(N48289));
    NOR2X1 U35418 (.A1(n23414), .A2(n26464), .ZN(N48290));
    NANDX1 U35419 (.A1(n25065), .A2(n37472), .ZN(N48291));
    NANDX1 U35420 (.A1(N5832), .A2(n41693), .ZN(N48292));
    INVX1 U35421 (.I(n18289), .ZN(N48293));
    NOR2X1 U35422 (.A1(n30058), .A2(n13986), .ZN(N48294));
    INVX1 U35423 (.I(N620), .ZN(N48295));
    INVX1 U35424 (.I(N702), .ZN(N48296));
    NOR2X1 U35425 (.A1(n23647), .A2(N4024), .ZN(N48297));
    INVX1 U35426 (.I(n25957), .ZN(N48298));
    INVX1 U35427 (.I(N7475), .ZN(N48299));
    NOR2X1 U35428 (.A1(n13236), .A2(n18311), .ZN(N48300));
    NANDX1 U35429 (.A1(n42666), .A2(N4783), .ZN(n48301));
    INVX1 U35430 (.I(N12287), .ZN(N48302));
    INVX1 U35431 (.I(N6074), .ZN(N48303));
    INVX1 U35432 (.I(n25246), .ZN(n48304));
    INVX1 U35433 (.I(n22543), .ZN(n48305));
    NOR2X1 U35434 (.A1(n38320), .A2(n30511), .ZN(N48306));
    NOR2X1 U35435 (.A1(n24905), .A2(N1024), .ZN(N48307));
    INVX1 U35436 (.I(n25524), .ZN(N48308));
    NANDX1 U35437 (.A1(n30711), .A2(n18216), .ZN(N48309));
    INVX1 U35438 (.I(n34734), .ZN(n48310));
    NOR2X1 U35439 (.A1(n36079), .A2(N6098), .ZN(N48311));
    NOR2X1 U35440 (.A1(N2009), .A2(n19333), .ZN(N48312));
    NANDX1 U35441 (.A1(N8462), .A2(N8206), .ZN(N48313));
    INVX1 U35442 (.I(n41771), .ZN(N48314));
    INVX1 U35443 (.I(N6646), .ZN(N48315));
    INVX1 U35444 (.I(n37203), .ZN(N48316));
    INVX1 U35445 (.I(N10965), .ZN(N48317));
    NOR2X1 U35446 (.A1(n34716), .A2(N5813), .ZN(N48318));
    NOR2X1 U35447 (.A1(n24485), .A2(n20397), .ZN(N48319));
    NOR2X1 U35448 (.A1(N11023), .A2(N2449), .ZN(N48320));
    INVX1 U35449 (.I(n31413), .ZN(N48321));
    INVX1 U35450 (.I(N932), .ZN(n48322));
    NOR2X1 U35451 (.A1(N8970), .A2(n37010), .ZN(N48323));
    NOR2X1 U35452 (.A1(N4749), .A2(n39018), .ZN(n48324));
    NOR2X1 U35453 (.A1(n18839), .A2(n37160), .ZN(N48325));
    INVX1 U35454 (.I(n27391), .ZN(N48326));
    NOR2X1 U35455 (.A1(N2368), .A2(n23717), .ZN(N48327));
    INVX1 U35456 (.I(n29250), .ZN(N48328));
    NOR2X1 U35457 (.A1(n40473), .A2(n35202), .ZN(N48329));
    INVX1 U35458 (.I(N2813), .ZN(n48330));
    INVX1 U35459 (.I(N7223), .ZN(N48331));
    INVX1 U35460 (.I(n22205), .ZN(N48332));
    NANDX1 U35461 (.A1(n15338), .A2(N2694), .ZN(N48333));
    NANDX1 U35462 (.A1(n25681), .A2(N3625), .ZN(N48334));
    INVX1 U35463 (.I(n24330), .ZN(N48335));
    NANDX1 U35464 (.A1(n16351), .A2(n29079), .ZN(N48336));
    NOR2X1 U35465 (.A1(N342), .A2(n37597), .ZN(N48337));
    INVX1 U35466 (.I(n36010), .ZN(N48338));
    NOR2X1 U35467 (.A1(N1212), .A2(n28057), .ZN(N48339));
    NANDX1 U35468 (.A1(n30720), .A2(n13835), .ZN(N48340));
    INVX1 U35469 (.I(n17401), .ZN(N48341));
    NANDX1 U35470 (.A1(n29784), .A2(n20213), .ZN(N48342));
    INVX1 U35471 (.I(n26687), .ZN(N48343));
    NOR2X1 U35472 (.A1(n35320), .A2(n34611), .ZN(N48344));
    NOR2X1 U35473 (.A1(n38014), .A2(n20156), .ZN(N48345));
    NANDX1 U35474 (.A1(n31318), .A2(n18055), .ZN(N48346));
    INVX1 U35475 (.I(n18160), .ZN(N48347));
    NANDX1 U35476 (.A1(n19943), .A2(N548), .ZN(n48348));
    NANDX1 U35477 (.A1(n14068), .A2(N9774), .ZN(N48349));
    INVX1 U35478 (.I(n25263), .ZN(N48350));
    NOR2X1 U35479 (.A1(n34700), .A2(n27022), .ZN(N48351));
    NOR2X1 U35480 (.A1(N5062), .A2(n20275), .ZN(N48352));
    NOR2X1 U35481 (.A1(N305), .A2(n39739), .ZN(N48353));
    NOR2X1 U35482 (.A1(n23740), .A2(n22953), .ZN(N48354));
    NOR2X1 U35483 (.A1(n15588), .A2(N3771), .ZN(n48355));
    NOR2X1 U35484 (.A1(N10129), .A2(n23927), .ZN(N48356));
    INVX1 U35485 (.I(n31126), .ZN(N48357));
    INVX1 U35486 (.I(n23185), .ZN(N48358));
    NANDX1 U35487 (.A1(n22594), .A2(n43128), .ZN(N48359));
    NANDX1 U35488 (.A1(N3547), .A2(N3403), .ZN(N48360));
    NANDX1 U35489 (.A1(N10190), .A2(n18345), .ZN(n48361));
    INVX1 U35490 (.I(N1417), .ZN(N48362));
    INVX1 U35491 (.I(n27544), .ZN(N48363));
    NANDX1 U35492 (.A1(N11848), .A2(n22536), .ZN(N48364));
    INVX1 U35493 (.I(N8114), .ZN(N48365));
    NANDX1 U35494 (.A1(n20202), .A2(n20746), .ZN(N48366));
    NANDX1 U35495 (.A1(n35789), .A2(n24517), .ZN(N48367));
    NANDX1 U35496 (.A1(n35597), .A2(n38123), .ZN(N48368));
    NOR2X1 U35497 (.A1(n23250), .A2(n36631), .ZN(N48369));
    INVX1 U35498 (.I(n29063), .ZN(N48370));
    NANDX1 U35499 (.A1(N2144), .A2(n25103), .ZN(N48371));
    NANDX1 U35500 (.A1(n38698), .A2(n20597), .ZN(N48372));
    NANDX1 U35501 (.A1(n13570), .A2(n16755), .ZN(n48373));
    INVX1 U35502 (.I(N5143), .ZN(N48374));
    NOR2X1 U35503 (.A1(n16741), .A2(N6671), .ZN(N48375));
    NANDX1 U35504 (.A1(n13202), .A2(n14784), .ZN(n48376));
    INVX1 U35505 (.I(n33403), .ZN(N48377));
    NOR2X1 U35506 (.A1(n41757), .A2(n15399), .ZN(n48378));
    INVX1 U35507 (.I(n42533), .ZN(N48379));
    NOR2X1 U35508 (.A1(N904), .A2(n21837), .ZN(N48380));
    INVX1 U35509 (.I(n27214), .ZN(n48381));
    NOR2X1 U35510 (.A1(N6043), .A2(n32646), .ZN(N48382));
    NANDX1 U35511 (.A1(n31146), .A2(n41624), .ZN(N48383));
    NOR2X1 U35512 (.A1(n41422), .A2(n17319), .ZN(N48384));
    NOR2X1 U35513 (.A1(n14704), .A2(n37902), .ZN(N48385));
    NANDX1 U35514 (.A1(N5210), .A2(N850), .ZN(N48386));
    INVX1 U35515 (.I(N7931), .ZN(N48387));
    NANDX1 U35516 (.A1(n20580), .A2(n38072), .ZN(N48388));
    NANDX1 U35517 (.A1(N2317), .A2(n36357), .ZN(N48389));
    NANDX1 U35518 (.A1(n41722), .A2(n25097), .ZN(N48390));
    NOR2X1 U35519 (.A1(n42625), .A2(n36614), .ZN(N48391));
    NOR2X1 U35520 (.A1(n16047), .A2(n17467), .ZN(N48392));
    NANDX1 U35521 (.A1(N5220), .A2(n33615), .ZN(N48393));
    NANDX1 U35522 (.A1(N3371), .A2(n34669), .ZN(N48394));
    INVX1 U35523 (.I(n20689), .ZN(N48395));
    NOR2X1 U35524 (.A1(n22763), .A2(N4798), .ZN(N48396));
    INVX1 U35525 (.I(n17652), .ZN(N48397));
    NOR2X1 U35526 (.A1(N10743), .A2(n25582), .ZN(N48398));
    INVX1 U35527 (.I(n31322), .ZN(N48399));
    NANDX1 U35528 (.A1(n36190), .A2(n23319), .ZN(N48400));
    NOR2X1 U35529 (.A1(n34930), .A2(n21568), .ZN(N48401));
    INVX1 U35530 (.I(n41192), .ZN(n48402));
    NANDX1 U35531 (.A1(N10663), .A2(n24434), .ZN(n48403));
    INVX1 U35532 (.I(n17809), .ZN(N48404));
    NOR2X1 U35533 (.A1(n21346), .A2(N7951), .ZN(N48405));
    NOR2X1 U35534 (.A1(n24716), .A2(n32300), .ZN(N48406));
    INVX1 U35535 (.I(n35084), .ZN(N48407));
    INVX1 U35536 (.I(n21496), .ZN(N48408));
    NOR2X1 U35537 (.A1(N12106), .A2(n39147), .ZN(N48409));
    NANDX1 U35538 (.A1(n22848), .A2(N10936), .ZN(N48410));
    NOR2X1 U35539 (.A1(N377), .A2(n20797), .ZN(N48411));
    INVX1 U35540 (.I(n13375), .ZN(N48412));
    NANDX1 U35541 (.A1(n41270), .A2(n24623), .ZN(N48413));
    NANDX1 U35542 (.A1(n38989), .A2(n35023), .ZN(N48414));
    NOR2X1 U35543 (.A1(n19950), .A2(N7677), .ZN(N48415));
    NOR2X1 U35544 (.A1(n33667), .A2(n29022), .ZN(N48416));
    NANDX1 U35545 (.A1(n14022), .A2(N10265), .ZN(N48417));
    NANDX1 U35546 (.A1(N12756), .A2(N1876), .ZN(N48418));
    NANDX1 U35547 (.A1(n23931), .A2(n31436), .ZN(N48419));
    INVX1 U35548 (.I(N9286), .ZN(N48420));
    INVX1 U35549 (.I(n23669), .ZN(N48421));
    NOR2X1 U35550 (.A1(n36792), .A2(n24045), .ZN(N48422));
    INVX1 U35551 (.I(N9980), .ZN(N48423));
    INVX1 U35552 (.I(N10766), .ZN(N48424));
    INVX1 U35553 (.I(N8250), .ZN(N48425));
    NANDX1 U35554 (.A1(n36445), .A2(n43272), .ZN(N48426));
    NOR2X1 U35555 (.A1(N2602), .A2(n40628), .ZN(N48427));
    NANDX1 U35556 (.A1(n25949), .A2(n26177), .ZN(N48428));
    NOR2X1 U35557 (.A1(n39970), .A2(n26121), .ZN(N48429));
    INVX1 U35558 (.I(n42405), .ZN(N48430));
    INVX1 U35559 (.I(n18181), .ZN(N48431));
    INVX1 U35560 (.I(N5639), .ZN(N48432));
    INVX1 U35561 (.I(n32149), .ZN(N48433));
    NOR2X1 U35562 (.A1(n42670), .A2(n42049), .ZN(n48434));
    NOR2X1 U35563 (.A1(n23243), .A2(n39594), .ZN(N48435));
    INVX1 U35564 (.I(n40022), .ZN(N48436));
    NANDX1 U35565 (.A1(N8923), .A2(N4799), .ZN(N48437));
    NOR2X1 U35566 (.A1(N1896), .A2(N4598), .ZN(N48438));
    NANDX1 U35567 (.A1(N4497), .A2(n34905), .ZN(N48439));
    INVX1 U35568 (.I(n30445), .ZN(N48440));
    NANDX1 U35569 (.A1(N11092), .A2(n16623), .ZN(N48441));
    INVX1 U35570 (.I(n19917), .ZN(N48442));
    NANDX1 U35571 (.A1(N7612), .A2(n27777), .ZN(N48443));
    NOR2X1 U35572 (.A1(N2930), .A2(N3307), .ZN(N48444));
    INVX1 U35573 (.I(N11097), .ZN(N48445));
    NOR2X1 U35574 (.A1(N5031), .A2(N2263), .ZN(N48446));
    NANDX1 U35575 (.A1(N1152), .A2(N3409), .ZN(N48447));
    INVX1 U35576 (.I(n30870), .ZN(N48448));
    NANDX1 U35577 (.A1(n16773), .A2(n15150), .ZN(N48449));
    INVX1 U35578 (.I(N11050), .ZN(N48450));
    INVX1 U35579 (.I(N8403), .ZN(N48451));
    NANDX1 U35580 (.A1(n35205), .A2(n28528), .ZN(N48452));
    INVX1 U35581 (.I(n35976), .ZN(n48453));
    NANDX1 U35582 (.A1(n43178), .A2(N2100), .ZN(N48454));
    INVX1 U35583 (.I(N7317), .ZN(N48455));
    NANDX1 U35584 (.A1(n24690), .A2(n43398), .ZN(N48456));
    NANDX1 U35585 (.A1(n31143), .A2(N11022), .ZN(N48457));
    INVX1 U35586 (.I(n36173), .ZN(n48458));
    INVX1 U35587 (.I(n30472), .ZN(N48459));
    NANDX1 U35588 (.A1(n16693), .A2(n32126), .ZN(n48460));
    NOR2X1 U35589 (.A1(n18704), .A2(N5427), .ZN(N48461));
    INVX1 U35590 (.I(n22610), .ZN(N48462));
    INVX1 U35591 (.I(n37459), .ZN(N48463));
    INVX1 U35592 (.I(n41790), .ZN(N48464));
    NANDX1 U35593 (.A1(n38900), .A2(N8087), .ZN(N48465));
    NOR2X1 U35594 (.A1(n30257), .A2(N7793), .ZN(N48466));
    NOR2X1 U35595 (.A1(n26848), .A2(N4789), .ZN(n48467));
    NANDX1 U35596 (.A1(n41217), .A2(N4715), .ZN(N48468));
    NOR2X1 U35597 (.A1(n28888), .A2(N5416), .ZN(N48469));
    INVX1 U35598 (.I(n21588), .ZN(N48470));
    INVX1 U35599 (.I(n37296), .ZN(N48471));
    NANDX1 U35600 (.A1(n14753), .A2(n25950), .ZN(N48472));
    INVX1 U35601 (.I(n33456), .ZN(N48473));
    INVX1 U35602 (.I(n28430), .ZN(N48474));
    NOR2X1 U35603 (.A1(n27211), .A2(N12096), .ZN(N48475));
    NOR2X1 U35604 (.A1(n25528), .A2(n20646), .ZN(N48476));
    NOR2X1 U35605 (.A1(n23295), .A2(n21700), .ZN(N48477));
    NANDX1 U35606 (.A1(n31087), .A2(n24853), .ZN(N48478));
    INVX1 U35607 (.I(n25555), .ZN(N48479));
    NOR2X1 U35608 (.A1(N9129), .A2(n30269), .ZN(N48480));
    NANDX1 U35609 (.A1(n27696), .A2(n25365), .ZN(N48481));
    NOR2X1 U35610 (.A1(n38963), .A2(n33744), .ZN(N48482));
    NANDX1 U35611 (.A1(n33762), .A2(N5024), .ZN(N48483));
    NANDX1 U35612 (.A1(n42962), .A2(n28160), .ZN(N48484));
    NOR2X1 U35613 (.A1(n17599), .A2(n30433), .ZN(N48485));
    INVX1 U35614 (.I(n29695), .ZN(N48486));
    NOR2X1 U35615 (.A1(n42467), .A2(N6868), .ZN(n48487));
    NOR2X1 U35616 (.A1(n22289), .A2(n28567), .ZN(N48488));
    NANDX1 U35617 (.A1(n43055), .A2(n43099), .ZN(N48489));
    NOR2X1 U35618 (.A1(n25137), .A2(n36868), .ZN(N48490));
    INVX1 U35619 (.I(N1614), .ZN(N48491));
    NOR2X1 U35620 (.A1(n30100), .A2(n26978), .ZN(N48492));
    INVX1 U35621 (.I(n25591), .ZN(N48493));
    NOR2X1 U35622 (.A1(N11305), .A2(N5560), .ZN(N48494));
    NANDX1 U35623 (.A1(n33770), .A2(n38201), .ZN(N48495));
    NOR2X1 U35624 (.A1(n23498), .A2(N12328), .ZN(N48496));
    INVX1 U35625 (.I(N7284), .ZN(N48497));
    NOR2X1 U35626 (.A1(N6037), .A2(n39430), .ZN(N48498));
    NANDX1 U35627 (.A1(n24034), .A2(n18246), .ZN(N48499));
    INVX1 U35628 (.I(n16247), .ZN(N48500));
    NOR2X1 U35629 (.A1(N2650), .A2(n19843), .ZN(N48501));
    INVX1 U35630 (.I(n29198), .ZN(N48502));
    NANDX1 U35631 (.A1(n34258), .A2(N8141), .ZN(N48503));
    INVX1 U35632 (.I(n17763), .ZN(N48504));
    INVX1 U35633 (.I(n13825), .ZN(N48505));
    INVX1 U35634 (.I(n23913), .ZN(N48506));
    NOR2X1 U35635 (.A1(n16003), .A2(N3890), .ZN(N48507));
    NANDX1 U35636 (.A1(N2322), .A2(n27387), .ZN(N48508));
    NOR2X1 U35637 (.A1(n41905), .A2(n24351), .ZN(n48509));
    NANDX1 U35638 (.A1(N4469), .A2(n20308), .ZN(n48510));
    NANDX1 U35639 (.A1(n18182), .A2(n38554), .ZN(N48511));
    NANDX1 U35640 (.A1(n34428), .A2(N2589), .ZN(N48512));
    NANDX1 U35641 (.A1(N479), .A2(n35233), .ZN(N48513));
    NOR2X1 U35642 (.A1(N12406), .A2(n26018), .ZN(n48514));
    NANDX1 U35643 (.A1(N640), .A2(n33460), .ZN(N48515));
    NOR2X1 U35644 (.A1(n14465), .A2(N4359), .ZN(N48516));
    NOR2X1 U35645 (.A1(n23529), .A2(n20361), .ZN(N48517));
    NANDX1 U35646 (.A1(n17001), .A2(N12363), .ZN(N48518));
    NANDX1 U35647 (.A1(n22801), .A2(N10795), .ZN(N48519));
    INVX1 U35648 (.I(n16829), .ZN(n48520));
    NOR2X1 U35649 (.A1(n26686), .A2(n28786), .ZN(N48521));
    INVX1 U35650 (.I(N11447), .ZN(n48522));
    INVX1 U35651 (.I(n14081), .ZN(N48523));
    NANDX1 U35652 (.A1(n38564), .A2(N4239), .ZN(N48524));
    NOR2X1 U35653 (.A1(N8766), .A2(n16644), .ZN(N48525));
    INVX1 U35654 (.I(N9941), .ZN(N48526));
    INVX1 U35655 (.I(N11481), .ZN(N48527));
    INVX1 U35656 (.I(n21427), .ZN(N48528));
    NOR2X1 U35657 (.A1(n28269), .A2(N1483), .ZN(N48529));
    INVX1 U35658 (.I(n26382), .ZN(N48530));
    NANDX1 U35659 (.A1(n17602), .A2(N8410), .ZN(N48531));
    INVX1 U35660 (.I(n18076), .ZN(N48532));
    INVX1 U35661 (.I(n37472), .ZN(N48533));
    NANDX1 U35662 (.A1(n31154), .A2(n22786), .ZN(N48534));
    NOR2X1 U35663 (.A1(n42600), .A2(n33399), .ZN(N48535));
    NOR2X1 U35664 (.A1(N2843), .A2(n28490), .ZN(N48536));
    NOR2X1 U35665 (.A1(n41791), .A2(n26936), .ZN(N48537));
    NANDX1 U35666 (.A1(n19812), .A2(n26556), .ZN(N48538));
    NOR2X1 U35667 (.A1(n31292), .A2(N6808), .ZN(N48539));
    NANDX1 U35668 (.A1(n26491), .A2(n35076), .ZN(N48540));
    INVX1 U35669 (.I(n42050), .ZN(N48541));
    NANDX1 U35670 (.A1(N11555), .A2(n16179), .ZN(N48542));
    NANDX1 U35671 (.A1(n32198), .A2(n34254), .ZN(N48543));
    INVX1 U35672 (.I(n26198), .ZN(n48544));
    NOR2X1 U35673 (.A1(N8224), .A2(N5511), .ZN(N48545));
    NANDX1 U35674 (.A1(n40503), .A2(n38909), .ZN(N48546));
    NANDX1 U35675 (.A1(n43346), .A2(n13607), .ZN(N48547));
    INVX1 U35676 (.I(n31344), .ZN(n48548));
    NANDX1 U35677 (.A1(N7092), .A2(N7683), .ZN(N48549));
    INVX1 U35678 (.I(n31046), .ZN(N48550));
    INVX1 U35679 (.I(N9793), .ZN(N48551));
    INVX1 U35680 (.I(N11672), .ZN(N48552));
    NOR2X1 U35681 (.A1(n26027), .A2(N10249), .ZN(N48553));
    INVX1 U35682 (.I(n27261), .ZN(n48554));
    INVX1 U35683 (.I(n14816), .ZN(N48555));
    INVX1 U35684 (.I(N6889), .ZN(n48556));
    INVX1 U35685 (.I(n42184), .ZN(N48557));
    INVX1 U35686 (.I(n33261), .ZN(N48558));
    NANDX1 U35687 (.A1(n26840), .A2(n19971), .ZN(N48559));
    NANDX1 U35688 (.A1(N6270), .A2(N9524), .ZN(N48560));
    NANDX1 U35689 (.A1(n29521), .A2(n40867), .ZN(N48561));
    INVX1 U35690 (.I(n36612), .ZN(N48562));
    INVX1 U35691 (.I(n15510), .ZN(N48563));
    INVX1 U35692 (.I(n23411), .ZN(N48564));
    NANDX1 U35693 (.A1(N3348), .A2(n24762), .ZN(N48565));
    NANDX1 U35694 (.A1(n29374), .A2(n35011), .ZN(N48566));
    INVX1 U35695 (.I(n13162), .ZN(N48567));
    NOR2X1 U35696 (.A1(n29933), .A2(n29148), .ZN(N48568));
    INVX1 U35697 (.I(N11498), .ZN(N48569));
    NANDX1 U35698 (.A1(n14581), .A2(n34438), .ZN(N48570));
    NOR2X1 U35699 (.A1(n31100), .A2(N10936), .ZN(N48571));
    NOR2X1 U35700 (.A1(n37369), .A2(n20460), .ZN(N48572));
    INVX1 U35701 (.I(n13097), .ZN(N48573));
    INVX1 U35702 (.I(N5926), .ZN(N48574));
    NANDX1 U35703 (.A1(N12611), .A2(n21435), .ZN(N48575));
    NOR2X1 U35704 (.A1(n25701), .A2(N3264), .ZN(N48576));
    INVX1 U35705 (.I(N6990), .ZN(n48577));
    NOR2X1 U35706 (.A1(n32181), .A2(n31680), .ZN(N48578));
    NOR2X1 U35707 (.A1(N1870), .A2(n29005), .ZN(N48579));
    INVX1 U35708 (.I(n20698), .ZN(n48580));
    INVX1 U35709 (.I(n22394), .ZN(N48581));
    NOR2X1 U35710 (.A1(n37478), .A2(N3039), .ZN(N48582));
    INVX1 U35711 (.I(n25105), .ZN(N48583));
    NOR2X1 U35712 (.A1(N6981), .A2(N8682), .ZN(N48584));
    INVX1 U35713 (.I(n33533), .ZN(N48585));
    NANDX1 U35714 (.A1(n41967), .A2(n39458), .ZN(N48586));
    NANDX1 U35715 (.A1(N785), .A2(N7100), .ZN(N48587));
    INVX1 U35716 (.I(n26485), .ZN(N48588));
    NANDX1 U35717 (.A1(n19961), .A2(n33475), .ZN(N48589));
    NOR2X1 U35718 (.A1(N8669), .A2(n21682), .ZN(N48590));
    NANDX1 U35719 (.A1(N218), .A2(N7214), .ZN(N48591));
    INVX1 U35720 (.I(n20915), .ZN(N48592));
    NANDX1 U35721 (.A1(n13297), .A2(N5359), .ZN(N48593));
    NANDX1 U35722 (.A1(n16336), .A2(N11562), .ZN(N48594));
    INVX1 U35723 (.I(n30310), .ZN(N48595));
    NANDX1 U35724 (.A1(N4109), .A2(N10951), .ZN(N48596));
    NANDX1 U35725 (.A1(n15567), .A2(n42597), .ZN(N48597));
    NANDX1 U35726 (.A1(n22940), .A2(n33062), .ZN(N48598));
    INVX1 U35727 (.I(n29773), .ZN(n48599));
    NOR2X1 U35728 (.A1(n34562), .A2(N6261), .ZN(N48600));
    NOR2X1 U35729 (.A1(N452), .A2(n14929), .ZN(N48601));
    NOR2X1 U35730 (.A1(N1098), .A2(n15146), .ZN(N48602));
    NOR2X1 U35731 (.A1(n35473), .A2(n25741), .ZN(N48603));
    NANDX1 U35732 (.A1(N5298), .A2(n31099), .ZN(N48604));
    INVX1 U35733 (.I(N11313), .ZN(N48605));
    NANDX1 U35734 (.A1(n43344), .A2(n31302), .ZN(N48606));
    INVX1 U35735 (.I(n37132), .ZN(N48607));
    NOR2X1 U35736 (.A1(N5690), .A2(N9226), .ZN(n48608));
    NOR2X1 U35737 (.A1(n43429), .A2(n21845), .ZN(N48609));
    NANDX1 U35738 (.A1(n34476), .A2(N8145), .ZN(N48610));
    NOR2X1 U35739 (.A1(n25565), .A2(N4085), .ZN(N48611));
    NANDX1 U35740 (.A1(n26016), .A2(n19013), .ZN(N48612));
    NANDX1 U35741 (.A1(n16793), .A2(n23839), .ZN(N48613));
    NANDX1 U35742 (.A1(n41946), .A2(N6107), .ZN(N48614));
    INVX1 U35743 (.I(N3771), .ZN(N48615));
    NANDX1 U35744 (.A1(n28374), .A2(n15083), .ZN(N48616));
    NOR2X1 U35745 (.A1(n28245), .A2(n36064), .ZN(N48617));
    NOR2X1 U35746 (.A1(N11584), .A2(n24523), .ZN(N48618));
    NANDX1 U35747 (.A1(n20810), .A2(N12106), .ZN(N48619));
    INVX1 U35748 (.I(n32334), .ZN(N48620));
    NANDX1 U35749 (.A1(n30129), .A2(n30159), .ZN(N48621));
    INVX1 U35750 (.I(N1901), .ZN(N48622));
    NANDX1 U35751 (.A1(n17190), .A2(n17596), .ZN(N48623));
    INVX1 U35752 (.I(N2989), .ZN(N48624));
    INVX1 U35753 (.I(n23302), .ZN(N48625));
    INVX1 U35754 (.I(n32861), .ZN(N48626));
    NANDX1 U35755 (.A1(n16727), .A2(n26311), .ZN(N48627));
    NOR2X1 U35756 (.A1(N1628), .A2(n31073), .ZN(N48628));
    NOR2X1 U35757 (.A1(n19552), .A2(n23664), .ZN(N48629));
    NOR2X1 U35758 (.A1(n31136), .A2(N4714), .ZN(N48630));
    NANDX1 U35759 (.A1(n41625), .A2(N6500), .ZN(N48631));
    NANDX1 U35760 (.A1(n20166), .A2(n28930), .ZN(N48632));
    NANDX1 U35761 (.A1(N6852), .A2(n23966), .ZN(N48633));
    INVX1 U35762 (.I(n30775), .ZN(N48634));
    NOR2X1 U35763 (.A1(n16078), .A2(n30238), .ZN(N48635));
    NANDX1 U35764 (.A1(n40146), .A2(N10067), .ZN(N48636));
    NANDX1 U35765 (.A1(n19214), .A2(n39474), .ZN(N48637));
    INVX1 U35766 (.I(N2053), .ZN(N48638));
    NOR2X1 U35767 (.A1(n34654), .A2(n22805), .ZN(N48639));
    NANDX1 U35768 (.A1(N414), .A2(n36149), .ZN(n48640));
    NANDX1 U35769 (.A1(n21229), .A2(n30542), .ZN(N48641));
    NOR2X1 U35770 (.A1(n19381), .A2(n37041), .ZN(N48642));
    NANDX1 U35771 (.A1(n39546), .A2(N12178), .ZN(N48643));
    INVX1 U35772 (.I(n36078), .ZN(N48644));
    NOR2X1 U35773 (.A1(n17057), .A2(n23380), .ZN(N48645));
    NOR2X1 U35774 (.A1(n33134), .A2(N10145), .ZN(N48646));
    INVX1 U35775 (.I(n29807), .ZN(N48647));
    NANDX1 U35776 (.A1(n30156), .A2(N5549), .ZN(n48648));
    NANDX1 U35777 (.A1(n19710), .A2(n40753), .ZN(N48649));
    NANDX1 U35778 (.A1(N571), .A2(N9765), .ZN(N48650));
    INVX1 U35779 (.I(N984), .ZN(N48651));
    INVX1 U35780 (.I(N8613), .ZN(N48652));
    NANDX1 U35781 (.A1(n22663), .A2(N37), .ZN(N48653));
    NOR2X1 U35782 (.A1(N5911), .A2(N11708), .ZN(N48654));
    NOR2X1 U35783 (.A1(n18089), .A2(n30282), .ZN(N48655));
    NANDX1 U35784 (.A1(n33591), .A2(N3866), .ZN(N48656));
    NOR2X1 U35785 (.A1(n13624), .A2(n26679), .ZN(N48657));
    NOR2X1 U35786 (.A1(n17160), .A2(n13014), .ZN(N48658));
    NANDX1 U35787 (.A1(N3843), .A2(N8242), .ZN(N48659));
    INVX1 U35788 (.I(n23552), .ZN(N48660));
    NOR2X1 U35789 (.A1(N9534), .A2(n13802), .ZN(N48661));
    NANDX1 U35790 (.A1(n18163), .A2(N4466), .ZN(N48662));
    INVX1 U35791 (.I(n16455), .ZN(N48663));
    NANDX1 U35792 (.A1(N9429), .A2(n16491), .ZN(N48664));
    NOR2X1 U35793 (.A1(n15339), .A2(n17879), .ZN(N48665));
    NANDX1 U35794 (.A1(n23107), .A2(N4688), .ZN(N48666));
    NOR2X1 U35795 (.A1(n13226), .A2(n41705), .ZN(N48667));
    NOR2X1 U35796 (.A1(n26849), .A2(n24911), .ZN(N48668));
    NOR2X1 U35797 (.A1(n33688), .A2(n27604), .ZN(N48669));
    NANDX1 U35798 (.A1(n37530), .A2(n25525), .ZN(N48670));
    NANDX1 U35799 (.A1(N7289), .A2(n20726), .ZN(N48671));
    NOR2X1 U35800 (.A1(N10771), .A2(n25692), .ZN(N48672));
    NANDX1 U35801 (.A1(n15236), .A2(N12458), .ZN(N48673));
    NANDX1 U35802 (.A1(n31592), .A2(n21886), .ZN(N48674));
    NOR2X1 U35803 (.A1(n35748), .A2(n37224), .ZN(N48675));
    NANDX1 U35804 (.A1(N3137), .A2(n16859), .ZN(N48676));
    INVX1 U35805 (.I(n23628), .ZN(N48677));
    INVX1 U35806 (.I(N467), .ZN(n48678));
    INVX1 U35807 (.I(n36292), .ZN(N48679));
    NOR2X1 U35808 (.A1(n22725), .A2(n26508), .ZN(N48680));
    NANDX1 U35809 (.A1(n21365), .A2(N10245), .ZN(N48681));
    NANDX1 U35810 (.A1(n25147), .A2(N7214), .ZN(N48682));
    NOR2X1 U35811 (.A1(n28142), .A2(n17984), .ZN(N48683));
    INVX1 U35812 (.I(n38979), .ZN(N48684));
    NANDX1 U35813 (.A1(n19475), .A2(n22798), .ZN(N48685));
    NANDX1 U35814 (.A1(n31040), .A2(N12788), .ZN(N48686));
    NOR2X1 U35815 (.A1(n14472), .A2(n20655), .ZN(N48687));
    INVX1 U35816 (.I(n31330), .ZN(N48688));
    INVX1 U35817 (.I(n30058), .ZN(N48689));
    NANDX1 U35818 (.A1(n13036), .A2(N9921), .ZN(N48690));
    NANDX1 U35819 (.A1(n28093), .A2(n32646), .ZN(N48691));
    INVX1 U35820 (.I(n16962), .ZN(N48692));
    INVX1 U35821 (.I(n26872), .ZN(N48693));
    NOR2X1 U35822 (.A1(n25365), .A2(n23765), .ZN(N48694));
    NANDX1 U35823 (.A1(n43186), .A2(n41748), .ZN(N48695));
    NOR2X1 U35824 (.A1(n38693), .A2(n31494), .ZN(N48696));
    NANDX1 U35825 (.A1(n18018), .A2(n42511), .ZN(N48697));
    NOR2X1 U35826 (.A1(n30805), .A2(N2332), .ZN(N48698));
    INVX1 U35827 (.I(N7988), .ZN(N48699));
    NANDX1 U35828 (.A1(N8429), .A2(n20557), .ZN(N48700));
    NANDX1 U35829 (.A1(n38881), .A2(n33592), .ZN(N48701));
    NOR2X1 U35830 (.A1(n29000), .A2(N7893), .ZN(N48702));
    INVX1 U35831 (.I(N2155), .ZN(n48703));
    NANDX1 U35832 (.A1(N7170), .A2(n18706), .ZN(N48704));
    INVX1 U35833 (.I(n22214), .ZN(N48705));
    INVX1 U35834 (.I(N4776), .ZN(N48706));
    NOR2X1 U35835 (.A1(n30425), .A2(n14154), .ZN(N48707));
    NANDX1 U35836 (.A1(N8126), .A2(n32687), .ZN(N48708));
    NOR2X1 U35837 (.A1(N7164), .A2(n38787), .ZN(N48709));
    NOR2X1 U35838 (.A1(n42648), .A2(n15886), .ZN(N48710));
    INVX1 U35839 (.I(n41089), .ZN(N48711));
    NANDX1 U35840 (.A1(n30400), .A2(N5475), .ZN(N48712));
    NANDX1 U35841 (.A1(n20520), .A2(n23253), .ZN(N48713));
    NOR2X1 U35842 (.A1(n28412), .A2(n19885), .ZN(N48714));
    NOR2X1 U35843 (.A1(n42945), .A2(n16734), .ZN(N48715));
    INVX1 U35844 (.I(n35040), .ZN(N48716));
    NANDX1 U35845 (.A1(n27297), .A2(n29495), .ZN(n48717));
    INVX1 U35846 (.I(n14249), .ZN(N48718));
    NOR2X1 U35847 (.A1(n13908), .A2(n22374), .ZN(n48719));
    INVX1 U35848 (.I(n38752), .ZN(N48720));
    INVX1 U35849 (.I(N7537), .ZN(N48721));
    NOR2X1 U35850 (.A1(n18393), .A2(n23422), .ZN(N48722));
    NANDX1 U35851 (.A1(N5689), .A2(n27095), .ZN(N48723));
    NOR2X1 U35852 (.A1(N11163), .A2(n36496), .ZN(N48724));
    NOR2X1 U35853 (.A1(n24095), .A2(n21104), .ZN(N48725));
    NANDX1 U35854 (.A1(N507), .A2(N7867), .ZN(N48726));
    NOR2X1 U35855 (.A1(N6920), .A2(n36166), .ZN(N48727));
    INVX1 U35856 (.I(n35546), .ZN(N48728));
    NANDX1 U35857 (.A1(N11771), .A2(n32307), .ZN(N48729));
    INVX1 U35858 (.I(N1627), .ZN(N48730));
    NOR2X1 U35859 (.A1(n13141), .A2(n13849), .ZN(N48731));
    NOR2X1 U35860 (.A1(n32358), .A2(n21385), .ZN(N48732));
    NOR2X1 U35861 (.A1(n40430), .A2(n34486), .ZN(n48733));
    INVX1 U35862 (.I(N2646), .ZN(N48734));
    NOR2X1 U35863 (.A1(n41706), .A2(N3488), .ZN(N48735));
    NANDX1 U35864 (.A1(n35491), .A2(n27582), .ZN(N48736));
    NOR2X1 U35865 (.A1(N3896), .A2(n17769), .ZN(N48737));
    NANDX1 U35866 (.A1(N4924), .A2(n24688), .ZN(N48738));
    NANDX1 U35867 (.A1(n40992), .A2(N6442), .ZN(N48739));
    NOR2X1 U35868 (.A1(N9290), .A2(n38748), .ZN(N48740));
    INVX1 U35869 (.I(N596), .ZN(N48741));
    INVX1 U35870 (.I(n25730), .ZN(N48742));
    INVX1 U35871 (.I(n18869), .ZN(n48743));
    NOR2X1 U35872 (.A1(n25508), .A2(n36856), .ZN(N48744));
    INVX1 U35873 (.I(N6201), .ZN(N48745));
    INVX1 U35874 (.I(n37049), .ZN(N48746));
    NANDX1 U35875 (.A1(n39416), .A2(n40536), .ZN(N48747));
    NOR2X1 U35876 (.A1(n21114), .A2(n14326), .ZN(N48748));
    NOR2X1 U35877 (.A1(n14689), .A2(n32094), .ZN(N48749));
    NOR2X1 U35878 (.A1(n19613), .A2(N2989), .ZN(N48750));
    INVX1 U35879 (.I(n17132), .ZN(N48751));
    NANDX1 U35880 (.A1(n26035), .A2(n16101), .ZN(N48752));
    NOR2X1 U35881 (.A1(n38624), .A2(n16696), .ZN(N48753));
    INVX1 U35882 (.I(N10562), .ZN(N48754));
    NOR2X1 U35883 (.A1(N949), .A2(n14856), .ZN(N48755));
    NANDX1 U35884 (.A1(n37805), .A2(N5788), .ZN(N48756));
    NOR2X1 U35885 (.A1(n35515), .A2(n42836), .ZN(N48757));
    NANDX1 U35886 (.A1(n31458), .A2(n39900), .ZN(N48758));
    INVX1 U35887 (.I(n42251), .ZN(N48759));
    NANDX1 U35888 (.A1(N116), .A2(n13468), .ZN(N48760));
    INVX1 U35889 (.I(n35646), .ZN(n48761));
    INVX1 U35890 (.I(n25194), .ZN(N48762));
    INVX1 U35891 (.I(n39891), .ZN(N48763));
    NOR2X1 U35892 (.A1(N1779), .A2(N2199), .ZN(N48764));
    NOR2X1 U35893 (.A1(n30083), .A2(n18894), .ZN(N48765));
    NANDX1 U35894 (.A1(n40644), .A2(n39712), .ZN(N48766));
    NOR2X1 U35895 (.A1(N1707), .A2(n32245), .ZN(N48767));
    NANDX1 U35896 (.A1(n40646), .A2(n41298), .ZN(N48768));
    INVX1 U35897 (.I(n40010), .ZN(N48769));
    INVX1 U35898 (.I(N9228), .ZN(N48770));
    INVX1 U35899 (.I(n27743), .ZN(N48771));
    NANDX1 U35900 (.A1(n26549), .A2(n17538), .ZN(N48772));
    INVX1 U35901 (.I(n15602), .ZN(N48773));
    NOR2X1 U35902 (.A1(n33913), .A2(n30475), .ZN(N48774));
    INVX1 U35903 (.I(n20011), .ZN(N48775));
    INVX1 U35904 (.I(n20387), .ZN(N48776));
    NANDX1 U35905 (.A1(n29994), .A2(N6997), .ZN(N48777));
    INVX1 U35906 (.I(n41082), .ZN(N48778));
    NOR2X1 U35907 (.A1(n16701), .A2(n42798), .ZN(N48779));
    NANDX1 U35908 (.A1(N5473), .A2(n38847), .ZN(N48780));
    NANDX1 U35909 (.A1(n36450), .A2(n26937), .ZN(N48781));
    INVX1 U35910 (.I(N3523), .ZN(N48782));
    NANDX1 U35911 (.A1(N5061), .A2(n20945), .ZN(N48783));
    INVX1 U35912 (.I(n31609), .ZN(N48784));
    INVX1 U35913 (.I(n34684), .ZN(N48785));
    NOR2X1 U35914 (.A1(n37873), .A2(n14804), .ZN(N48786));
    NOR2X1 U35915 (.A1(n13009), .A2(n24494), .ZN(N48787));
    NANDX1 U35916 (.A1(n33395), .A2(n36382), .ZN(N48788));
    NOR2X1 U35917 (.A1(n40391), .A2(n23691), .ZN(N48789));
    NANDX1 U35918 (.A1(n34238), .A2(n40391), .ZN(N48790));
    NANDX1 U35919 (.A1(n19471), .A2(n35543), .ZN(N48791));
    NOR2X1 U35920 (.A1(N12198), .A2(n28520), .ZN(N48792));
    NOR2X1 U35921 (.A1(n24294), .A2(n21722), .ZN(N48793));
    INVX1 U35922 (.I(n29354), .ZN(N48794));
    NOR2X1 U35923 (.A1(N5586), .A2(N7170), .ZN(N48795));
    INVX1 U35924 (.I(n40269), .ZN(N48796));
    INVX1 U35925 (.I(n21756), .ZN(N48797));
    INVX1 U35926 (.I(N3839), .ZN(N48798));
    NANDX1 U35927 (.A1(n25773), .A2(n28716), .ZN(N48799));
    INVX1 U35928 (.I(n18682), .ZN(N48800));
    NANDX1 U35929 (.A1(N11284), .A2(n42372), .ZN(N48801));
    NOR2X1 U35930 (.A1(n35201), .A2(n28970), .ZN(N48802));
    NANDX1 U35931 (.A1(N11199), .A2(N10720), .ZN(N48803));
    NANDX1 U35932 (.A1(n13077), .A2(n39239), .ZN(N48804));
    NANDX1 U35933 (.A1(n37370), .A2(n17488), .ZN(N48805));
    NANDX1 U35934 (.A1(n23252), .A2(N6361), .ZN(N48806));
    NOR2X1 U35935 (.A1(n20101), .A2(n33715), .ZN(N48807));
    NANDX1 U35936 (.A1(N10368), .A2(N1678), .ZN(N48808));
    NANDX1 U35937 (.A1(n14206), .A2(n26121), .ZN(N48809));
    INVX1 U35938 (.I(n32601), .ZN(N48810));
    INVX1 U35939 (.I(N6259), .ZN(N48811));
    INVX1 U35940 (.I(n41449), .ZN(N48812));
    INVX1 U35941 (.I(n24570), .ZN(N48813));
    INVX1 U35942 (.I(n13487), .ZN(N48814));
    NANDX1 U35943 (.A1(n34056), .A2(n24206), .ZN(N48815));
    NOR2X1 U35944 (.A1(N3660), .A2(n19972), .ZN(n48816));
    NANDX1 U35945 (.A1(n30709), .A2(n27139), .ZN(N48817));
    NOR2X1 U35946 (.A1(N168), .A2(n33499), .ZN(N48818));
    NOR2X1 U35947 (.A1(n20269), .A2(n23741), .ZN(N48819));
    NANDX1 U35948 (.A1(n20316), .A2(n15099), .ZN(N48820));
    INVX1 U35949 (.I(n24201), .ZN(N48821));
    NANDX1 U35950 (.A1(n17358), .A2(n13329), .ZN(N48822));
    INVX1 U35951 (.I(n13296), .ZN(N48823));
    INVX1 U35952 (.I(n25889), .ZN(N48824));
    NOR2X1 U35953 (.A1(n13347), .A2(N5274), .ZN(N48825));
    NOR2X1 U35954 (.A1(n31256), .A2(n29009), .ZN(N48826));
    NOR2X1 U35955 (.A1(n25573), .A2(n22348), .ZN(n48827));
    NOR2X1 U35956 (.A1(N6299), .A2(N9584), .ZN(N48828));
    NOR2X1 U35957 (.A1(n42435), .A2(N9752), .ZN(N48829));
    INVX1 U35958 (.I(N9148), .ZN(N48830));
    INVX1 U35959 (.I(n32268), .ZN(n48831));
    NOR2X1 U35960 (.A1(n40015), .A2(N3894), .ZN(N48832));
    NOR2X1 U35961 (.A1(n20743), .A2(n34792), .ZN(N48833));
    NANDX1 U35962 (.A1(n23751), .A2(n19232), .ZN(n48834));
    NANDX1 U35963 (.A1(N12528), .A2(n34801), .ZN(N48835));
    NOR2X1 U35964 (.A1(n25874), .A2(n29754), .ZN(N48836));
    NANDX1 U35965 (.A1(N3337), .A2(n15290), .ZN(N48837));
    NOR2X1 U35966 (.A1(n18589), .A2(n37637), .ZN(N48838));
    NANDX1 U35967 (.A1(n24888), .A2(N3748), .ZN(N48839));
    NOR2X1 U35968 (.A1(n13530), .A2(N3179), .ZN(N48840));
    NOR2X1 U35969 (.A1(N12357), .A2(n22878), .ZN(N48841));
    NANDX1 U35970 (.A1(n35688), .A2(n19420), .ZN(N48842));
    NANDX1 U35971 (.A1(n35008), .A2(n29842), .ZN(N48843));
    INVX1 U35972 (.I(n41365), .ZN(N48844));
    NOR2X1 U35973 (.A1(n21784), .A2(n17545), .ZN(N48845));
    NANDX1 U35974 (.A1(N2792), .A2(n35010), .ZN(N48846));
    INVX1 U35975 (.I(n32545), .ZN(N48847));
    NANDX1 U35976 (.A1(n31217), .A2(N4362), .ZN(N48848));
    INVX1 U35977 (.I(N6333), .ZN(N48849));
    INVX1 U35978 (.I(n22294), .ZN(N48850));
    INVX1 U35979 (.I(n35426), .ZN(N48851));
    NANDX1 U35980 (.A1(n34429), .A2(n28284), .ZN(N48852));
    NOR2X1 U35981 (.A1(N3314), .A2(N7690), .ZN(N48853));
    INVX1 U35982 (.I(n28681), .ZN(N48854));
    NOR2X1 U35983 (.A1(n23765), .A2(n20216), .ZN(N48855));
    INVX1 U35984 (.I(n15997), .ZN(N48856));
    INVX1 U35985 (.I(n36110), .ZN(N48857));
    NOR2X1 U35986 (.A1(n25333), .A2(N4965), .ZN(N48858));
    NOR2X1 U35987 (.A1(N6550), .A2(n32844), .ZN(N48859));
    INVX1 U35988 (.I(n16531), .ZN(N48860));
    NANDX1 U35989 (.A1(n23686), .A2(n26667), .ZN(N48861));
    INVX1 U35990 (.I(N11891), .ZN(N48862));
    NOR2X1 U35991 (.A1(N4348), .A2(n36996), .ZN(N48863));
    INVX1 U35992 (.I(n38777), .ZN(N48864));
    NOR2X1 U35993 (.A1(n32672), .A2(n31770), .ZN(N48865));
    NANDX1 U35994 (.A1(n34884), .A2(n16978), .ZN(N48866));
    NANDX1 U35995 (.A1(n15176), .A2(n26874), .ZN(N48867));
    NANDX1 U35996 (.A1(n20852), .A2(n34661), .ZN(N48868));
    NOR2X1 U35997 (.A1(N4839), .A2(N6201), .ZN(N48869));
    NANDX1 U35998 (.A1(n35090), .A2(N2431), .ZN(N48870));
    NANDX1 U35999 (.A1(N622), .A2(n18961), .ZN(N48871));
    INVX1 U36000 (.I(n13987), .ZN(N48872));
    NANDX1 U36001 (.A1(n42644), .A2(n15557), .ZN(N48873));
    INVX1 U36002 (.I(N3519), .ZN(N48874));
    NANDX1 U36003 (.A1(n24803), .A2(n31975), .ZN(N48875));
    INVX1 U36004 (.I(n14003), .ZN(N48876));
    NOR2X1 U36005 (.A1(n29424), .A2(N5414), .ZN(N48877));
    INVX1 U36006 (.I(N11596), .ZN(N48878));
    INVX1 U36007 (.I(N11), .ZN(N48879));
    NOR2X1 U36008 (.A1(n20800), .A2(n24351), .ZN(N48880));
    NOR2X1 U36009 (.A1(n25638), .A2(n30552), .ZN(N48881));
    INVX1 U36010 (.I(N6936), .ZN(N48882));
    NOR2X1 U36011 (.A1(n42098), .A2(N7557), .ZN(N48883));
    NANDX1 U36012 (.A1(n14349), .A2(n21543), .ZN(N48884));
    INVX1 U36013 (.I(n13520), .ZN(N48885));
    INVX1 U36014 (.I(n43292), .ZN(N48886));
    NOR2X1 U36015 (.A1(n35859), .A2(n24623), .ZN(N48887));
    NANDX1 U36016 (.A1(N2634), .A2(n28305), .ZN(N48888));
    NANDX1 U36017 (.A1(n21737), .A2(n23398), .ZN(N48889));
    NOR2X1 U36018 (.A1(n33333), .A2(n33666), .ZN(N48890));
    INVX1 U36019 (.I(N9619), .ZN(n48891));
    INVX1 U36020 (.I(N2670), .ZN(N48892));
    INVX1 U36021 (.I(n26310), .ZN(n48893));
    NOR2X1 U36022 (.A1(n33667), .A2(n22925), .ZN(N48894));
    NOR2X1 U36023 (.A1(n21972), .A2(n20161), .ZN(N48895));
    NOR2X1 U36024 (.A1(n26001), .A2(n41703), .ZN(n48896));
    NOR2X1 U36025 (.A1(n39520), .A2(n25010), .ZN(N48897));
    NANDX1 U36026 (.A1(N2766), .A2(N7076), .ZN(N48898));
    NOR2X1 U36027 (.A1(n31139), .A2(n42862), .ZN(N48899));
    NOR2X1 U36028 (.A1(n36311), .A2(n21126), .ZN(N48900));
    NOR2X1 U36029 (.A1(n24940), .A2(N666), .ZN(N48901));
    NOR2X1 U36030 (.A1(n36411), .A2(n43436), .ZN(N48902));
    NOR2X1 U36031 (.A1(n39080), .A2(n40460), .ZN(N48903));
    INVX1 U36032 (.I(N8189), .ZN(N48904));
    INVX1 U36033 (.I(N1074), .ZN(N48905));
    NOR2X1 U36034 (.A1(n31986), .A2(n21234), .ZN(N48906));
    NANDX1 U36035 (.A1(n14514), .A2(N9145), .ZN(N48907));
    NOR2X1 U36036 (.A1(N10561), .A2(n23834), .ZN(n48908));
    NANDX1 U36037 (.A1(N3007), .A2(n30909), .ZN(N48909));
    INVX1 U36038 (.I(n23825), .ZN(N48910));
    NOR2X1 U36039 (.A1(n34354), .A2(n16663), .ZN(N48911));
    INVX1 U36040 (.I(n15968), .ZN(N48912));
    NANDX1 U36041 (.A1(n31449), .A2(n20927), .ZN(N48913));
    INVX1 U36042 (.I(n31413), .ZN(N48914));
    NANDX1 U36043 (.A1(n19827), .A2(n18080), .ZN(N48915));
    NANDX1 U36044 (.A1(n28015), .A2(n38414), .ZN(N48916));
    INVX1 U36045 (.I(n27973), .ZN(N48917));
    NOR2X1 U36046 (.A1(n16693), .A2(n28169), .ZN(N48918));
    NOR2X1 U36047 (.A1(n25837), .A2(n20781), .ZN(N48919));
    NANDX1 U36048 (.A1(N6198), .A2(n26268), .ZN(N48920));
    NOR2X1 U36049 (.A1(n26786), .A2(N5140), .ZN(N48921));
    INVX1 U36050 (.I(N3292), .ZN(N48922));
    NOR2X1 U36051 (.A1(n31380), .A2(n34075), .ZN(N48923));
    NOR2X1 U36052 (.A1(n19189), .A2(n22051), .ZN(N48924));
    INVX1 U36053 (.I(n43408), .ZN(N48925));
    NOR2X1 U36054 (.A1(n28511), .A2(N9443), .ZN(N48926));
    NANDX1 U36055 (.A1(n22897), .A2(n27137), .ZN(N48927));
    INVX1 U36056 (.I(N8035), .ZN(N48928));
    NANDX1 U36057 (.A1(n29298), .A2(n24727), .ZN(N48929));
    NOR2X1 U36058 (.A1(n16945), .A2(n40243), .ZN(N48930));
    NANDX1 U36059 (.A1(N4832), .A2(n36120), .ZN(n48931));
    INVX1 U36060 (.I(n39198), .ZN(N48932));
    NOR2X1 U36061 (.A1(n17561), .A2(N123), .ZN(N48933));
    NANDX1 U36062 (.A1(N3262), .A2(n21183), .ZN(N48934));
    NANDX1 U36063 (.A1(n38081), .A2(n30051), .ZN(N48935));
    INVX1 U36064 (.I(n40035), .ZN(N48936));
    NANDX1 U36065 (.A1(N4088), .A2(n14753), .ZN(N48937));
    INVX1 U36066 (.I(n21838), .ZN(N48938));
    INVX1 U36067 (.I(N12773), .ZN(N48939));
    NOR2X1 U36068 (.A1(n35364), .A2(n14090), .ZN(N48940));
    INVX1 U36069 (.I(n16618), .ZN(N48941));
    NOR2X1 U36070 (.A1(n26978), .A2(N3069), .ZN(n48942));
    INVX1 U36071 (.I(n31809), .ZN(N48943));
    INVX1 U36072 (.I(n19317), .ZN(N48944));
    NOR2X1 U36073 (.A1(N4829), .A2(n36878), .ZN(N48945));
    INVX1 U36074 (.I(n17233), .ZN(N48946));
    INVX1 U36075 (.I(n28199), .ZN(N48947));
    NOR2X1 U36076 (.A1(n34747), .A2(n14777), .ZN(N48948));
    NANDX1 U36077 (.A1(n20989), .A2(n24123), .ZN(N48949));
    NOR2X1 U36078 (.A1(n35742), .A2(N9759), .ZN(N48950));
    NANDX1 U36079 (.A1(n19598), .A2(N12212), .ZN(N48951));
    NANDX1 U36080 (.A1(N11489), .A2(n15981), .ZN(N48952));
    NOR2X1 U36081 (.A1(n17787), .A2(n16083), .ZN(n48953));
    INVX1 U36082 (.I(n20855), .ZN(N48954));
    NANDX1 U36083 (.A1(n25702), .A2(n16570), .ZN(N48955));
    INVX1 U36084 (.I(n32596), .ZN(N48956));
    NOR2X1 U36085 (.A1(n15060), .A2(n39612), .ZN(N48957));
    NANDX1 U36086 (.A1(N11726), .A2(n24338), .ZN(N48958));
    NOR2X1 U36087 (.A1(n36152), .A2(n28794), .ZN(N48959));
    INVX1 U36088 (.I(n13669), .ZN(N48960));
    INVX1 U36089 (.I(N6875), .ZN(N48961));
    INVX1 U36090 (.I(N8883), .ZN(N48962));
    NOR2X1 U36091 (.A1(n15215), .A2(N10774), .ZN(N48963));
    NANDX1 U36092 (.A1(n26704), .A2(n26754), .ZN(N48964));
    INVX1 U36093 (.I(N1018), .ZN(N48965));
    NANDX1 U36094 (.A1(n18618), .A2(n21872), .ZN(N48966));
    NANDX1 U36095 (.A1(n33999), .A2(n38441), .ZN(N48967));
    NANDX1 U36096 (.A1(n23122), .A2(N6047), .ZN(n48968));
    INVX1 U36097 (.I(N8941), .ZN(N48969));
    NOR2X1 U36098 (.A1(N6668), .A2(n33278), .ZN(n48970));
    NANDX1 U36099 (.A1(n32499), .A2(N8280), .ZN(N48971));
    NOR2X1 U36100 (.A1(N2695), .A2(n17724), .ZN(N48972));
    INVX1 U36101 (.I(n41784), .ZN(N48973));
    INVX1 U36102 (.I(n30294), .ZN(N48974));
    INVX1 U36103 (.I(n27060), .ZN(N48975));
    NANDX1 U36104 (.A1(n29910), .A2(N21), .ZN(n48976));
    NOR2X1 U36105 (.A1(n30927), .A2(n32537), .ZN(N48977));
    INVX1 U36106 (.I(n42478), .ZN(N48978));
    NANDX1 U36107 (.A1(n37217), .A2(n27126), .ZN(N48979));
    INVX1 U36108 (.I(N6547), .ZN(N48980));
    NANDX1 U36109 (.A1(n19383), .A2(n15487), .ZN(N48981));
    NANDX1 U36110 (.A1(n15730), .A2(N5293), .ZN(N48982));
    INVX1 U36111 (.I(N4756), .ZN(N48983));
    NANDX1 U36112 (.A1(n29458), .A2(n40603), .ZN(N48984));
    NANDX1 U36113 (.A1(n22938), .A2(n28594), .ZN(N48985));
    NOR2X1 U36114 (.A1(N9759), .A2(n31800), .ZN(N48986));
    NANDX1 U36115 (.A1(N596), .A2(n18237), .ZN(n48987));
    NOR2X1 U36116 (.A1(n38989), .A2(n38843), .ZN(N48988));
    NOR2X1 U36117 (.A1(N9055), .A2(n37848), .ZN(N48989));
    NANDX1 U36118 (.A1(n35951), .A2(n21502), .ZN(N48990));
    NANDX1 U36119 (.A1(n42497), .A2(N882), .ZN(N48991));
    NOR2X1 U36120 (.A1(n14512), .A2(n14619), .ZN(N48992));
    INVX1 U36121 (.I(N9484), .ZN(n48993));
    INVX1 U36122 (.I(N3083), .ZN(N48994));
    NOR2X1 U36123 (.A1(N12495), .A2(N213), .ZN(N48995));
    NANDX1 U36124 (.A1(n35432), .A2(n18487), .ZN(N48996));
    INVX1 U36125 (.I(N1718), .ZN(N48997));
    NOR2X1 U36126 (.A1(n40215), .A2(n35465), .ZN(N48998));
    INVX1 U36127 (.I(n40442), .ZN(N48999));
    INVX1 U36128 (.I(n20421), .ZN(N49000));
    NOR2X1 U36129 (.A1(n29715), .A2(n14797), .ZN(N49001));
    INVX1 U36130 (.I(n22193), .ZN(N49002));
    NANDX1 U36131 (.A1(n16477), .A2(n21218), .ZN(N49003));
    INVX1 U36132 (.I(N9395), .ZN(N49004));
    NANDX1 U36133 (.A1(n41477), .A2(N7722), .ZN(N49005));
    NOR2X1 U36134 (.A1(n24514), .A2(N10804), .ZN(N49006));
    NANDX1 U36135 (.A1(n37008), .A2(N697), .ZN(N49007));
    INVX1 U36136 (.I(n18647), .ZN(N49008));
    NANDX1 U36137 (.A1(n24077), .A2(N10044), .ZN(N49009));
    INVX1 U36138 (.I(n20819), .ZN(n49010));
    NOR2X1 U36139 (.A1(n40726), .A2(N7468), .ZN(N49011));
    INVX1 U36140 (.I(N7355), .ZN(N49012));
    INVX1 U36141 (.I(n42090), .ZN(N49013));
    NANDX1 U36142 (.A1(N5708), .A2(N10490), .ZN(N49014));
    NOR2X1 U36143 (.A1(N11864), .A2(n21387), .ZN(N49015));
    NOR2X1 U36144 (.A1(N10938), .A2(N3323), .ZN(N49016));
    INVX1 U36145 (.I(N8339), .ZN(N49017));
    NOR2X1 U36146 (.A1(n33391), .A2(n19143), .ZN(N49018));
    NANDX1 U36147 (.A1(n16606), .A2(N9519), .ZN(N49019));
    NANDX1 U36148 (.A1(n24932), .A2(n28701), .ZN(N49020));
    INVX1 U36149 (.I(n34975), .ZN(N49021));
    INVX1 U36150 (.I(n19731), .ZN(N49022));
    INVX1 U36151 (.I(n41630), .ZN(N49023));
    INVX1 U36152 (.I(N5913), .ZN(N49024));
    NOR2X1 U36153 (.A1(n33438), .A2(n37682), .ZN(N49025));
    INVX1 U36154 (.I(n39146), .ZN(N49026));
    NOR2X1 U36155 (.A1(N1357), .A2(n40689), .ZN(n49027));
    NANDX1 U36156 (.A1(n22550), .A2(n41307), .ZN(N49028));
    NANDX1 U36157 (.A1(n21107), .A2(N6173), .ZN(n49029));
    NANDX1 U36158 (.A1(N705), .A2(n25315), .ZN(N49030));
    INVX1 U36159 (.I(N6990), .ZN(n49031));
    NOR2X1 U36160 (.A1(N72), .A2(n31921), .ZN(n49032));
    NOR2X1 U36161 (.A1(n42456), .A2(n23423), .ZN(N49033));
    INVX1 U36162 (.I(n18714), .ZN(N49034));
    INVX1 U36163 (.I(N8802), .ZN(N49035));
    NANDX1 U36164 (.A1(N2232), .A2(N3993), .ZN(N49036));
    NOR2X1 U36165 (.A1(n29593), .A2(N11014), .ZN(N49037));
    NANDX1 U36166 (.A1(n23971), .A2(N12370), .ZN(N49038));
    INVX1 U36167 (.I(n29416), .ZN(N49039));
    NOR2X1 U36168 (.A1(n39113), .A2(n38184), .ZN(N49040));
    INVX1 U36169 (.I(N1814), .ZN(N49041));
    NOR2X1 U36170 (.A1(N2937), .A2(n16808), .ZN(N49042));
    NOR2X1 U36171 (.A1(N9926), .A2(N8169), .ZN(N49043));
    NOR2X1 U36172 (.A1(n31526), .A2(N7589), .ZN(N49044));
    NOR2X1 U36173 (.A1(N11476), .A2(n18233), .ZN(N49045));
    NANDX1 U36174 (.A1(N7795), .A2(n16714), .ZN(N49046));
    INVX1 U36175 (.I(n43178), .ZN(n49047));
    NOR2X1 U36176 (.A1(n30132), .A2(n29298), .ZN(N49048));
    NOR2X1 U36177 (.A1(n30722), .A2(n42948), .ZN(N49049));
    NOR2X1 U36178 (.A1(n28529), .A2(n28892), .ZN(N49050));
    NOR2X1 U36179 (.A1(n24169), .A2(n23603), .ZN(N49051));
    NOR2X1 U36180 (.A1(n15662), .A2(n34335), .ZN(N49052));
    NOR2X1 U36181 (.A1(n32470), .A2(n16510), .ZN(N49053));
    NOR2X1 U36182 (.A1(n30318), .A2(n31909), .ZN(N49054));
    NOR2X1 U36183 (.A1(n37906), .A2(n35970), .ZN(N49055));
    NOR2X1 U36184 (.A1(N2347), .A2(n25593), .ZN(N49056));
    NANDX1 U36185 (.A1(N8740), .A2(n30168), .ZN(N49057));
    NANDX1 U36186 (.A1(n19126), .A2(n16827), .ZN(N49058));
    NOR2X1 U36187 (.A1(n40524), .A2(n37229), .ZN(N49059));
    INVX1 U36188 (.I(n30820), .ZN(N49060));
    NOR2X1 U36189 (.A1(N9926), .A2(n35393), .ZN(N49061));
    INVX1 U36190 (.I(n23208), .ZN(N49062));
    INVX1 U36191 (.I(N8323), .ZN(N49063));
    NANDX1 U36192 (.A1(n18788), .A2(n40792), .ZN(N49064));
    INVX1 U36193 (.I(n28135), .ZN(N49065));
    NANDX1 U36194 (.A1(N8695), .A2(n25534), .ZN(N49066));
    NOR2X1 U36195 (.A1(N1193), .A2(n24089), .ZN(n49067));
    INVX1 U36196 (.I(n16465), .ZN(N49068));
    NANDX1 U36197 (.A1(n22836), .A2(n36312), .ZN(N49069));
    NANDX1 U36198 (.A1(n41961), .A2(n42819), .ZN(N49070));
    INVX1 U36199 (.I(n28692), .ZN(N49071));
    NANDX1 U36200 (.A1(N11595), .A2(N5719), .ZN(N49072));
    NANDX1 U36201 (.A1(n21520), .A2(n41112), .ZN(N49073));
    NANDX1 U36202 (.A1(n34407), .A2(N6686), .ZN(N49074));
    INVX1 U36203 (.I(n38156), .ZN(N49075));
    INVX1 U36204 (.I(n36520), .ZN(N49076));
    INVX1 U36205 (.I(n32967), .ZN(N49077));
    INVX1 U36206 (.I(n13317), .ZN(N49078));
    INVX1 U36207 (.I(n22114), .ZN(N49079));
    INVX1 U36208 (.I(n18477), .ZN(N49080));
    NANDX1 U36209 (.A1(N10334), .A2(n38593), .ZN(N49081));
    NANDX1 U36210 (.A1(N3173), .A2(N10971), .ZN(N49082));
    NOR2X1 U36211 (.A1(n35671), .A2(N8380), .ZN(N49083));
    NANDX1 U36212 (.A1(n28773), .A2(n19974), .ZN(N49084));
    INVX1 U36213 (.I(n23519), .ZN(N49085));
    INVX1 U36214 (.I(n15149), .ZN(N49086));
    INVX1 U36215 (.I(N11788), .ZN(N49087));
    NANDX1 U36216 (.A1(n27294), .A2(N6472), .ZN(N49088));
    INVX1 U36217 (.I(N10022), .ZN(n49089));
    NOR2X1 U36218 (.A1(N5841), .A2(n20385), .ZN(N49090));
    NANDX1 U36219 (.A1(N10549), .A2(n32178), .ZN(N49091));
    NOR2X1 U36220 (.A1(n29025), .A2(n14595), .ZN(N49092));
    NOR2X1 U36221 (.A1(n13826), .A2(n42678), .ZN(N49093));
    NANDX1 U36222 (.A1(n24796), .A2(n25778), .ZN(N49094));
    INVX1 U36223 (.I(n22855), .ZN(N49095));
    INVX1 U36224 (.I(n32115), .ZN(n49096));
    INVX1 U36225 (.I(N1286), .ZN(N49097));
    NOR2X1 U36226 (.A1(N9890), .A2(N6115), .ZN(N49098));
    NOR2X1 U36227 (.A1(n21677), .A2(N7308), .ZN(N49099));
    INVX1 U36228 (.I(n17828), .ZN(N49100));
    NOR2X1 U36229 (.A1(N6609), .A2(n28921), .ZN(N49101));
    NANDX1 U36230 (.A1(n26994), .A2(N9859), .ZN(N49102));
    NOR2X1 U36231 (.A1(n15699), .A2(n28137), .ZN(N49103));
    INVX1 U36232 (.I(n19973), .ZN(N49104));
    NANDX1 U36233 (.A1(N8461), .A2(n19179), .ZN(N49105));
    NOR2X1 U36234 (.A1(n22936), .A2(N1484), .ZN(n49106));
    INVX1 U36235 (.I(N2319), .ZN(N49107));
    NANDX1 U36236 (.A1(n16404), .A2(n24507), .ZN(N49108));
    INVX1 U36237 (.I(n28565), .ZN(N49109));
    NANDX1 U36238 (.A1(n15491), .A2(N8179), .ZN(N49110));
    NANDX1 U36239 (.A1(n22799), .A2(N4766), .ZN(N49111));
    INVX1 U36240 (.I(n36132), .ZN(N49112));
    NOR2X1 U36241 (.A1(N5556), .A2(N11834), .ZN(N49113));
    NANDX1 U36242 (.A1(N5094), .A2(n31237), .ZN(N49114));
    NOR2X1 U36243 (.A1(n33230), .A2(n25872), .ZN(N49115));
    NOR2X1 U36244 (.A1(n36185), .A2(n24012), .ZN(n49116));
    INVX1 U36245 (.I(n17132), .ZN(n49117));
    INVX1 U36246 (.I(N9948), .ZN(N49118));
    INVX1 U36247 (.I(n38945), .ZN(N49119));
    INVX1 U36248 (.I(n17823), .ZN(N49120));
    INVX1 U36249 (.I(n37735), .ZN(N49121));
    NANDX1 U36250 (.A1(N582), .A2(N9754), .ZN(n49122));
    INVX1 U36251 (.I(n36014), .ZN(N49123));
    NOR2X1 U36252 (.A1(n28371), .A2(N12649), .ZN(N49124));
    NANDX1 U36253 (.A1(n29425), .A2(N7884), .ZN(N49125));
    NOR2X1 U36254 (.A1(N3680), .A2(n12978), .ZN(N49126));
    NOR2X1 U36255 (.A1(n37105), .A2(n35887), .ZN(N49127));
    INVX1 U36256 (.I(n26391), .ZN(N49128));
    INVX1 U36257 (.I(n23091), .ZN(n49129));
    NOR2X1 U36258 (.A1(N2259), .A2(n16245), .ZN(N49130));
    NANDX1 U36259 (.A1(N3678), .A2(N11718), .ZN(N49131));
    NOR2X1 U36260 (.A1(N11181), .A2(n21376), .ZN(N49132));
    NANDX1 U36261 (.A1(N3775), .A2(N11638), .ZN(N49133));
    NOR2X1 U36262 (.A1(n37700), .A2(N4179), .ZN(n49134));
    NOR2X1 U36263 (.A1(n22598), .A2(N6507), .ZN(N49135));
    INVX1 U36264 (.I(n41702), .ZN(N49136));
    NOR2X1 U36265 (.A1(n14989), .A2(N1909), .ZN(N49137));
    INVX1 U36266 (.I(n41989), .ZN(N49138));
    NOR2X1 U36267 (.A1(n19782), .A2(n30748), .ZN(N49139));
    NANDX1 U36268 (.A1(n38061), .A2(N10366), .ZN(N49140));
    INVX1 U36269 (.I(n29999), .ZN(N49141));
    NANDX1 U36270 (.A1(n27156), .A2(n33676), .ZN(N49142));
    NOR2X1 U36271 (.A1(n36203), .A2(N1384), .ZN(N49143));
    NOR2X1 U36272 (.A1(n39513), .A2(n38311), .ZN(N49144));
    NOR2X1 U36273 (.A1(n31936), .A2(n32538), .ZN(N49145));
    NOR2X1 U36274 (.A1(N3118), .A2(N1343), .ZN(N49146));
    NANDX1 U36275 (.A1(N12023), .A2(n32724), .ZN(N49147));
    NOR2X1 U36276 (.A1(n27011), .A2(n34632), .ZN(N49148));
    INVX1 U36277 (.I(n15208), .ZN(N49149));
    INVX1 U36278 (.I(n38169), .ZN(N49150));
    NOR2X1 U36279 (.A1(n21143), .A2(n32757), .ZN(N49151));
    NOR2X1 U36280 (.A1(n13817), .A2(n19283), .ZN(n49152));
    INVX1 U36281 (.I(n40972), .ZN(N49153));
    NANDX1 U36282 (.A1(N3354), .A2(n33702), .ZN(N49154));
    NANDX1 U36283 (.A1(n32096), .A2(n19423), .ZN(N49155));
    INVX1 U36284 (.I(n29004), .ZN(N49156));
    NOR2X1 U36285 (.A1(N7285), .A2(n30089), .ZN(N49157));
    NOR2X1 U36286 (.A1(n41779), .A2(n27361), .ZN(N49158));
    INVX1 U36287 (.I(n31030), .ZN(N49159));
    INVX1 U36288 (.I(n39716), .ZN(N49160));
    NANDX1 U36289 (.A1(n13937), .A2(N11451), .ZN(N49161));
    INVX1 U36290 (.I(N8634), .ZN(N49162));
    NANDX1 U36291 (.A1(n42543), .A2(n31070), .ZN(N49163));
    NANDX1 U36292 (.A1(n12887), .A2(N6881), .ZN(N49164));
    NANDX1 U36293 (.A1(N66), .A2(n39199), .ZN(N49165));
    NOR2X1 U36294 (.A1(n23448), .A2(n29428), .ZN(N49166));
    NOR2X1 U36295 (.A1(n42870), .A2(N4176), .ZN(N49167));
    INVX1 U36296 (.I(N7283), .ZN(N49168));
    NANDX1 U36297 (.A1(n32556), .A2(N7966), .ZN(N49169));
    NOR2X1 U36298 (.A1(N6124), .A2(n20671), .ZN(N49170));
    NOR2X1 U36299 (.A1(n34825), .A2(n16915), .ZN(N49171));
    NOR2X1 U36300 (.A1(N5289), .A2(n28365), .ZN(N49172));
    INVX1 U36301 (.I(N3602), .ZN(N49173));
    INVX1 U36302 (.I(n19343), .ZN(N49174));
    NOR2X1 U36303 (.A1(N4967), .A2(n21910), .ZN(N49175));
    INVX1 U36304 (.I(n40246), .ZN(N49176));
    INVX1 U36305 (.I(n26958), .ZN(N49177));
    INVX1 U36306 (.I(N1950), .ZN(N49178));
    NOR2X1 U36307 (.A1(N8870), .A2(N1347), .ZN(n49179));
    NOR2X1 U36308 (.A1(N11336), .A2(n41782), .ZN(N49180));
    NANDX1 U36309 (.A1(N419), .A2(n39427), .ZN(N49181));
    NANDX1 U36310 (.A1(N6542), .A2(n16626), .ZN(N49182));
    INVX1 U36311 (.I(n31046), .ZN(N49183));
    NANDX1 U36312 (.A1(n26381), .A2(n36335), .ZN(n49184));
    NANDX1 U36313 (.A1(N3181), .A2(n29616), .ZN(N49185));
    INVX1 U36314 (.I(N12204), .ZN(N49186));
    NOR2X1 U36315 (.A1(n34736), .A2(n34113), .ZN(N49187));
    NOR2X1 U36316 (.A1(n31510), .A2(N2295), .ZN(N49188));
    NANDX1 U36317 (.A1(n23443), .A2(N4245), .ZN(N49189));
    NOR2X1 U36318 (.A1(n21992), .A2(n38743), .ZN(N49190));
    NANDX1 U36319 (.A1(n33328), .A2(n26732), .ZN(N49191));
    INVX1 U36320 (.I(n23426), .ZN(N49192));
    NOR2X1 U36321 (.A1(n16679), .A2(n19648), .ZN(N49193));
    NOR2X1 U36322 (.A1(N716), .A2(N7221), .ZN(n49194));
    NANDX1 U36323 (.A1(n27096), .A2(n33235), .ZN(N49195));
    NOR2X1 U36324 (.A1(n19957), .A2(n19379), .ZN(N49196));
    NOR2X1 U36325 (.A1(n21840), .A2(n40193), .ZN(N49197));
    INVX1 U36326 (.I(N12480), .ZN(N49198));
    INVX1 U36327 (.I(n38432), .ZN(N49199));
    NOR2X1 U36328 (.A1(n20185), .A2(N8082), .ZN(N49200));
    NOR2X1 U36329 (.A1(N4516), .A2(n30074), .ZN(N49201));
    NOR2X1 U36330 (.A1(N5935), .A2(N9609), .ZN(N49202));
    INVX1 U36331 (.I(N4940), .ZN(n49203));
    NANDX1 U36332 (.A1(n32746), .A2(N11299), .ZN(N49204));
    INVX1 U36333 (.I(N7945), .ZN(N49205));
    NOR2X1 U36334 (.A1(n16430), .A2(n39515), .ZN(N49206));
    INVX1 U36335 (.I(n39344), .ZN(N49207));
    NOR2X1 U36336 (.A1(n38425), .A2(n15250), .ZN(N49208));
    NOR2X1 U36337 (.A1(n16792), .A2(N1651), .ZN(N49209));
    NOR2X1 U36338 (.A1(n18951), .A2(n40097), .ZN(N49210));
    INVX1 U36339 (.I(n23405), .ZN(N49211));
    NOR2X1 U36340 (.A1(N7554), .A2(n21782), .ZN(N49212));
    NOR2X1 U36341 (.A1(n37627), .A2(n15430), .ZN(N49213));
    NANDX1 U36342 (.A1(N3763), .A2(n25490), .ZN(N49214));
    NANDX1 U36343 (.A1(n36796), .A2(N4443), .ZN(N49215));
    INVX1 U36344 (.I(n35685), .ZN(N49216));
    NOR2X1 U36345 (.A1(n24549), .A2(n41794), .ZN(N49217));
    NANDX1 U36346 (.A1(N9866), .A2(n37665), .ZN(N49218));
    NANDX1 U36347 (.A1(N4818), .A2(n42595), .ZN(n49219));
    NANDX1 U36348 (.A1(N11290), .A2(N773), .ZN(N49220));
    NANDX1 U36349 (.A1(n30240), .A2(n30549), .ZN(n49221));
    INVX1 U36350 (.I(n43324), .ZN(N49222));
    INVX1 U36351 (.I(n42962), .ZN(N49223));
    NANDX1 U36352 (.A1(N4569), .A2(n37116), .ZN(N49224));
    NOR2X1 U36353 (.A1(n21507), .A2(n30558), .ZN(N49225));
    NANDX1 U36354 (.A1(n22745), .A2(n13561), .ZN(N49226));
    INVX1 U36355 (.I(N2128), .ZN(N49227));
    NOR2X1 U36356 (.A1(n38102), .A2(n26677), .ZN(N49228));
    NOR2X1 U36357 (.A1(n36211), .A2(n26222), .ZN(N49229));
    NANDX1 U36358 (.A1(N5933), .A2(n20719), .ZN(N49230));
    NANDX1 U36359 (.A1(n27037), .A2(n32008), .ZN(N49231));
    INVX1 U36360 (.I(n19501), .ZN(N49232));
    NANDX1 U36361 (.A1(n41241), .A2(N11437), .ZN(N49233));
    INVX1 U36362 (.I(n34805), .ZN(N49234));
    INVX1 U36363 (.I(n19620), .ZN(N49235));
    NOR2X1 U36364 (.A1(n37721), .A2(N2891), .ZN(N49236));
    NANDX1 U36365 (.A1(n24806), .A2(N1330), .ZN(N49237));
    NOR2X1 U36366 (.A1(n38367), .A2(n37364), .ZN(n49238));
    NANDX1 U36367 (.A1(n33819), .A2(n31993), .ZN(N49239));
    NANDX1 U36368 (.A1(n27593), .A2(n14412), .ZN(N49240));
    INVX1 U36369 (.I(N5239), .ZN(N49241));
    INVX1 U36370 (.I(n41463), .ZN(N49242));
    INVX1 U36371 (.I(N3908), .ZN(N49243));
    NANDX1 U36372 (.A1(n36171), .A2(n13088), .ZN(N49244));
    NOR2X1 U36373 (.A1(n33939), .A2(n24525), .ZN(N49245));
    INVX1 U36374 (.I(n14951), .ZN(N49246));
    NANDX1 U36375 (.A1(n35420), .A2(N10852), .ZN(N49247));
    NOR2X1 U36376 (.A1(n38310), .A2(n17940), .ZN(N49248));
    NOR2X1 U36377 (.A1(n29319), .A2(n37451), .ZN(N49249));
    NOR2X1 U36378 (.A1(n23211), .A2(n15618), .ZN(N49250));
    NANDX1 U36379 (.A1(N11731), .A2(n20461), .ZN(N49251));
    NANDX1 U36380 (.A1(n15822), .A2(n41205), .ZN(N49252));
    NANDX1 U36381 (.A1(n36165), .A2(n28876), .ZN(N49253));
    NANDX1 U36382 (.A1(n29752), .A2(N5082), .ZN(N49254));
    INVX1 U36383 (.I(n42840), .ZN(N49255));
    NOR2X1 U36384 (.A1(n39937), .A2(n23892), .ZN(N49256));
    NOR2X1 U36385 (.A1(N11415), .A2(N5549), .ZN(N49257));
    INVX1 U36386 (.I(N11947), .ZN(N49258));
    NOR2X1 U36387 (.A1(n25478), .A2(n19566), .ZN(N49259));
    NOR2X1 U36388 (.A1(N11325), .A2(n13544), .ZN(N49260));
    NOR2X1 U36389 (.A1(n24215), .A2(n29162), .ZN(N49261));
    INVX1 U36390 (.I(n35945), .ZN(N49262));
    NOR2X1 U36391 (.A1(n33252), .A2(n41447), .ZN(N49263));
    INVX1 U36392 (.I(n31394), .ZN(n49264));
    NANDX1 U36393 (.A1(n22438), .A2(N1222), .ZN(N49265));
    NANDX1 U36394 (.A1(n27519), .A2(N7220), .ZN(N49266));
    NANDX1 U36395 (.A1(N6941), .A2(n36836), .ZN(N49267));
    NOR2X1 U36396 (.A1(N2162), .A2(n37931), .ZN(N49268));
    NANDX1 U36397 (.A1(n32803), .A2(N6405), .ZN(N49269));
    NOR2X1 U36398 (.A1(n14808), .A2(n15650), .ZN(N49270));
    NANDX1 U36399 (.A1(n15812), .A2(n29193), .ZN(N49271));
    INVX1 U36400 (.I(n40026), .ZN(N49272));
    INVX1 U36401 (.I(N12517), .ZN(n49273));
    INVX1 U36402 (.I(N10712), .ZN(N49274));
    INVX1 U36403 (.I(n20153), .ZN(N49275));
    NOR2X1 U36404 (.A1(n13050), .A2(N499), .ZN(N49276));
    INVX1 U36405 (.I(N3951), .ZN(N49277));
    NOR2X1 U36406 (.A1(n33589), .A2(N11171), .ZN(n49278));
    INVX1 U36407 (.I(n30209), .ZN(N49279));
    NANDX1 U36408 (.A1(N12138), .A2(n22050), .ZN(N49280));
    NANDX1 U36409 (.A1(n20083), .A2(N11380), .ZN(N49281));
    NANDX1 U36410 (.A1(N9482), .A2(n15868), .ZN(N49282));
    INVX1 U36411 (.I(n14199), .ZN(n49283));
    NANDX1 U36412 (.A1(n29598), .A2(n29839), .ZN(N49284));
    NOR2X1 U36413 (.A1(n34159), .A2(n32035), .ZN(N49285));
    NOR2X1 U36414 (.A1(n34550), .A2(n24011), .ZN(N49286));
    NOR2X1 U36415 (.A1(n28503), .A2(n26740), .ZN(N49287));
    NOR2X1 U36416 (.A1(n34573), .A2(n30690), .ZN(N49288));
    INVX1 U36417 (.I(n14369), .ZN(N49289));
    INVX1 U36418 (.I(n39799), .ZN(N49290));
    NOR2X1 U36419 (.A1(n25754), .A2(n41617), .ZN(N49291));
    NANDX1 U36420 (.A1(N4105), .A2(n18227), .ZN(N49292));
    NANDX1 U36421 (.A1(n22013), .A2(n17388), .ZN(N49293));
    NOR2X1 U36422 (.A1(n22417), .A2(n21266), .ZN(N49294));
    NOR2X1 U36423 (.A1(n41694), .A2(N7632), .ZN(N49295));
    NANDX1 U36424 (.A1(n22061), .A2(n39667), .ZN(N49296));
    NANDX1 U36425 (.A1(n13138), .A2(N9885), .ZN(N49297));
    INVX1 U36426 (.I(n41641), .ZN(N49298));
    NANDX1 U36427 (.A1(N4616), .A2(n22421), .ZN(n49299));
    NOR2X1 U36428 (.A1(N1521), .A2(n36790), .ZN(N49300));
    NANDX1 U36429 (.A1(n41320), .A2(n27574), .ZN(N49301));
    NANDX1 U36430 (.A1(n29144), .A2(n30088), .ZN(N49302));
    NOR2X1 U36431 (.A1(n37050), .A2(n33662), .ZN(N49303));
    INVX1 U36432 (.I(N645), .ZN(N49304));
    INVX1 U36433 (.I(N1443), .ZN(N49305));
    NANDX1 U36434 (.A1(N6957), .A2(n32816), .ZN(N49306));
    NOR2X1 U36435 (.A1(n22196), .A2(N11404), .ZN(n49307));
    NANDX1 U36436 (.A1(n23733), .A2(n24542), .ZN(N49308));
    INVX1 U36437 (.I(n21400), .ZN(N49309));
    INVX1 U36438 (.I(N8130), .ZN(N49310));
    INVX1 U36439 (.I(n24490), .ZN(N49311));
    NOR2X1 U36440 (.A1(n27536), .A2(n17807), .ZN(N49312));
    NANDX1 U36441 (.A1(n15063), .A2(n35061), .ZN(N49313));
    NOR2X1 U36442 (.A1(N734), .A2(N11356), .ZN(N49314));
    NOR2X1 U36443 (.A1(n27463), .A2(N1545), .ZN(N49315));
    NANDX1 U36444 (.A1(n28107), .A2(N11175), .ZN(n49316));
    NANDX1 U36445 (.A1(N6544), .A2(n18131), .ZN(N49317));
    INVX1 U36446 (.I(n36085), .ZN(N49318));
    INVX1 U36447 (.I(n24152), .ZN(N49319));
    NOR2X1 U36448 (.A1(n43419), .A2(n38373), .ZN(N49320));
    INVX1 U36449 (.I(n21347), .ZN(N49321));
    INVX1 U36450 (.I(n41455), .ZN(N49322));
    NOR2X1 U36451 (.A1(n31779), .A2(N9313), .ZN(N49323));
    INVX1 U36452 (.I(n39266), .ZN(N49324));
    INVX1 U36453 (.I(n36168), .ZN(N49325));
    NANDX1 U36454 (.A1(N10890), .A2(n26581), .ZN(N49326));
    NOR2X1 U36455 (.A1(n20675), .A2(N10572), .ZN(N49327));
    NANDX1 U36456 (.A1(N9485), .A2(n38678), .ZN(N49328));
    NANDX1 U36457 (.A1(n32889), .A2(n34902), .ZN(n49329));
    INVX1 U36458 (.I(N2164), .ZN(N49330));
    NANDX1 U36459 (.A1(n18312), .A2(n15995), .ZN(N49331));
    INVX1 U36460 (.I(N7939), .ZN(n49332));
    NANDX1 U36461 (.A1(N4753), .A2(n29285), .ZN(N49333));
    NANDX1 U36462 (.A1(n35888), .A2(n22854), .ZN(N49334));
    INVX1 U36463 (.I(n34880), .ZN(N49335));
    INVX1 U36464 (.I(n25116), .ZN(N49336));
    INVX1 U36465 (.I(n26333), .ZN(n49337));
    NOR2X1 U36466 (.A1(N3888), .A2(N9442), .ZN(N49338));
    NANDX1 U36467 (.A1(n24562), .A2(N9693), .ZN(N49339));
    INVX1 U36468 (.I(n23726), .ZN(N49340));
    NANDX1 U36469 (.A1(N6713), .A2(N2822), .ZN(N49341));
    NANDX1 U36470 (.A1(n28171), .A2(n38138), .ZN(N49342));
    INVX1 U36471 (.I(N3010), .ZN(N49343));
    NANDX1 U36472 (.A1(n18100), .A2(N628), .ZN(N49344));
    INVX1 U36473 (.I(N12532), .ZN(N49345));
    NOR2X1 U36474 (.A1(n29418), .A2(N4947), .ZN(N49346));
    INVX1 U36475 (.I(n25588), .ZN(N49347));
    NOR2X1 U36476 (.A1(n42931), .A2(n40383), .ZN(N49348));
    INVX1 U36477 (.I(n15471), .ZN(N49349));
    NOR2X1 U36478 (.A1(n36712), .A2(n14592), .ZN(N49350));
    NOR2X1 U36479 (.A1(N7482), .A2(n24284), .ZN(N49351));
    NOR2X1 U36480 (.A1(n20887), .A2(N8542), .ZN(N49352));
    NOR2X1 U36481 (.A1(n23709), .A2(n27700), .ZN(N49353));
    NOR2X1 U36482 (.A1(n18374), .A2(n20580), .ZN(N49354));
    INVX1 U36483 (.I(n29033), .ZN(N49355));
    INVX1 U36484 (.I(n35969), .ZN(N49356));
    INVX1 U36485 (.I(n40890), .ZN(N49357));
    INVX1 U36486 (.I(n26213), .ZN(N49358));
    NANDX1 U36487 (.A1(N11061), .A2(n41480), .ZN(N49359));
    INVX1 U36488 (.I(N199), .ZN(N49360));
    NANDX1 U36489 (.A1(n21223), .A2(n15669), .ZN(n49361));
    NANDX1 U36490 (.A1(N4142), .A2(n30261), .ZN(n49362));
    INVX1 U36491 (.I(N11623), .ZN(N49363));
    NANDX1 U36492 (.A1(n16477), .A2(n22190), .ZN(N49364));
    INVX1 U36493 (.I(n30958), .ZN(n49365));
    INVX1 U36494 (.I(n36993), .ZN(N49366));
    NOR2X1 U36495 (.A1(N10479), .A2(N3780), .ZN(N49367));
    INVX1 U36496 (.I(n29191), .ZN(N49368));
    NOR2X1 U36497 (.A1(N4181), .A2(n25986), .ZN(N49369));
    INVX1 U36498 (.I(n16269), .ZN(N49370));
    INVX1 U36499 (.I(n31919), .ZN(N49371));
    INVX1 U36500 (.I(N6733), .ZN(N49372));
    INVX1 U36501 (.I(N6887), .ZN(N49373));
    NOR2X1 U36502 (.A1(n41539), .A2(n22555), .ZN(N49374));
    NANDX1 U36503 (.A1(N2209), .A2(n42495), .ZN(N49375));
    NOR2X1 U36504 (.A1(N3511), .A2(n32927), .ZN(n49376));
    INVX1 U36505 (.I(n25700), .ZN(N49377));
    NANDX1 U36506 (.A1(N10516), .A2(n17805), .ZN(N49378));
    INVX1 U36507 (.I(n30332), .ZN(n49379));
    INVX1 U36508 (.I(n29198), .ZN(N49380));
    NANDX1 U36509 (.A1(N3682), .A2(n17863), .ZN(N49381));
    NOR2X1 U36510 (.A1(n29667), .A2(N3946), .ZN(N49382));
    NANDX1 U36511 (.A1(n28072), .A2(n25544), .ZN(N49383));
    NOR2X1 U36512 (.A1(n24484), .A2(N2389), .ZN(N49384));
    INVX1 U36513 (.I(n15815), .ZN(N49385));
    NANDX1 U36514 (.A1(n34482), .A2(n13662), .ZN(N49386));
    NANDX1 U36515 (.A1(n23184), .A2(n20216), .ZN(N49387));
    INVX1 U36516 (.I(N12638), .ZN(N49388));
    NOR2X1 U36517 (.A1(N913), .A2(N1065), .ZN(N49389));
    INVX1 U36518 (.I(n18718), .ZN(N49390));
    INVX1 U36519 (.I(n19982), .ZN(N49391));
    NANDX1 U36520 (.A1(n35041), .A2(N8206), .ZN(N49392));
    NOR2X1 U36521 (.A1(n42583), .A2(N610), .ZN(N49393));
    NANDX1 U36522 (.A1(n36208), .A2(n32115), .ZN(N49394));
    INVX1 U36523 (.I(n18280), .ZN(N49395));
    NOR2X1 U36524 (.A1(n14998), .A2(N10348), .ZN(N49396));
    INVX1 U36525 (.I(n30812), .ZN(N49397));
    INVX1 U36526 (.I(n29771), .ZN(N49398));
    NOR2X1 U36527 (.A1(n25977), .A2(n42634), .ZN(N49399));
    INVX1 U36528 (.I(N1190), .ZN(N49400));
    INVX1 U36529 (.I(N350), .ZN(N49401));
    NANDX1 U36530 (.A1(n35696), .A2(n33472), .ZN(N49402));
    NOR2X1 U36531 (.A1(N8386), .A2(N9981), .ZN(N49403));
    NOR2X1 U36532 (.A1(n33106), .A2(N7866), .ZN(N49404));
    NOR2X1 U36533 (.A1(n21897), .A2(n41627), .ZN(N49405));
    NOR2X1 U36534 (.A1(n14632), .A2(n30269), .ZN(N49406));
    INVX1 U36535 (.I(n22591), .ZN(N49407));
    NOR2X1 U36536 (.A1(n34852), .A2(n32938), .ZN(N49408));
    INVX1 U36537 (.I(N11871), .ZN(N49409));
    INVX1 U36538 (.I(n28371), .ZN(N49410));
    NANDX1 U36539 (.A1(N5604), .A2(n27532), .ZN(N49411));
    INVX1 U36540 (.I(n39945), .ZN(N49412));
    NOR2X1 U36541 (.A1(n36628), .A2(n31726), .ZN(N49413));
    NOR2X1 U36542 (.A1(n26627), .A2(n31905), .ZN(N49414));
    NANDX1 U36543 (.A1(n26287), .A2(n25291), .ZN(N49415));
    INVX1 U36544 (.I(n34152), .ZN(N49416));
    NOR2X1 U36545 (.A1(n20509), .A2(n32307), .ZN(N49417));
    NANDX1 U36546 (.A1(n35141), .A2(N8783), .ZN(N49418));
    INVX1 U36547 (.I(N3939), .ZN(N49419));
    NOR2X1 U36548 (.A1(n25180), .A2(n26557), .ZN(N49420));
    NOR2X1 U36549 (.A1(n26731), .A2(N6184), .ZN(n49421));
    INVX1 U36550 (.I(n29281), .ZN(N49422));
    INVX1 U36551 (.I(n33444), .ZN(N49423));
    NOR2X1 U36552 (.A1(n41411), .A2(N8662), .ZN(N49424));
    NANDX1 U36553 (.A1(n29664), .A2(n29896), .ZN(N49425));
    NOR2X1 U36554 (.A1(n18096), .A2(n38875), .ZN(N49426));
    NOR2X1 U36555 (.A1(n33066), .A2(n37487), .ZN(n49427));
    NANDX1 U36556 (.A1(n17671), .A2(n14524), .ZN(N49428));
    INVX1 U36557 (.I(n31616), .ZN(N49429));
    INVX1 U36558 (.I(n35812), .ZN(N49430));
    NOR2X1 U36559 (.A1(n43282), .A2(N4433), .ZN(N49431));
    INVX1 U36560 (.I(n26366), .ZN(N49432));
    NANDX1 U36561 (.A1(n20062), .A2(n32549), .ZN(N49433));
    NOR2X1 U36562 (.A1(n39022), .A2(n34015), .ZN(N49434));
    NANDX1 U36563 (.A1(n17637), .A2(n21633), .ZN(N49435));
    INVX1 U36564 (.I(n22559), .ZN(N49436));
    NANDX1 U36565 (.A1(N6094), .A2(N10635), .ZN(N49437));
    NANDX1 U36566 (.A1(N1496), .A2(n24998), .ZN(N49438));
    NANDX1 U36567 (.A1(n38982), .A2(n19721), .ZN(N49439));
    NOR2X1 U36568 (.A1(N10033), .A2(N3277), .ZN(n49440));
    NANDX1 U36569 (.A1(n39056), .A2(n39088), .ZN(N49441));
    NANDX1 U36570 (.A1(n38866), .A2(N49), .ZN(N49442));
    NANDX1 U36571 (.A1(N11439), .A2(n25495), .ZN(N49443));
    NOR2X1 U36572 (.A1(n33668), .A2(n13380), .ZN(N49444));
    NANDX1 U36573 (.A1(n13890), .A2(n34709), .ZN(N49445));
    NANDX1 U36574 (.A1(n35523), .A2(N10907), .ZN(N49446));
    NOR2X1 U36575 (.A1(n43347), .A2(n17000), .ZN(N49447));
    NANDX1 U36576 (.A1(N5154), .A2(N8175), .ZN(N49448));
    INVX1 U36577 (.I(N27), .ZN(N49449));
    INVX1 U36578 (.I(n42366), .ZN(N49450));
    NOR2X1 U36579 (.A1(N3397), .A2(N2171), .ZN(N49451));
    NANDX1 U36580 (.A1(n42452), .A2(n30938), .ZN(N49452));
    INVX1 U36581 (.I(n27525), .ZN(N49453));
    INVX1 U36582 (.I(n31208), .ZN(N49454));
    NANDX1 U36583 (.A1(N2688), .A2(n13438), .ZN(n49455));
    NOR2X1 U36584 (.A1(N5748), .A2(n24369), .ZN(N49456));
    NANDX1 U36585 (.A1(n30136), .A2(N9465), .ZN(N49457));
    NOR2X1 U36586 (.A1(n41042), .A2(N6798), .ZN(n49458));
    NOR2X1 U36587 (.A1(N4249), .A2(n14766), .ZN(N49459));
    NOR2X1 U36588 (.A1(N12423), .A2(n37412), .ZN(N49460));
    NOR2X1 U36589 (.A1(n16106), .A2(n36305), .ZN(N49461));
    NOR2X1 U36590 (.A1(N9182), .A2(n38475), .ZN(N49462));
    NANDX1 U36591 (.A1(n41314), .A2(n25941), .ZN(N49463));
    NANDX1 U36592 (.A1(n15046), .A2(N3134), .ZN(N49464));
    INVX1 U36593 (.I(N217), .ZN(N49465));
    INVX1 U36594 (.I(N7964), .ZN(n49466));
    NOR2X1 U36595 (.A1(N1249), .A2(n32332), .ZN(N49467));
    NOR2X1 U36596 (.A1(n31384), .A2(n31476), .ZN(N49468));
    NOR2X1 U36597 (.A1(n28953), .A2(n38274), .ZN(N49469));
    INVX1 U36598 (.I(n33201), .ZN(N49470));
    NOR2X1 U36599 (.A1(n25625), .A2(N2151), .ZN(N49471));
    NANDX1 U36600 (.A1(n24496), .A2(N7936), .ZN(n49472));
    NOR2X1 U36601 (.A1(n35937), .A2(N6798), .ZN(N49473));
    NANDX1 U36602 (.A1(n17162), .A2(N4639), .ZN(N49474));
    INVX1 U36603 (.I(n23953), .ZN(N49475));
    NANDX1 U36604 (.A1(n22607), .A2(N8159), .ZN(N49476));
    INVX1 U36605 (.I(n18108), .ZN(N49477));
    NANDX1 U36606 (.A1(n18315), .A2(n19356), .ZN(N49478));
    NANDX1 U36607 (.A1(n16305), .A2(n40419), .ZN(N49479));
    NOR2X1 U36608 (.A1(n18433), .A2(n25899), .ZN(N49480));
    NANDX1 U36609 (.A1(n34892), .A2(N5307), .ZN(N49481));
    NANDX1 U36610 (.A1(N6724), .A2(n40609), .ZN(n49482));
    INVX1 U36611 (.I(n20899), .ZN(N49483));
    NANDX1 U36612 (.A1(N1580), .A2(n13364), .ZN(N49484));
    NOR2X1 U36613 (.A1(N5433), .A2(n30525), .ZN(N49485));
    NOR2X1 U36614 (.A1(n24905), .A2(N686), .ZN(N49486));
    NOR2X1 U36615 (.A1(N4039), .A2(N8844), .ZN(N49487));
    NOR2X1 U36616 (.A1(N11826), .A2(n14646), .ZN(N49488));
    NOR2X1 U36617 (.A1(n20861), .A2(n32139), .ZN(N49489));
    INVX1 U36618 (.I(n17807), .ZN(N49490));
    NOR2X1 U36619 (.A1(n14070), .A2(N233), .ZN(N49491));
    NOR2X1 U36620 (.A1(n38641), .A2(n38691), .ZN(N49492));
    INVX1 U36621 (.I(n35044), .ZN(N49493));
    NOR2X1 U36622 (.A1(N9566), .A2(N12470), .ZN(N49494));
    NANDX1 U36623 (.A1(N826), .A2(n25833), .ZN(N49495));
    NANDX1 U36624 (.A1(N6258), .A2(n12886), .ZN(N49496));
    NANDX1 U36625 (.A1(n31162), .A2(N3251), .ZN(N49497));
    INVX1 U36626 (.I(n24881), .ZN(N49498));
    INVX1 U36627 (.I(n17074), .ZN(N49499));
    NANDX1 U36628 (.A1(n16419), .A2(N6726), .ZN(N49500));
    INVX1 U36629 (.I(N5085), .ZN(N49501));
    NOR2X1 U36630 (.A1(n31901), .A2(n42720), .ZN(N49502));
    INVX1 U36631 (.I(n21814), .ZN(N49503));
    NOR2X1 U36632 (.A1(N1280), .A2(n17032), .ZN(N49504));
    INVX1 U36633 (.I(n36323), .ZN(n49505));
    INVX1 U36634 (.I(n30429), .ZN(N49506));
    NANDX1 U36635 (.A1(N9005), .A2(n31254), .ZN(N49507));
    INVX1 U36636 (.I(n20491), .ZN(N49508));
    NOR2X1 U36637 (.A1(n23398), .A2(n17524), .ZN(N49509));
    NOR2X1 U36638 (.A1(n26648), .A2(n30107), .ZN(N49510));
    INVX1 U36639 (.I(n28422), .ZN(N49511));
    NOR2X1 U36640 (.A1(n22674), .A2(N1368), .ZN(N49512));
    INVX1 U36641 (.I(n26448), .ZN(N49513));
    NANDX1 U36642 (.A1(n35628), .A2(N4557), .ZN(N49514));
    NOR2X1 U36643 (.A1(n41740), .A2(n26370), .ZN(N49515));
    NANDX1 U36644 (.A1(n32699), .A2(n33081), .ZN(N49516));
    NOR2X1 U36645 (.A1(n15230), .A2(n21827), .ZN(N49517));
    INVX1 U36646 (.I(N10230), .ZN(N49518));
    NOR2X1 U36647 (.A1(n40672), .A2(n20742), .ZN(N49519));
    INVX1 U36648 (.I(n24390), .ZN(N49520));
    INVX1 U36649 (.I(n15053), .ZN(N49521));
    INVX1 U36650 (.I(n16995), .ZN(N49522));
    INVX1 U36651 (.I(N4598), .ZN(N49523));
    NANDX1 U36652 (.A1(n28227), .A2(n16952), .ZN(N49524));
    INVX1 U36653 (.I(n18020), .ZN(N49525));
    INVX1 U36654 (.I(n22276), .ZN(N49526));
    NOR2X1 U36655 (.A1(N4483), .A2(N7335), .ZN(N49527));
    INVX1 U36656 (.I(n20532), .ZN(N49528));
    NOR2X1 U36657 (.A1(n41141), .A2(n43293), .ZN(N49529));
    NOR2X1 U36658 (.A1(n12898), .A2(N11327), .ZN(N49530));
    NOR2X1 U36659 (.A1(N12807), .A2(n31838), .ZN(N49531));
    NOR2X1 U36660 (.A1(n33549), .A2(n29367), .ZN(N49532));
    NANDX1 U36661 (.A1(n34216), .A2(n34099), .ZN(N49533));
    NOR2X1 U36662 (.A1(N7738), .A2(n15146), .ZN(N49534));
    NANDX1 U36663 (.A1(n42834), .A2(n33053), .ZN(N49535));
    NOR2X1 U36664 (.A1(n35825), .A2(N7600), .ZN(N49536));
    INVX1 U36665 (.I(n14628), .ZN(N49537));
    INVX1 U36666 (.I(n20043), .ZN(N49538));
    INVX1 U36667 (.I(n15897), .ZN(N49539));
    NOR2X1 U36668 (.A1(n30894), .A2(N3246), .ZN(N49540));
    NOR2X1 U36669 (.A1(n39455), .A2(N5823), .ZN(N49541));
    INVX1 U36670 (.I(n24281), .ZN(N49542));
    NANDX1 U36671 (.A1(n29766), .A2(n29139), .ZN(N49543));
    INVX1 U36672 (.I(N5340), .ZN(N49544));
    INVX1 U36673 (.I(n32601), .ZN(N49545));
    NOR2X1 U36674 (.A1(n29638), .A2(n30018), .ZN(N49546));
    NANDX1 U36675 (.A1(n38640), .A2(n19059), .ZN(N49547));
    NOR2X1 U36676 (.A1(n21121), .A2(N11411), .ZN(N49548));
    INVX1 U36677 (.I(n36681), .ZN(N49549));
    NANDX1 U36678 (.A1(n38578), .A2(n13251), .ZN(N49550));
    NANDX1 U36679 (.A1(N11002), .A2(N32), .ZN(N49551));
    NANDX1 U36680 (.A1(n14247), .A2(n30106), .ZN(N49552));
    INVX1 U36681 (.I(n20070), .ZN(n49553));
    NOR2X1 U36682 (.A1(n24723), .A2(n28379), .ZN(n49554));
    NOR2X1 U36683 (.A1(N10389), .A2(n26764), .ZN(N49555));
    NANDX1 U36684 (.A1(n25302), .A2(N5572), .ZN(N49556));
    INVX1 U36685 (.I(N1147), .ZN(N49557));
    INVX1 U36686 (.I(n18614), .ZN(N49558));
    NANDX1 U36687 (.A1(N856), .A2(n42137), .ZN(N49559));
    NANDX1 U36688 (.A1(N1946), .A2(n19468), .ZN(N49560));
    NOR2X1 U36689 (.A1(n17664), .A2(n14573), .ZN(n49561));
    NANDX1 U36690 (.A1(n34702), .A2(n25574), .ZN(N49562));
    INVX1 U36691 (.I(N6010), .ZN(N49563));
    NANDX1 U36692 (.A1(n33390), .A2(N6451), .ZN(N49564));
    NOR2X1 U36693 (.A1(N7631), .A2(n31173), .ZN(N49565));
    INVX1 U36694 (.I(N1317), .ZN(N49566));
    NOR2X1 U36695 (.A1(N7447), .A2(n33494), .ZN(N49567));
    NOR2X1 U36696 (.A1(n13018), .A2(n18164), .ZN(N49568));
    NANDX1 U36697 (.A1(n38286), .A2(n26458), .ZN(N49569));
    INVX1 U36698 (.I(n39141), .ZN(N49570));
    NOR2X1 U36699 (.A1(N7325), .A2(n41087), .ZN(N49571));
    INVX1 U36700 (.I(N7648), .ZN(N49572));
    NANDX1 U36701 (.A1(N5369), .A2(N10900), .ZN(N49573));
    INVX1 U36702 (.I(n30943), .ZN(N49574));
    NANDX1 U36703 (.A1(n35348), .A2(N6651), .ZN(N49575));
    INVX1 U36704 (.I(n41799), .ZN(N49576));
    INVX1 U36705 (.I(N1411), .ZN(N49577));
    NOR2X1 U36706 (.A1(n26583), .A2(n35879), .ZN(N49578));
    NOR2X1 U36707 (.A1(n34029), .A2(n25900), .ZN(N49579));
    NOR2X1 U36708 (.A1(n36726), .A2(n33744), .ZN(N49580));
    NANDX1 U36709 (.A1(n31539), .A2(n16729), .ZN(N49581));
    NANDX1 U36710 (.A1(n16888), .A2(n31530), .ZN(N49582));
    INVX1 U36711 (.I(N4182), .ZN(N49583));
    NOR2X1 U36712 (.A1(n18455), .A2(N9139), .ZN(N49584));
    NANDX1 U36713 (.A1(n29354), .A2(n38477), .ZN(N49585));
    NANDX1 U36714 (.A1(N66), .A2(n30353), .ZN(N49586));
    NOR2X1 U36715 (.A1(n37318), .A2(n18359), .ZN(N49587));
    INVX1 U36716 (.I(n38729), .ZN(n49588));
    INVX1 U36717 (.I(n40504), .ZN(N49589));
    NANDX1 U36718 (.A1(n34164), .A2(n20740), .ZN(N49590));
    INVX1 U36719 (.I(n33541), .ZN(N49591));
    NANDX1 U36720 (.A1(n36986), .A2(N3661), .ZN(N49592));
    INVX1 U36721 (.I(N10242), .ZN(N49593));
    INVX1 U36722 (.I(N8627), .ZN(N49594));
    INVX1 U36723 (.I(n28271), .ZN(N49595));
    NOR2X1 U36724 (.A1(N10305), .A2(N3253), .ZN(N49596));
    NANDX1 U36725 (.A1(n27680), .A2(n22286), .ZN(N49597));
    NOR2X1 U36726 (.A1(n32524), .A2(N12031), .ZN(N49598));
    INVX1 U36727 (.I(n33699), .ZN(N49599));
    NOR2X1 U36728 (.A1(n34700), .A2(N4148), .ZN(N49600));
    NOR2X1 U36729 (.A1(N8125), .A2(n34332), .ZN(N49601));
    INVX1 U36730 (.I(n31968), .ZN(N49602));
    NOR2X1 U36731 (.A1(n14869), .A2(n22036), .ZN(N49603));
    NANDX1 U36732 (.A1(n41534), .A2(n25697), .ZN(N49604));
    NOR2X1 U36733 (.A1(N8303), .A2(n32840), .ZN(N49605));
    NOR2X1 U36734 (.A1(n29434), .A2(n17638), .ZN(N49606));
    NOR2X1 U36735 (.A1(n39738), .A2(N10570), .ZN(N49607));
    INVX1 U36736 (.I(n23945), .ZN(N49608));
    NOR2X1 U36737 (.A1(N5418), .A2(N2677), .ZN(N49609));
    NOR2X1 U36738 (.A1(n21760), .A2(n36375), .ZN(N49610));
    NANDX1 U36739 (.A1(N2667), .A2(n30202), .ZN(N49611));
    NANDX1 U36740 (.A1(N10791), .A2(n21061), .ZN(N49612));
    NANDX1 U36741 (.A1(n42759), .A2(n32660), .ZN(N49613));
    INVX1 U36742 (.I(n21322), .ZN(N49614));
    NANDX1 U36743 (.A1(n35170), .A2(n36698), .ZN(n49615));
    INVX1 U36744 (.I(n33153), .ZN(N49616));
    NANDX1 U36745 (.A1(n16785), .A2(n19114), .ZN(N49617));
    NOR2X1 U36746 (.A1(n24588), .A2(N5059), .ZN(N49618));
    NANDX1 U36747 (.A1(n33696), .A2(n18684), .ZN(N49619));
    NANDX1 U36748 (.A1(n28793), .A2(n21360), .ZN(N49620));
    NANDX1 U36749 (.A1(N7080), .A2(n14262), .ZN(n49621));
    INVX1 U36750 (.I(n42899), .ZN(N49622));
    INVX1 U36751 (.I(N1049), .ZN(n49623));
    NANDX1 U36752 (.A1(N11732), .A2(n23288), .ZN(N49624));
    NOR2X1 U36753 (.A1(N919), .A2(n16924), .ZN(N49625));
    NANDX1 U36754 (.A1(n38529), .A2(n41774), .ZN(N49626));
    NANDX1 U36755 (.A1(n39677), .A2(n31454), .ZN(n49627));
    INVX1 U36756 (.I(N2669), .ZN(N49628));
    INVX1 U36757 (.I(N9064), .ZN(N49629));
    NANDX1 U36758 (.A1(N1833), .A2(n42695), .ZN(N49630));
    NOR2X1 U36759 (.A1(n20516), .A2(N1596), .ZN(N49631));
    INVX1 U36760 (.I(n31555), .ZN(N49632));
    INVX1 U36761 (.I(n32711), .ZN(N49633));
    INVX1 U36762 (.I(N8329), .ZN(N49634));
    INVX1 U36763 (.I(n36487), .ZN(N49635));
    NANDX1 U36764 (.A1(n32033), .A2(N4746), .ZN(N49636));
    NANDX1 U36765 (.A1(n31216), .A2(n38816), .ZN(N49637));
    INVX1 U36766 (.I(N8248), .ZN(N49638));
    NANDX1 U36767 (.A1(n37569), .A2(N11657), .ZN(N49639));
    NANDX1 U36768 (.A1(n15230), .A2(n30811), .ZN(N49640));
    INVX1 U36769 (.I(N12004), .ZN(N49641));
    NOR2X1 U36770 (.A1(n29039), .A2(N3516), .ZN(n49642));
    NANDX1 U36771 (.A1(n25877), .A2(n13712), .ZN(N49643));
    INVX1 U36772 (.I(N8035), .ZN(N49644));
    NOR2X1 U36773 (.A1(N4793), .A2(n30425), .ZN(N49645));
    NANDX1 U36774 (.A1(n13121), .A2(n19089), .ZN(N49646));
    NANDX1 U36775 (.A1(N12177), .A2(n40802), .ZN(N49647));
    NANDX1 U36776 (.A1(n34520), .A2(n28545), .ZN(N49648));
    INVX1 U36777 (.I(n30315), .ZN(N49649));
    NANDX1 U36778 (.A1(n33303), .A2(n24411), .ZN(N49650));
    NANDX1 U36779 (.A1(n42738), .A2(n39640), .ZN(N49651));
    INVX1 U36780 (.I(N11369), .ZN(N49652));
    NOR2X1 U36781 (.A1(n34381), .A2(n40407), .ZN(N49653));
    INVX1 U36782 (.I(N9365), .ZN(n49654));
    NANDX1 U36783 (.A1(N4758), .A2(n29416), .ZN(N49655));
    NOR2X1 U36784 (.A1(N6551), .A2(n34208), .ZN(N49656));
    NANDX1 U36785 (.A1(n33520), .A2(n37008), .ZN(N49657));
    INVX1 U36786 (.I(N10031), .ZN(N49658));
    NANDX1 U36787 (.A1(n13575), .A2(n34759), .ZN(n49659));
    INVX1 U36788 (.I(n31799), .ZN(N49660));
    NOR2X1 U36789 (.A1(n16754), .A2(n14798), .ZN(N49661));
    NANDX1 U36790 (.A1(n30844), .A2(n32286), .ZN(N49662));
    NANDX1 U36791 (.A1(n27012), .A2(n37112), .ZN(N49663));
    NANDX1 U36792 (.A1(n14542), .A2(n28020), .ZN(N49664));
    INVX1 U36793 (.I(N5588), .ZN(N49665));
    INVX1 U36794 (.I(n23437), .ZN(N49666));
    NANDX1 U36795 (.A1(n13007), .A2(N490), .ZN(N49667));
    INVX1 U36796 (.I(n36894), .ZN(N49668));
    NANDX1 U36797 (.A1(n40095), .A2(n30429), .ZN(N49669));
    NANDX1 U36798 (.A1(N6654), .A2(n25820), .ZN(N49670));
    NOR2X1 U36799 (.A1(n31092), .A2(N12258), .ZN(n49671));
    NANDX1 U36800 (.A1(N11490), .A2(n29011), .ZN(N49672));
    INVX1 U36801 (.I(n25189), .ZN(N49673));
    INVX1 U36802 (.I(n42236), .ZN(N49674));
    INVX1 U36803 (.I(n33074), .ZN(N49675));
    NANDX1 U36804 (.A1(N8694), .A2(n37295), .ZN(N49676));
    NANDX1 U36805 (.A1(n19641), .A2(n42883), .ZN(N49677));
    NOR2X1 U36806 (.A1(n32757), .A2(n42907), .ZN(N49678));
    NANDX1 U36807 (.A1(n33246), .A2(n39162), .ZN(N49679));
    NOR2X1 U36808 (.A1(n30892), .A2(n25465), .ZN(N49680));
    INVX1 U36809 (.I(n34464), .ZN(N49681));
    NANDX1 U36810 (.A1(n35727), .A2(N8138), .ZN(N49682));
    NANDX1 U36811 (.A1(N4512), .A2(N3290), .ZN(N49683));
    NOR2X1 U36812 (.A1(n23203), .A2(N2920), .ZN(N49684));
    NANDX1 U36813 (.A1(n29265), .A2(n34835), .ZN(N49685));
    NOR2X1 U36814 (.A1(N8546), .A2(n16917), .ZN(n49686));
    NANDX1 U36815 (.A1(N2368), .A2(N6378), .ZN(N49687));
    NOR2X1 U36816 (.A1(n34930), .A2(n33222), .ZN(N49688));
    INVX1 U36817 (.I(n24045), .ZN(N49689));
    NANDX1 U36818 (.A1(N6887), .A2(n19734), .ZN(N49690));
    INVX1 U36819 (.I(n27459), .ZN(N49691));
    INVX1 U36820 (.I(n18986), .ZN(N49692));
    NOR2X1 U36821 (.A1(n23523), .A2(N920), .ZN(N49693));
    NOR2X1 U36822 (.A1(n22620), .A2(n38584), .ZN(N49694));
    NANDX1 U36823 (.A1(n33205), .A2(n18314), .ZN(N49695));
    NANDX1 U36824 (.A1(n25507), .A2(n37258), .ZN(N49696));
    NANDX1 U36825 (.A1(N2170), .A2(N2331), .ZN(N49697));
    NANDX1 U36826 (.A1(n20679), .A2(n37850), .ZN(N49698));
    NANDX1 U36827 (.A1(n15355), .A2(n29308), .ZN(N49699));
    NOR2X1 U36828 (.A1(n32468), .A2(n43032), .ZN(N49700));
    INVX1 U36829 (.I(n39355), .ZN(N49701));
    NANDX1 U36830 (.A1(n13960), .A2(n23341), .ZN(N49702));
    INVX1 U36831 (.I(n32945), .ZN(N49703));
    INVX1 U36832 (.I(n23901), .ZN(n49704));
    NANDX1 U36833 (.A1(N4264), .A2(N3048), .ZN(N49705));
    NANDX1 U36834 (.A1(n13499), .A2(n36253), .ZN(N49706));
    INVX1 U36835 (.I(n25654), .ZN(N49707));
    NANDX1 U36836 (.A1(n20434), .A2(n18852), .ZN(N49708));
    NANDX1 U36837 (.A1(N12444), .A2(n28966), .ZN(N49709));
    INVX1 U36838 (.I(N6821), .ZN(N49710));
    NOR2X1 U36839 (.A1(n25529), .A2(n25808), .ZN(N49711));
    NANDX1 U36840 (.A1(n14525), .A2(n25367), .ZN(N49712));
    INVX1 U36841 (.I(N87), .ZN(N49713));
    INVX1 U36842 (.I(N6426), .ZN(N49714));
    INVX1 U36843 (.I(n34718), .ZN(N49715));
    NANDX1 U36844 (.A1(n21744), .A2(n15146), .ZN(N49716));
    NOR2X1 U36845 (.A1(n15687), .A2(n18194), .ZN(N49717));
    NANDX1 U36846 (.A1(n29185), .A2(N654), .ZN(N49718));
    NANDX1 U36847 (.A1(N1047), .A2(n41772), .ZN(N49719));
    NOR2X1 U36848 (.A1(n19898), .A2(n31268), .ZN(N49720));
    NANDX1 U36849 (.A1(n38543), .A2(n41442), .ZN(N49721));
    INVX1 U36850 (.I(n30207), .ZN(N49722));
    INVX1 U36851 (.I(N12345), .ZN(N49723));
    NOR2X1 U36852 (.A1(n17383), .A2(n27392), .ZN(N49724));
    NOR2X1 U36853 (.A1(n17469), .A2(N7939), .ZN(N49725));
    NANDX1 U36854 (.A1(n40895), .A2(n42656), .ZN(N49726));
    INVX1 U36855 (.I(N8846), .ZN(N49727));
    NANDX1 U36856 (.A1(N1063), .A2(n24532), .ZN(N49728));
    INVX1 U36857 (.I(n28839), .ZN(N49729));
    NANDX1 U36858 (.A1(n22855), .A2(n29472), .ZN(N49730));
    NANDX1 U36859 (.A1(N10835), .A2(N7065), .ZN(N49731));
    INVX1 U36860 (.I(n42102), .ZN(N49732));
    NANDX1 U36861 (.A1(N5617), .A2(n40072), .ZN(N49733));
    NOR2X1 U36862 (.A1(n35824), .A2(n42930), .ZN(N49734));
    NOR2X1 U36863 (.A1(n32976), .A2(n16840), .ZN(N49735));
    INVX1 U36864 (.I(n32914), .ZN(N49736));
    NANDX1 U36865 (.A1(n20992), .A2(n28957), .ZN(N49737));
    NANDX1 U36866 (.A1(n20175), .A2(n20897), .ZN(n49738));
    NANDX1 U36867 (.A1(n24184), .A2(N11639), .ZN(N49739));
    INVX1 U36868 (.I(N2913), .ZN(N49740));
    NOR2X1 U36869 (.A1(N917), .A2(n15448), .ZN(N49741));
    NANDX1 U36870 (.A1(N1887), .A2(n26282), .ZN(N49742));
    INVX1 U36871 (.I(N12433), .ZN(N49743));
    NANDX1 U36872 (.A1(N10002), .A2(n18050), .ZN(N49744));
    INVX1 U36873 (.I(n37112), .ZN(N49745));
    NOR2X1 U36874 (.A1(N10647), .A2(n22775), .ZN(N49746));
    INVX1 U36875 (.I(n27486), .ZN(N49747));
    NOR2X1 U36876 (.A1(n22497), .A2(N8001), .ZN(N49748));
    NOR2X1 U36877 (.A1(n41133), .A2(n29410), .ZN(N49749));
    NOR2X1 U36878 (.A1(N8237), .A2(n16192), .ZN(N49750));
    NOR2X1 U36879 (.A1(n19876), .A2(N6865), .ZN(N49751));
    NOR2X1 U36880 (.A1(N6561), .A2(N7782), .ZN(N49752));
    INVX1 U36881 (.I(N12397), .ZN(N49753));
    NOR2X1 U36882 (.A1(n27914), .A2(n35617), .ZN(N49754));
    NANDX1 U36883 (.A1(n42504), .A2(N2147), .ZN(N49755));
    NANDX1 U36884 (.A1(N10222), .A2(n28938), .ZN(N49756));
    INVX1 U36885 (.I(n20868), .ZN(N49757));
    INVX1 U36886 (.I(N9172), .ZN(N49758));
    INVX1 U36887 (.I(n33748), .ZN(N49759));
    NOR2X1 U36888 (.A1(N2562), .A2(n26455), .ZN(N49760));
    NOR2X1 U36889 (.A1(n31972), .A2(n29016), .ZN(N49761));
    INVX1 U36890 (.I(n37843), .ZN(n49762));
    INVX1 U36891 (.I(n36800), .ZN(N49763));
    NANDX1 U36892 (.A1(n41946), .A2(n43360), .ZN(n49764));
    INVX1 U36893 (.I(n33258), .ZN(N49765));
    NANDX1 U36894 (.A1(N8364), .A2(N7379), .ZN(n49766));
    NOR2X1 U36895 (.A1(n20143), .A2(N6410), .ZN(N49767));
    INVX1 U36896 (.I(n39652), .ZN(N49768));
    INVX1 U36897 (.I(n14872), .ZN(N49769));
    NOR2X1 U36898 (.A1(n37499), .A2(N12791), .ZN(N49770));
    NANDX1 U36899 (.A1(n32060), .A2(n36218), .ZN(N49771));
    INVX1 U36900 (.I(n34621), .ZN(N49772));
    NOR2X1 U36901 (.A1(n21823), .A2(N12800), .ZN(N49773));
    NANDX1 U36902 (.A1(N5595), .A2(N7171), .ZN(N49774));
    NANDX1 U36903 (.A1(n32074), .A2(N8406), .ZN(n49775));
    NANDX1 U36904 (.A1(n31961), .A2(N7102), .ZN(N49776));
    NOR2X1 U36905 (.A1(n33924), .A2(n15465), .ZN(N49777));
    NOR2X1 U36906 (.A1(n28031), .A2(n25287), .ZN(N49778));
    INVX1 U36907 (.I(N3645), .ZN(N49779));
    NOR2X1 U36908 (.A1(N4748), .A2(n18516), .ZN(N49780));
    NOR2X1 U36909 (.A1(n31926), .A2(n31306), .ZN(N49781));
    NANDX1 U36910 (.A1(n20513), .A2(n13732), .ZN(N49782));
    NANDX1 U36911 (.A1(N1341), .A2(n22611), .ZN(N49783));
    NANDX1 U36912 (.A1(n14141), .A2(n17034), .ZN(N49784));
    NOR2X1 U36913 (.A1(n21311), .A2(n13425), .ZN(N49785));
    INVX1 U36914 (.I(n19396), .ZN(n49786));
    NOR2X1 U36915 (.A1(n38532), .A2(n26497), .ZN(N49787));
    NANDX1 U36916 (.A1(n28983), .A2(n31641), .ZN(N49788));
    NANDX1 U36917 (.A1(N3222), .A2(n13455), .ZN(N49789));
    NOR2X1 U36918 (.A1(N6866), .A2(n24601), .ZN(N49790));
    NANDX1 U36919 (.A1(n15061), .A2(N8042), .ZN(N49791));
    NOR2X1 U36920 (.A1(n36046), .A2(n16422), .ZN(N49792));
    NANDX1 U36921 (.A1(N6305), .A2(n27616), .ZN(n49793));
    NOR2X1 U36922 (.A1(n28916), .A2(N6841), .ZN(N49794));
    INVX1 U36923 (.I(N2477), .ZN(N49795));
    NANDX1 U36924 (.A1(n27968), .A2(n15902), .ZN(N49796));
    INVX1 U36925 (.I(N3891), .ZN(N49797));
    NANDX1 U36926 (.A1(n36762), .A2(n30387), .ZN(N49798));
    NANDX1 U36927 (.A1(N11953), .A2(N8235), .ZN(N49799));
    NOR2X1 U36928 (.A1(N4854), .A2(n21690), .ZN(N49800));
    NOR2X1 U36929 (.A1(N1399), .A2(N2818), .ZN(N49801));
    INVX1 U36930 (.I(n16459), .ZN(N49802));
    INVX1 U36931 (.I(n27506), .ZN(N49803));
    NANDX1 U36932 (.A1(n27280), .A2(n39323), .ZN(N49804));
    INVX1 U36933 (.I(N1103), .ZN(N49805));
    NOR2X1 U36934 (.A1(n33932), .A2(N7943), .ZN(N49806));
    NOR2X1 U36935 (.A1(n26088), .A2(n43074), .ZN(N49807));
    NANDX1 U36936 (.A1(n31669), .A2(n30984), .ZN(N49808));
    NOR2X1 U36937 (.A1(n35219), .A2(n13953), .ZN(N49809));
    NOR2X1 U36938 (.A1(N11066), .A2(n25905), .ZN(N49810));
    NOR2X1 U36939 (.A1(n38181), .A2(n20438), .ZN(N49811));
    NOR2X1 U36940 (.A1(n30250), .A2(n21836), .ZN(N49812));
    INVX1 U36941 (.I(N2338), .ZN(N49813));
    NOR2X1 U36942 (.A1(n13925), .A2(n29844), .ZN(N49814));
    NANDX1 U36943 (.A1(n30884), .A2(n25694), .ZN(N49815));
    NOR2X1 U36944 (.A1(n31987), .A2(n24382), .ZN(N49816));
    INVX1 U36945 (.I(n29609), .ZN(N49817));
    NOR2X1 U36946 (.A1(n27608), .A2(n29210), .ZN(N49818));
    NANDX1 U36947 (.A1(N5485), .A2(N6401), .ZN(N49819));
    INVX1 U36948 (.I(n40703), .ZN(N49820));
    NANDX1 U36949 (.A1(n35226), .A2(N8296), .ZN(N49821));
    NOR2X1 U36950 (.A1(n24107), .A2(n36156), .ZN(N49822));
    NANDX1 U36951 (.A1(n24356), .A2(N12613), .ZN(N49823));
    NOR2X1 U36952 (.A1(n27423), .A2(n14951), .ZN(N49824));
    INVX1 U36953 (.I(n41347), .ZN(N49825));
    NANDX1 U36954 (.A1(n25286), .A2(n18439), .ZN(N49826));
    NANDX1 U36955 (.A1(N3195), .A2(n40105), .ZN(N49827));
    NANDX1 U36956 (.A1(N4715), .A2(n26241), .ZN(N49828));
    NANDX1 U36957 (.A1(n22002), .A2(N1659), .ZN(N49829));
    INVX1 U36958 (.I(n27486), .ZN(N49830));
    NANDX1 U36959 (.A1(N2023), .A2(n14396), .ZN(N49831));
    NOR2X1 U36960 (.A1(n26929), .A2(n22691), .ZN(N49832));
    INVX1 U36961 (.I(N7563), .ZN(n49833));
    INVX1 U36962 (.I(n33781), .ZN(n49834));
    NOR2X1 U36963 (.A1(n17667), .A2(n14727), .ZN(N49835));
    NOR2X1 U36964 (.A1(n22297), .A2(n23647), .ZN(N49836));
    NANDX1 U36965 (.A1(n13298), .A2(N5460), .ZN(N49837));
    INVX1 U36966 (.I(n29993), .ZN(N49838));
    NOR2X1 U36967 (.A1(N8173), .A2(n17277), .ZN(N49839));
    INVX1 U36968 (.I(n24093), .ZN(N49840));
    NOR2X1 U36969 (.A1(n25050), .A2(n25751), .ZN(N49841));
    NOR2X1 U36970 (.A1(n42215), .A2(n33810), .ZN(N49842));
    INVX1 U36971 (.I(n13139), .ZN(N49843));
    NANDX1 U36972 (.A1(N10681), .A2(n25509), .ZN(N49844));
    NANDX1 U36973 (.A1(N7923), .A2(n20243), .ZN(N49845));
    NOR2X1 U36974 (.A1(n29521), .A2(n37910), .ZN(N49846));
    NOR2X1 U36975 (.A1(n35068), .A2(n16734), .ZN(N49847));
    INVX1 U36976 (.I(n28170), .ZN(N49848));
    NANDX1 U36977 (.A1(n42807), .A2(n39710), .ZN(N49849));
    NOR2X1 U36978 (.A1(n41140), .A2(n37562), .ZN(N49850));
    INVX1 U36979 (.I(n33868), .ZN(N49851));
    NANDX1 U36980 (.A1(N4003), .A2(N5125), .ZN(N49852));
    NANDX1 U36981 (.A1(n29205), .A2(N3867), .ZN(N49853));
    NOR2X1 U36982 (.A1(n12957), .A2(n17005), .ZN(N49854));
    NOR2X1 U36983 (.A1(n13318), .A2(n32194), .ZN(N49855));
    INVX1 U36984 (.I(N10920), .ZN(N49856));
    NOR2X1 U36985 (.A1(n17186), .A2(n40440), .ZN(N49857));
    INVX1 U36986 (.I(n41206), .ZN(N49858));
    NOR2X1 U36987 (.A1(n42967), .A2(n35080), .ZN(n49859));
    NANDX1 U36988 (.A1(n19206), .A2(n24094), .ZN(N49860));
    NOR2X1 U36989 (.A1(n15117), .A2(N11442), .ZN(N49861));
    NOR2X1 U36990 (.A1(n28304), .A2(N1837), .ZN(N49862));
    NANDX1 U36991 (.A1(n21986), .A2(n40113), .ZN(N49863));
    INVX1 U36992 (.I(N7718), .ZN(N49864));
    NOR2X1 U36993 (.A1(n41524), .A2(n20674), .ZN(N49865));
    INVX1 U36994 (.I(n20110), .ZN(N49866));
    NOR2X1 U36995 (.A1(n39385), .A2(n17682), .ZN(N49867));
    INVX1 U36996 (.I(n38028), .ZN(N49868));
    INVX1 U36997 (.I(n31558), .ZN(N49869));
    NOR2X1 U36998 (.A1(n22280), .A2(N9801), .ZN(N49870));
    NANDX1 U36999 (.A1(N3567), .A2(N5894), .ZN(N49871));
    NANDX1 U37000 (.A1(n17341), .A2(n41696), .ZN(N49872));
    NANDX1 U37001 (.A1(n28782), .A2(n17795), .ZN(N49873));
    NOR2X1 U37002 (.A1(n20298), .A2(N12077), .ZN(N49874));
    INVX1 U37003 (.I(n16938), .ZN(N49875));
    NANDX1 U37004 (.A1(n25665), .A2(N7124), .ZN(N49876));
    NOR2X1 U37005 (.A1(n36018), .A2(n14315), .ZN(N49877));
    INVX1 U37006 (.I(n16217), .ZN(N49878));
    NANDX1 U37007 (.A1(N1381), .A2(n40487), .ZN(N49879));
    INVX1 U37008 (.I(n25927), .ZN(N49880));
    NOR2X1 U37009 (.A1(n25571), .A2(n37886), .ZN(N49881));
    INVX1 U37010 (.I(N2381), .ZN(N49882));
    NOR2X1 U37011 (.A1(n23626), .A2(n41868), .ZN(N49883));
    NANDX1 U37012 (.A1(N11529), .A2(N9527), .ZN(N49884));
    NOR2X1 U37013 (.A1(n29323), .A2(N5489), .ZN(N49885));
    NANDX1 U37014 (.A1(n31079), .A2(n13116), .ZN(N49886));
    NANDX1 U37015 (.A1(N6937), .A2(n28460), .ZN(N49887));
    NANDX1 U37016 (.A1(n24319), .A2(n21005), .ZN(N49888));
    NANDX1 U37017 (.A1(N8018), .A2(n26901), .ZN(N49889));
    INVX1 U37018 (.I(n42550), .ZN(N49890));
    NANDX1 U37019 (.A1(N2070), .A2(n14684), .ZN(N49891));
    NANDX1 U37020 (.A1(n17320), .A2(N9097), .ZN(N49892));
    NANDX1 U37021 (.A1(n19700), .A2(n40228), .ZN(n49893));
    INVX1 U37022 (.I(n18095), .ZN(N49894));
    NANDX1 U37023 (.A1(n30940), .A2(n27621), .ZN(N49895));
    INVX1 U37024 (.I(n16790), .ZN(N49896));
    INVX1 U37025 (.I(N4862), .ZN(n49897));
    INVX1 U37026 (.I(n35904), .ZN(N49898));
    NOR2X1 U37027 (.A1(N1013), .A2(N10571), .ZN(N49899));
    INVX1 U37028 (.I(n15011), .ZN(n49900));
    INVX1 U37029 (.I(n23171), .ZN(N49901));
    NANDX1 U37030 (.A1(N4684), .A2(n30778), .ZN(n49902));
    INVX1 U37031 (.I(n18278), .ZN(N49903));
    NOR2X1 U37032 (.A1(n26468), .A2(N6652), .ZN(N49904));
    INVX1 U37033 (.I(n25244), .ZN(N49905));
    NANDX1 U37034 (.A1(n26393), .A2(N11680), .ZN(N49906));
    NOR2X1 U37035 (.A1(n34167), .A2(N3115), .ZN(N49907));
    NANDX1 U37036 (.A1(N7995), .A2(N7690), .ZN(N49908));
    INVX1 U37037 (.I(n30783), .ZN(N49909));
    NOR2X1 U37038 (.A1(n20182), .A2(n12894), .ZN(N49910));
    NOR2X1 U37039 (.A1(N10874), .A2(n23464), .ZN(N49911));
    INVX1 U37040 (.I(n25885), .ZN(N49912));
    NOR2X1 U37041 (.A1(n42314), .A2(n38592), .ZN(N49913));
    INVX1 U37042 (.I(n29619), .ZN(N49914));
    INVX1 U37043 (.I(N3567), .ZN(N49915));
    NANDX1 U37044 (.A1(n23052), .A2(n43370), .ZN(n49916));
    NANDX1 U37045 (.A1(N4824), .A2(N2336), .ZN(N49917));
    NANDX1 U37046 (.A1(n16503), .A2(n24184), .ZN(N49918));
    NANDX1 U37047 (.A1(N9297), .A2(n23180), .ZN(N49919));
    NOR2X1 U37048 (.A1(n16986), .A2(N5813), .ZN(N49920));
    NANDX1 U37049 (.A1(n19217), .A2(n15674), .ZN(N49921));
    NOR2X1 U37050 (.A1(n22891), .A2(n16227), .ZN(n49922));
    NOR2X1 U37051 (.A1(n42034), .A2(n42111), .ZN(N49923));
    INVX1 U37052 (.I(n30556), .ZN(N49924));
    NANDX1 U37053 (.A1(n42518), .A2(N6382), .ZN(N49925));
    NANDX1 U37054 (.A1(N2612), .A2(n15055), .ZN(N49926));
    NOR2X1 U37055 (.A1(n35662), .A2(n20100), .ZN(N49927));
    NOR2X1 U37056 (.A1(n37997), .A2(n41218), .ZN(N49928));
    NANDX1 U37057 (.A1(N8388), .A2(N9557), .ZN(N49929));
    NOR2X1 U37058 (.A1(n21247), .A2(n29363), .ZN(N49930));
    INVX1 U37059 (.I(n27059), .ZN(N49931));
    INVX1 U37060 (.I(n16105), .ZN(N49932));
    NANDX1 U37061 (.A1(n15207), .A2(n38995), .ZN(N49933));
    INVX1 U37062 (.I(n38038), .ZN(N49934));
    NOR2X1 U37063 (.A1(n36957), .A2(n41475), .ZN(N49935));
    NOR2X1 U37064 (.A1(n20395), .A2(n40521), .ZN(N49936));
    INVX1 U37065 (.I(N417), .ZN(N49937));
    NOR2X1 U37066 (.A1(n15115), .A2(N3491), .ZN(N49938));
    NOR2X1 U37067 (.A1(n35214), .A2(N11387), .ZN(N49939));
    NOR2X1 U37068 (.A1(n32959), .A2(n25466), .ZN(N49940));
    NOR2X1 U37069 (.A1(n32196), .A2(n15688), .ZN(N49941));
    NOR2X1 U37070 (.A1(N7766), .A2(N12576), .ZN(N49942));
    NOR2X1 U37071 (.A1(n23603), .A2(n28680), .ZN(N49943));
    NANDX1 U37072 (.A1(n38809), .A2(n13882), .ZN(N49944));
    NANDX1 U37073 (.A1(n23055), .A2(n41118), .ZN(N49945));
    INVX1 U37074 (.I(n21057), .ZN(N49946));
    INVX1 U37075 (.I(N11962), .ZN(N49947));
    INVX1 U37076 (.I(N12024), .ZN(N49948));
    INVX1 U37077 (.I(n40597), .ZN(N49949));
    NOR2X1 U37078 (.A1(N5549), .A2(N11805), .ZN(N49950));
    INVX1 U37079 (.I(n16935), .ZN(N49951));
    INVX1 U37080 (.I(n31198), .ZN(N49952));
    INVX1 U37081 (.I(n28282), .ZN(N49953));
    NOR2X1 U37082 (.A1(N4296), .A2(N3008), .ZN(N49954));
    INVX1 U37083 (.I(N6551), .ZN(N49955));
    NANDX1 U37084 (.A1(N7817), .A2(n24911), .ZN(N49956));
    INVX1 U37085 (.I(n36305), .ZN(N49957));
    INVX1 U37086 (.I(N3920), .ZN(N49958));
    INVX1 U37087 (.I(n26117), .ZN(N49959));
    NANDX1 U37088 (.A1(n26624), .A2(n27761), .ZN(N49960));
    NANDX1 U37089 (.A1(n34408), .A2(n39784), .ZN(N49961));
    NOR2X1 U37090 (.A1(n21212), .A2(n13130), .ZN(N49962));
    NANDX1 U37091 (.A1(n33017), .A2(n21689), .ZN(N49963));
    NANDX1 U37092 (.A1(N234), .A2(n42566), .ZN(N49964));
    NOR2X1 U37093 (.A1(n18195), .A2(n19015), .ZN(N49965));
    INVX1 U37094 (.I(n21202), .ZN(N49966));
    NANDX1 U37095 (.A1(N10802), .A2(n25995), .ZN(N49967));
    NANDX1 U37096 (.A1(n35712), .A2(N872), .ZN(n49968));
    NANDX1 U37097 (.A1(n20712), .A2(N4791), .ZN(N49969));
    NOR2X1 U37098 (.A1(n36508), .A2(N278), .ZN(N49970));
    INVX1 U37099 (.I(n20796), .ZN(n49971));
    INVX1 U37100 (.I(n39514), .ZN(N49972));
    NANDX1 U37101 (.A1(n27552), .A2(n17253), .ZN(N49973));
    NANDX1 U37102 (.A1(N9454), .A2(n39949), .ZN(N49974));
    NANDX1 U37103 (.A1(n31122), .A2(n29862), .ZN(N49975));
    NANDX1 U37104 (.A1(N8246), .A2(N4584), .ZN(N49976));
    NOR2X1 U37105 (.A1(N12497), .A2(n15466), .ZN(N49977));
    NANDX1 U37106 (.A1(n23299), .A2(n31140), .ZN(n49978));
    NOR2X1 U37107 (.A1(N5218), .A2(n32011), .ZN(N49979));
    NANDX1 U37108 (.A1(n15609), .A2(n36801), .ZN(N49980));
    NANDX1 U37109 (.A1(N8645), .A2(n26758), .ZN(N49981));
    NOR2X1 U37110 (.A1(n19120), .A2(n34483), .ZN(N49982));
    NOR2X1 U37111 (.A1(n15587), .A2(n18562), .ZN(N49983));
    INVX1 U37112 (.I(n25183), .ZN(n49984));
    NOR2X1 U37113 (.A1(N11489), .A2(n35827), .ZN(N49985));
    NOR2X1 U37114 (.A1(n41351), .A2(N12413), .ZN(N49986));
    NANDX1 U37115 (.A1(n35614), .A2(n41164), .ZN(N49987));
    NANDX1 U37116 (.A1(n40759), .A2(N9031), .ZN(N49988));
    INVX1 U37117 (.I(n28426), .ZN(N49989));
    NANDX1 U37118 (.A1(n33962), .A2(n16964), .ZN(n49990));
    INVX1 U37119 (.I(N6099), .ZN(N49991));
    NOR2X1 U37120 (.A1(N2685), .A2(N4423), .ZN(N49992));
    NANDX1 U37121 (.A1(n14724), .A2(n23542), .ZN(N49993));
    NANDX1 U37122 (.A1(n22803), .A2(n28809), .ZN(N49994));
    INVX1 U37123 (.I(n37815), .ZN(N49995));
    NOR2X1 U37124 (.A1(n33357), .A2(N5832), .ZN(N49996));
    INVX1 U37125 (.I(n38701), .ZN(N49997));
    NANDX1 U37126 (.A1(N4966), .A2(n31650), .ZN(N49998));
    NANDX1 U37127 (.A1(n35809), .A2(N3944), .ZN(N49999));
    NANDX1 U37128 (.A1(N1368), .A2(n32688), .ZN(N50000));
    NOR2X1 U37129 (.A1(N12141), .A2(N12858), .ZN(N50001));
    NANDX1 U37130 (.A1(n41044), .A2(n18956), .ZN(n50002));
    INVX1 U37131 (.I(n33409), .ZN(N50003));
    NANDX1 U37132 (.A1(n34268), .A2(n37812), .ZN(N50004));
    NANDX1 U37133 (.A1(n41688), .A2(n17142), .ZN(N50005));
    NOR2X1 U37134 (.A1(n13878), .A2(N11485), .ZN(N50006));
    INVX1 U37135 (.I(N3762), .ZN(N50007));
    NANDX1 U37136 (.A1(n14687), .A2(n32142), .ZN(N50008));
    NOR2X1 U37137 (.A1(n19652), .A2(n20319), .ZN(N50009));
    NANDX1 U37138 (.A1(N11988), .A2(n13943), .ZN(N50010));
    NOR2X1 U37139 (.A1(N3035), .A2(n36310), .ZN(N50011));
    INVX1 U37140 (.I(n15175), .ZN(N50012));
    INVX1 U37141 (.I(n22885), .ZN(N50013));
    NOR2X1 U37142 (.A1(n14330), .A2(n30423), .ZN(N50014));
    NANDX1 U37143 (.A1(n27387), .A2(N10898), .ZN(N50015));
    NOR2X1 U37144 (.A1(n20514), .A2(n42266), .ZN(N50016));
    INVX1 U37145 (.I(n32128), .ZN(N50017));
    NOR2X1 U37146 (.A1(n27839), .A2(N10789), .ZN(N50018));
    NOR2X1 U37147 (.A1(n34834), .A2(n25475), .ZN(N50019));
    INVX1 U37148 (.I(n24898), .ZN(N50020));
    NANDX1 U37149 (.A1(N4779), .A2(n33645), .ZN(N50021));
    INVX1 U37150 (.I(N8401), .ZN(N50022));
    NOR2X1 U37151 (.A1(N6356), .A2(N1239), .ZN(N50023));
    INVX1 U37152 (.I(N11211), .ZN(N50024));
    NANDX1 U37153 (.A1(n32450), .A2(N3317), .ZN(N50025));
    INVX1 U37154 (.I(N9080), .ZN(N50026));
    INVX1 U37155 (.I(n28009), .ZN(N50027));
    NOR2X1 U37156 (.A1(n38364), .A2(N5050), .ZN(N50028));
    NANDX1 U37157 (.A1(N11246), .A2(n37178), .ZN(n50029));
    INVX1 U37158 (.I(n39085), .ZN(N50030));
    INVX1 U37159 (.I(N6592), .ZN(N50031));
    NANDX1 U37160 (.A1(n19649), .A2(n34524), .ZN(N50032));
    INVX1 U37161 (.I(N10982), .ZN(N50033));
    NOR2X1 U37162 (.A1(n24876), .A2(N3983), .ZN(N50034));
    NANDX1 U37163 (.A1(n29443), .A2(N10339), .ZN(N50035));
    NOR2X1 U37164 (.A1(n39009), .A2(n21549), .ZN(N50036));
    NANDX1 U37165 (.A1(n17666), .A2(n24865), .ZN(N50037));
    NANDX1 U37166 (.A1(n26746), .A2(n43375), .ZN(N50038));
    INVX1 U37167 (.I(n26083), .ZN(N50039));
    NOR2X1 U37168 (.A1(n15121), .A2(n24213), .ZN(N50040));
    INVX1 U37169 (.I(n41978), .ZN(N50041));
    NOR2X1 U37170 (.A1(n34803), .A2(n25832), .ZN(N50042));
    INVX1 U37171 (.I(n21777), .ZN(N50043));
    INVX1 U37172 (.I(n22335), .ZN(N50044));
    NANDX1 U37173 (.A1(N2669), .A2(N7844), .ZN(N50045));
    NOR2X1 U37174 (.A1(N6652), .A2(N12074), .ZN(N50046));
    NANDX1 U37175 (.A1(N6670), .A2(n40374), .ZN(N50047));
    NOR2X1 U37176 (.A1(n28218), .A2(n21815), .ZN(N50048));
    INVX1 U37177 (.I(n42762), .ZN(N50049));
    INVX1 U37178 (.I(n32840), .ZN(N50050));
    NANDX1 U37179 (.A1(n13948), .A2(n15450), .ZN(N50051));
    INVX1 U37180 (.I(n18749), .ZN(n50052));
    INVX1 U37181 (.I(n22855), .ZN(N50053));
    INVX1 U37182 (.I(n20882), .ZN(N50054));
    NANDX1 U37183 (.A1(n43085), .A2(N8693), .ZN(N50055));
    INVX1 U37184 (.I(n24452), .ZN(N50056));
    NOR2X1 U37185 (.A1(n38649), .A2(n27121), .ZN(N50057));
    INVX1 U37186 (.I(n33059), .ZN(N50058));
    INVX1 U37187 (.I(n30304), .ZN(N50059));
    INVX1 U37188 (.I(n30121), .ZN(N50060));
    INVX1 U37189 (.I(N1868), .ZN(N50061));
    INVX1 U37190 (.I(N5547), .ZN(N50062));
    NANDX1 U37191 (.A1(n36987), .A2(n42576), .ZN(N50063));
    INVX1 U37192 (.I(n25858), .ZN(N50064));
    NANDX1 U37193 (.A1(N12778), .A2(n42674), .ZN(N50065));
    NOR2X1 U37194 (.A1(n42119), .A2(N11736), .ZN(N50066));
    NANDX1 U37195 (.A1(n19528), .A2(n15601), .ZN(N50067));
    INVX1 U37196 (.I(n17900), .ZN(N50068));
    NOR2X1 U37197 (.A1(N9005), .A2(n38606), .ZN(N50069));
    NOR2X1 U37198 (.A1(n25805), .A2(n23683), .ZN(N50070));
    NANDX1 U37199 (.A1(n38936), .A2(N10514), .ZN(N50071));
    NOR2X1 U37200 (.A1(n15264), .A2(n37719), .ZN(N50072));
    NANDX1 U37201 (.A1(N9489), .A2(n32945), .ZN(N50073));
    NOR2X1 U37202 (.A1(N3003), .A2(n21728), .ZN(N50074));
    NOR2X1 U37203 (.A1(n18540), .A2(n34779), .ZN(N50075));
    NANDX1 U37204 (.A1(n17741), .A2(N12785), .ZN(N50076));
    INVX1 U37205 (.I(n19156), .ZN(N50077));
    NOR2X1 U37206 (.A1(n36269), .A2(n34757), .ZN(N50078));
    INVX1 U37207 (.I(N376), .ZN(N50079));
    INVX1 U37208 (.I(n24434), .ZN(N50080));
    NOR2X1 U37209 (.A1(n37984), .A2(N6766), .ZN(N50081));
    NANDX1 U37210 (.A1(n43347), .A2(N2229), .ZN(N50082));
    NOR2X1 U37211 (.A1(n41509), .A2(n17492), .ZN(n50083));
    NANDX1 U37212 (.A1(n41538), .A2(n26980), .ZN(N50084));
    NANDX1 U37213 (.A1(N6056), .A2(n19662), .ZN(N50085));
    INVX1 U37214 (.I(N11374), .ZN(N50086));
    NOR2X1 U37215 (.A1(N5817), .A2(n19149), .ZN(N50087));
    NOR2X1 U37216 (.A1(n18601), .A2(n35890), .ZN(n50088));
    NOR2X1 U37217 (.A1(N6006), .A2(n18366), .ZN(N50089));
    INVX1 U37218 (.I(n31755), .ZN(N50090));
    NOR2X1 U37219 (.A1(n14154), .A2(N12716), .ZN(N50091));
    NANDX1 U37220 (.A1(n41817), .A2(N9161), .ZN(N50092));
    NANDX1 U37221 (.A1(n41691), .A2(N1069), .ZN(N50093));
    INVX1 U37222 (.I(n39728), .ZN(N50094));
    INVX1 U37223 (.I(n22982), .ZN(N50095));
    INVX1 U37224 (.I(n35219), .ZN(N50096));
    INVX1 U37225 (.I(n23209), .ZN(n50097));
    NANDX1 U37226 (.A1(n30274), .A2(n34582), .ZN(N50098));
    INVX1 U37227 (.I(n36090), .ZN(N50099));
    NOR2X1 U37228 (.A1(n20796), .A2(N899), .ZN(N50100));
    NOR2X1 U37229 (.A1(n31779), .A2(N6904), .ZN(N50101));
    INVX1 U37230 (.I(n13407), .ZN(N50102));
    NANDX1 U37231 (.A1(n19142), .A2(n27560), .ZN(N50103));
    NOR2X1 U37232 (.A1(n23071), .A2(n25904), .ZN(N50104));
    NOR2X1 U37233 (.A1(N2718), .A2(n13802), .ZN(N50105));
    NANDX1 U37234 (.A1(N1749), .A2(n43209), .ZN(N50106));
    NOR2X1 U37235 (.A1(n14410), .A2(n27210), .ZN(n50107));
    INVX1 U37236 (.I(n30173), .ZN(N50108));
    NOR2X1 U37237 (.A1(n31713), .A2(N6655), .ZN(N50109));
    NANDX1 U37238 (.A1(N6888), .A2(n42744), .ZN(N50110));
    NANDX1 U37239 (.A1(n27683), .A2(n33322), .ZN(N50111));
    NOR2X1 U37240 (.A1(N5669), .A2(n29905), .ZN(n50112));
    NOR2X1 U37241 (.A1(n19075), .A2(N4450), .ZN(N50113));
    NANDX1 U37242 (.A1(n36314), .A2(n35182), .ZN(n50114));
    NANDX1 U37243 (.A1(N8425), .A2(n31602), .ZN(N50115));
    NOR2X1 U37244 (.A1(n22227), .A2(n18770), .ZN(N50116));
    INVX1 U37245 (.I(N11643), .ZN(N50117));
    INVX1 U37246 (.I(N10555), .ZN(n50118));
    NANDX1 U37247 (.A1(N1330), .A2(n30408), .ZN(N50119));
    NANDX1 U37248 (.A1(n22722), .A2(n37062), .ZN(N50120));
    INVX1 U37249 (.I(n29609), .ZN(N50121));
    NOR2X1 U37250 (.A1(n33716), .A2(N3499), .ZN(N50122));
    INVX1 U37251 (.I(N3424), .ZN(N50123));
    NOR2X1 U37252 (.A1(n25127), .A2(n17005), .ZN(N50124));
    NOR2X1 U37253 (.A1(n29577), .A2(n39408), .ZN(N50125));
    INVX1 U37254 (.I(n21286), .ZN(N50126));
    NOR2X1 U37255 (.A1(N8868), .A2(n42568), .ZN(n50127));
    NOR2X1 U37256 (.A1(n20774), .A2(N7545), .ZN(n50128));
    INVX1 U37257 (.I(n32417), .ZN(N50129));
    NANDX1 U37258 (.A1(N11546), .A2(n17476), .ZN(N50130));
    NANDX1 U37259 (.A1(n31633), .A2(n42633), .ZN(N50131));
    NOR2X1 U37260 (.A1(n14902), .A2(N1732), .ZN(N50132));
    NANDX1 U37261 (.A1(n30594), .A2(n35447), .ZN(N50133));
    NOR2X1 U37262 (.A1(n36136), .A2(n28551), .ZN(N50134));
    NANDX1 U37263 (.A1(n17791), .A2(n35235), .ZN(N50135));
    NANDX1 U37264 (.A1(n37047), .A2(n20850), .ZN(N50136));
    NANDX1 U37265 (.A1(N4540), .A2(n41618), .ZN(N50137));
    NANDX1 U37266 (.A1(N3635), .A2(n13311), .ZN(N50138));
    INVX1 U37267 (.I(N860), .ZN(N50139));
    INVX1 U37268 (.I(n29924), .ZN(N50140));
    NOR2X1 U37269 (.A1(n25846), .A2(N3928), .ZN(n50141));
    NANDX1 U37270 (.A1(n14006), .A2(n36240), .ZN(N50142));
    INVX1 U37271 (.I(n28907), .ZN(N50143));
    INVX1 U37272 (.I(n38560), .ZN(N50144));
    NANDX1 U37273 (.A1(n19625), .A2(n43007), .ZN(N50145));
    NANDX1 U37274 (.A1(N4703), .A2(n13149), .ZN(N50146));
    NANDX1 U37275 (.A1(n29618), .A2(n24044), .ZN(N50147));
    NANDX1 U37276 (.A1(N6995), .A2(N2231), .ZN(N50148));
    NOR2X1 U37277 (.A1(N5140), .A2(n22437), .ZN(N50149));
    NOR2X1 U37278 (.A1(n18450), .A2(n19944), .ZN(N50150));
    INVX1 U37279 (.I(n32751), .ZN(N50151));
    INVX1 U37280 (.I(N10389), .ZN(N50152));
    NOR2X1 U37281 (.A1(n33155), .A2(N2228), .ZN(N50153));
    INVX1 U37282 (.I(n25922), .ZN(N50154));
    INVX1 U37283 (.I(n37396), .ZN(n50155));
    NANDX1 U37284 (.A1(N3965), .A2(n43104), .ZN(n50156));
    NOR2X1 U37285 (.A1(N3499), .A2(n31156), .ZN(N50157));
    NOR2X1 U37286 (.A1(N6327), .A2(n36997), .ZN(N50158));
    INVX1 U37287 (.I(n30371), .ZN(N50159));
    NOR2X1 U37288 (.A1(n17246), .A2(n22281), .ZN(N50160));
    NOR2X1 U37289 (.A1(N12066), .A2(N1245), .ZN(N50161));
    NOR2X1 U37290 (.A1(n20195), .A2(N10868), .ZN(N50162));
    NANDX1 U37291 (.A1(N9473), .A2(n40095), .ZN(N50163));
    NANDX1 U37292 (.A1(n14277), .A2(n29777), .ZN(N50164));
    INVX1 U37293 (.I(n22766), .ZN(N50165));
    INVX1 U37294 (.I(n15979), .ZN(N50166));
    NANDX1 U37295 (.A1(N12005), .A2(n19943), .ZN(N50167));
    NANDX1 U37296 (.A1(n41729), .A2(n13122), .ZN(N50168));
    NOR2X1 U37297 (.A1(n32683), .A2(n19448), .ZN(N50169));
    NANDX1 U37298 (.A1(n42934), .A2(n39498), .ZN(N50170));
    NANDX1 U37299 (.A1(N6387), .A2(n18306), .ZN(N50171));
    INVX1 U37300 (.I(n18452), .ZN(N50172));
    NOR2X1 U37301 (.A1(n19064), .A2(n38647), .ZN(N50173));
    NOR2X1 U37302 (.A1(n13549), .A2(n37799), .ZN(N50174));
    NANDX1 U37303 (.A1(n18422), .A2(n41755), .ZN(N50175));
    NANDX1 U37304 (.A1(n15203), .A2(n21048), .ZN(n50176));
    NANDX1 U37305 (.A1(n31181), .A2(n27417), .ZN(N50177));
    NANDX1 U37306 (.A1(n40803), .A2(n33417), .ZN(n50178));
    NANDX1 U37307 (.A1(N132), .A2(n27100), .ZN(N50179));
    NANDX1 U37308 (.A1(N9260), .A2(N3987), .ZN(N50180));
    NANDX1 U37309 (.A1(N5285), .A2(N6967), .ZN(N50181));
    INVX1 U37310 (.I(n13271), .ZN(N50182));
    NOR2X1 U37311 (.A1(n30892), .A2(N12180), .ZN(N50183));
    INVX1 U37312 (.I(n15746), .ZN(n50184));
    INVX1 U37313 (.I(n41644), .ZN(N50185));
    INVX1 U37314 (.I(n18037), .ZN(N50186));
    NANDX1 U37315 (.A1(n41507), .A2(N421), .ZN(N50187));
    INVX1 U37316 (.I(N8762), .ZN(N50188));
    INVX1 U37317 (.I(N9184), .ZN(N50189));
    INVX1 U37318 (.I(n14156), .ZN(N50190));
    NANDX1 U37319 (.A1(n26122), .A2(n41858), .ZN(N50191));
    NANDX1 U37320 (.A1(n42901), .A2(n15298), .ZN(N50192));
    NOR2X1 U37321 (.A1(n36568), .A2(n21351), .ZN(N50193));
    NOR2X1 U37322 (.A1(n33214), .A2(n33791), .ZN(N50194));
    INVX1 U37323 (.I(N9094), .ZN(N50195));
    INVX1 U37324 (.I(n15679), .ZN(N50196));
    INVX1 U37325 (.I(n26635), .ZN(N50197));
    INVX1 U37326 (.I(n35361), .ZN(n50198));
    NANDX1 U37327 (.A1(N1879), .A2(n41634), .ZN(n50199));
    NANDX1 U37328 (.A1(n35451), .A2(n19637), .ZN(N50200));
    NOR2X1 U37329 (.A1(N9841), .A2(n28820), .ZN(N50201));
    NOR2X1 U37330 (.A1(n13676), .A2(n25014), .ZN(n50202));
    NOR2X1 U37331 (.A1(N12062), .A2(N11019), .ZN(N50203));
    NANDX1 U37332 (.A1(n17039), .A2(n16603), .ZN(N50204));
    NANDX1 U37333 (.A1(n38390), .A2(N6831), .ZN(N50205));
    INVX1 U37334 (.I(n28708), .ZN(N50206));
    NANDX1 U37335 (.A1(N12407), .A2(n39597), .ZN(n50207));
    NANDX1 U37336 (.A1(n39276), .A2(N12439), .ZN(N50208));
    NOR2X1 U37337 (.A1(n20844), .A2(n38824), .ZN(N50209));
    NANDX1 U37338 (.A1(n19006), .A2(n42604), .ZN(N50210));
    NANDX1 U37339 (.A1(n38642), .A2(n21993), .ZN(N50211));
    INVX1 U37340 (.I(n13670), .ZN(N50212));
    NOR2X1 U37341 (.A1(n16903), .A2(n28363), .ZN(N50213));
    NOR2X1 U37342 (.A1(n28964), .A2(n39381), .ZN(N50214));
    NOR2X1 U37343 (.A1(N2530), .A2(N2191), .ZN(N50215));
    INVX1 U37344 (.I(n30599), .ZN(N50216));
    NANDX1 U37345 (.A1(n19344), .A2(N5514), .ZN(N50217));
    INVX1 U37346 (.I(n21430), .ZN(N50218));
    INVX1 U37347 (.I(n35037), .ZN(n50219));
    NANDX1 U37348 (.A1(n14076), .A2(N1415), .ZN(N50220));
    NANDX1 U37349 (.A1(n42580), .A2(N2823), .ZN(N50221));
    INVX1 U37350 (.I(n41711), .ZN(N50222));
    NANDX1 U37351 (.A1(n31611), .A2(N9911), .ZN(N50223));
    NOR2X1 U37352 (.A1(N1808), .A2(N3997), .ZN(N50224));
    NANDX1 U37353 (.A1(n19850), .A2(N8812), .ZN(N50225));
    INVX1 U37354 (.I(n15758), .ZN(N50226));
    NANDX1 U37355 (.A1(n37510), .A2(N7628), .ZN(N50227));
    NOR2X1 U37356 (.A1(n14317), .A2(N6328), .ZN(n50228));
    NOR2X1 U37357 (.A1(n19830), .A2(n15358), .ZN(N50229));
    NOR2X1 U37358 (.A1(N11148), .A2(N6922), .ZN(N50230));
    NANDX1 U37359 (.A1(n25223), .A2(n41488), .ZN(N50231));
    INVX1 U37360 (.I(n14010), .ZN(N50232));
    INVX1 U37361 (.I(n21277), .ZN(n50233));
    NANDX1 U37362 (.A1(N7367), .A2(n42567), .ZN(N50234));
    INVX1 U37363 (.I(N6802), .ZN(N50235));
    NOR2X1 U37364 (.A1(N5515), .A2(n23139), .ZN(N50236));
    INVX1 U37365 (.I(n14326), .ZN(N50237));
    NANDX1 U37366 (.A1(n15868), .A2(N4956), .ZN(N50238));
    NOR2X1 U37367 (.A1(n23495), .A2(N11616), .ZN(N50239));
    NOR2X1 U37368 (.A1(n19503), .A2(n27300), .ZN(N50240));
    NOR2X1 U37369 (.A1(n34860), .A2(N10620), .ZN(N50241));
    INVX1 U37370 (.I(n31461), .ZN(N50242));
    NOR2X1 U37371 (.A1(n15087), .A2(n29477), .ZN(N50243));
    INVX1 U37372 (.I(n18777), .ZN(N50244));
    INVX1 U37373 (.I(n40117), .ZN(n50245));
    NANDX1 U37374 (.A1(n17040), .A2(n39212), .ZN(N50246));
    INVX1 U37375 (.I(n23841), .ZN(N50247));
    NOR2X1 U37376 (.A1(n27736), .A2(n36659), .ZN(N50248));
    NANDX1 U37377 (.A1(n31741), .A2(n40985), .ZN(N50249));
    NOR2X1 U37378 (.A1(n26376), .A2(n39349), .ZN(N50250));
    NOR2X1 U37379 (.A1(n37991), .A2(N8556), .ZN(N50251));
    NANDX1 U37380 (.A1(N11498), .A2(n30745), .ZN(N50252));
    NANDX1 U37381 (.A1(n22118), .A2(n30929), .ZN(N50253));
    INVX1 U37382 (.I(n33290), .ZN(N50254));
    NOR2X1 U37383 (.A1(N12867), .A2(N8658), .ZN(N50255));
    NOR2X1 U37384 (.A1(n32861), .A2(N5302), .ZN(N50256));
    NANDX1 U37385 (.A1(N6428), .A2(N1041), .ZN(n50257));
    NANDX1 U37386 (.A1(n19949), .A2(n20514), .ZN(N50258));
    NOR2X1 U37387 (.A1(n13135), .A2(N6945), .ZN(N50259));
    INVX1 U37388 (.I(N328), .ZN(N50260));
    NOR2X1 U37389 (.A1(n21870), .A2(n39676), .ZN(n50261));
    NANDX1 U37390 (.A1(N6069), .A2(N4759), .ZN(N50262));
    INVX1 U37391 (.I(n17566), .ZN(N50263));
    NOR2X1 U37392 (.A1(N11621), .A2(n39683), .ZN(N50264));
    NANDX1 U37393 (.A1(n38484), .A2(n19180), .ZN(N50265));
    INVX1 U37394 (.I(N7878), .ZN(N50266));
    INVX1 U37395 (.I(N5542), .ZN(N50267));
    NANDX1 U37396 (.A1(n33139), .A2(n26925), .ZN(N50268));
    NANDX1 U37397 (.A1(n23859), .A2(n16736), .ZN(n50269));
    INVX1 U37398 (.I(N900), .ZN(N50270));
    NANDX1 U37399 (.A1(n16136), .A2(n40996), .ZN(n50271));
    NANDX1 U37400 (.A1(n16463), .A2(n39919), .ZN(N50272));
    NOR2X1 U37401 (.A1(N2346), .A2(N10842), .ZN(N50273));
    NOR2X1 U37402 (.A1(n40257), .A2(N6421), .ZN(N50274));
    NOR2X1 U37403 (.A1(n21968), .A2(N7721), .ZN(n50275));
    NOR2X1 U37404 (.A1(n34607), .A2(N2732), .ZN(N50276));
    NANDX1 U37405 (.A1(n29150), .A2(N290), .ZN(N50277));
    NOR2X1 U37406 (.A1(n34691), .A2(n30707), .ZN(N50278));
    INVX1 U37407 (.I(N7823), .ZN(N50279));
    INVX1 U37408 (.I(n14127), .ZN(N50280));
    NANDX1 U37409 (.A1(n27081), .A2(n15027), .ZN(N50281));
    NOR2X1 U37410 (.A1(n32897), .A2(N12550), .ZN(N50282));
    NANDX1 U37411 (.A1(n39039), .A2(n42148), .ZN(N50283));
    NANDX1 U37412 (.A1(n41385), .A2(N9518), .ZN(N50284));
    INVX1 U37413 (.I(n38169), .ZN(N50285));
    NANDX1 U37414 (.A1(n37449), .A2(n16664), .ZN(N50286));
    INVX1 U37415 (.I(N1355), .ZN(N50287));
    NANDX1 U37416 (.A1(n38902), .A2(n27912), .ZN(N50288));
    NANDX1 U37417 (.A1(n39191), .A2(n28514), .ZN(N50289));
    NANDX1 U37418 (.A1(n16105), .A2(n29102), .ZN(N50290));
    NANDX1 U37419 (.A1(n40185), .A2(n43229), .ZN(N50291));
    NOR2X1 U37420 (.A1(n13473), .A2(N4463), .ZN(N50292));
    NOR2X1 U37421 (.A1(N2897), .A2(N6692), .ZN(N50293));
    NOR2X1 U37422 (.A1(n31616), .A2(N5368), .ZN(N50294));
    INVX1 U37423 (.I(n29528), .ZN(N50295));
    NOR2X1 U37424 (.A1(N10514), .A2(n13904), .ZN(N50296));
    NANDX1 U37425 (.A1(n37642), .A2(n20247), .ZN(N50297));
    NOR2X1 U37426 (.A1(n38996), .A2(n17724), .ZN(N50298));
    NOR2X1 U37427 (.A1(n13115), .A2(n23711), .ZN(N50299));
    INVX1 U37428 (.I(n41629), .ZN(N50300));
    NOR2X1 U37429 (.A1(n32963), .A2(n16938), .ZN(N50301));
    INVX1 U37430 (.I(n19355), .ZN(N50302));
    NANDX1 U37431 (.A1(N12057), .A2(n32827), .ZN(N50303));
    INVX1 U37432 (.I(n36370), .ZN(N50304));
    NOR2X1 U37433 (.A1(N7208), .A2(N8564), .ZN(N50305));
    NOR2X1 U37434 (.A1(N2255), .A2(n36269), .ZN(N50306));
    NOR2X1 U37435 (.A1(n39971), .A2(n36462), .ZN(N50307));
    INVX1 U37436 (.I(n39832), .ZN(N50308));
    NOR2X1 U37437 (.A1(n13111), .A2(n32390), .ZN(N50309));
    NANDX1 U37438 (.A1(n20514), .A2(N10058), .ZN(N50310));
    NANDX1 U37439 (.A1(N752), .A2(n16595), .ZN(n50311));
    NANDX1 U37440 (.A1(n21667), .A2(n39237), .ZN(N50312));
    INVX1 U37441 (.I(N4138), .ZN(N50313));
    INVX1 U37442 (.I(n29775), .ZN(n50314));
    NOR2X1 U37443 (.A1(n37626), .A2(n30291), .ZN(N50315));
    NOR2X1 U37444 (.A1(n19557), .A2(n27178), .ZN(N50316));
    INVX1 U37445 (.I(n33103), .ZN(N50317));
    NANDX1 U37446 (.A1(n22963), .A2(n22384), .ZN(N50318));
    INVX1 U37447 (.I(n15952), .ZN(N50319));
    INVX1 U37448 (.I(N11969), .ZN(N50320));
    NOR2X1 U37449 (.A1(n28358), .A2(n34038), .ZN(N50321));
    INVX1 U37450 (.I(N5399), .ZN(n50322));
    NANDX1 U37451 (.A1(n37570), .A2(N6151), .ZN(N50323));
    NANDX1 U37452 (.A1(N10882), .A2(n27817), .ZN(N50324));
    NANDX1 U37453 (.A1(n34283), .A2(n21634), .ZN(N50325));
    NOR2X1 U37454 (.A1(n20585), .A2(n27507), .ZN(N50326));
    NANDX1 U37455 (.A1(n40555), .A2(n15958), .ZN(N50327));
    NOR2X1 U37456 (.A1(n24260), .A2(N2652), .ZN(N50328));
    INVX1 U37457 (.I(n43371), .ZN(N50329));
    NOR2X1 U37458 (.A1(n22863), .A2(n15508), .ZN(N50330));
    INVX1 U37459 (.I(n38110), .ZN(N50331));
    NOR2X1 U37460 (.A1(n34354), .A2(N12675), .ZN(N50332));
    NANDX1 U37461 (.A1(n42976), .A2(N7753), .ZN(N50333));
    NOR2X1 U37462 (.A1(n37073), .A2(n13903), .ZN(N50334));
    NANDX1 U37463 (.A1(n37634), .A2(n31400), .ZN(N50335));
    INVX1 U37464 (.I(n28444), .ZN(N50336));
    NOR2X1 U37465 (.A1(n35683), .A2(n38709), .ZN(N50337));
    NANDX1 U37466 (.A1(n37296), .A2(n25471), .ZN(N50338));
    NANDX1 U37467 (.A1(n14993), .A2(N6259), .ZN(N50339));
    NANDX1 U37468 (.A1(n15472), .A2(n39309), .ZN(N50340));
    NANDX1 U37469 (.A1(n38334), .A2(N11345), .ZN(N50341));
    NANDX1 U37470 (.A1(n22651), .A2(n38820), .ZN(N50342));
    NANDX1 U37471 (.A1(n35325), .A2(n13389), .ZN(N50343));
    NOR2X1 U37472 (.A1(n43077), .A2(n21733), .ZN(N50344));
    NOR2X1 U37473 (.A1(N3188), .A2(n36973), .ZN(N50345));
    NANDX1 U37474 (.A1(n24267), .A2(N1083), .ZN(N50346));
    NOR2X1 U37475 (.A1(n23507), .A2(n26445), .ZN(N50347));
    INVX1 U37476 (.I(n39934), .ZN(n50348));
    INVX1 U37477 (.I(n13797), .ZN(N50349));
    NOR2X1 U37478 (.A1(n24940), .A2(N9735), .ZN(N50350));
    NANDX1 U37479 (.A1(n40411), .A2(N5571), .ZN(N50351));
    NOR2X1 U37480 (.A1(n35272), .A2(N6595), .ZN(N50352));
    NANDX1 U37481 (.A1(n14450), .A2(N1943), .ZN(N50353));
    INVX1 U37482 (.I(n39454), .ZN(N50354));
    INVX1 U37483 (.I(n17438), .ZN(N50355));
    NOR2X1 U37484 (.A1(n16423), .A2(N8563), .ZN(N50356));
    INVX1 U37485 (.I(n43076), .ZN(N50357));
    INVX1 U37486 (.I(N2400), .ZN(N50358));
    INVX1 U37487 (.I(n30410), .ZN(N50359));
    INVX1 U37488 (.I(n27131), .ZN(N50360));
    NANDX1 U37489 (.A1(N12048), .A2(n37078), .ZN(N50361));
    NOR2X1 U37490 (.A1(n30573), .A2(n18546), .ZN(N50362));
    INVX1 U37491 (.I(n30342), .ZN(N50363));
    NOR2X1 U37492 (.A1(n37516), .A2(n36966), .ZN(N50364));
    NANDX1 U37493 (.A1(N639), .A2(n38219), .ZN(n50365));
    NOR2X1 U37494 (.A1(n35733), .A2(N4340), .ZN(N50366));
    NOR2X1 U37495 (.A1(n40743), .A2(N11458), .ZN(N50367));
    NOR2X1 U37496 (.A1(N3374), .A2(n20020), .ZN(N50368));
    NOR2X1 U37497 (.A1(N2977), .A2(N3548), .ZN(N50369));
    NOR2X1 U37498 (.A1(n36814), .A2(n33957), .ZN(N50370));
    INVX1 U37499 (.I(n20472), .ZN(N50371));
    NANDX1 U37500 (.A1(N3017), .A2(N3758), .ZN(N50372));
    INVX1 U37501 (.I(n23270), .ZN(N50373));
    NOR2X1 U37502 (.A1(n19904), .A2(N10139), .ZN(N50374));
    NOR2X1 U37503 (.A1(n13948), .A2(N3632), .ZN(N50375));
    INVX1 U37504 (.I(N4266), .ZN(N50376));
    NANDX1 U37505 (.A1(n25522), .A2(n39998), .ZN(N50377));
    NANDX1 U37506 (.A1(N12276), .A2(n37268), .ZN(N50378));
    INVX1 U37507 (.I(n27768), .ZN(N50379));
    NANDX1 U37508 (.A1(N3234), .A2(n21393), .ZN(N50380));
    NANDX1 U37509 (.A1(N6781), .A2(N7097), .ZN(N50381));
    NANDX1 U37510 (.A1(n30417), .A2(N8386), .ZN(N50382));
    NOR2X1 U37511 (.A1(n29317), .A2(N1083), .ZN(N50383));
    INVX1 U37512 (.I(N6955), .ZN(N50384));
    NANDX1 U37513 (.A1(N9057), .A2(n26859), .ZN(N50385));
    NANDX1 U37514 (.A1(n36523), .A2(n30486), .ZN(N50386));
    INVX1 U37515 (.I(N7159), .ZN(N50387));
    NOR2X1 U37516 (.A1(n26179), .A2(n32680), .ZN(N50388));
    NANDX1 U37517 (.A1(n41408), .A2(N1483), .ZN(N50389));
    INVX1 U37518 (.I(n34942), .ZN(N50390));
    NANDX1 U37519 (.A1(N1600), .A2(n27855), .ZN(N50391));
    NOR2X1 U37520 (.A1(n24576), .A2(n34635), .ZN(N50392));
    NANDX1 U37521 (.A1(n40894), .A2(N11259), .ZN(N50393));
    INVX1 U37522 (.I(n23892), .ZN(n50394));
    NOR2X1 U37523 (.A1(N3094), .A2(N10646), .ZN(n50395));
    NANDX1 U37524 (.A1(n27445), .A2(n19703), .ZN(N50396));
    NOR2X1 U37525 (.A1(N8142), .A2(N2433), .ZN(N50397));
    NOR2X1 U37526 (.A1(n35942), .A2(N9591), .ZN(N50398));
    NANDX1 U37527 (.A1(n18648), .A2(n31951), .ZN(N50399));
    INVX1 U37528 (.I(N6263), .ZN(N50400));
    INVX1 U37529 (.I(n13952), .ZN(N50401));
    INVX1 U37530 (.I(n42043), .ZN(N50402));
    INVX1 U37531 (.I(n15266), .ZN(N50403));
    NOR2X1 U37532 (.A1(n29807), .A2(n39580), .ZN(N50404));
    NANDX1 U37533 (.A1(n16908), .A2(N7367), .ZN(N50405));
    NOR2X1 U37534 (.A1(n40799), .A2(n27301), .ZN(N50406));
    INVX1 U37535 (.I(n41125), .ZN(N50407));
    INVX1 U37536 (.I(n23786), .ZN(N50408));
    NANDX1 U37537 (.A1(n20993), .A2(n31927), .ZN(N50409));
    NOR2X1 U37538 (.A1(N7961), .A2(n24396), .ZN(N50410));
    INVX1 U37539 (.I(n19359), .ZN(N50411));
    NOR2X1 U37540 (.A1(N7535), .A2(n18560), .ZN(N50412));
    NANDX1 U37541 (.A1(n30648), .A2(n22192), .ZN(N50413));
    INVX1 U37542 (.I(n18898), .ZN(N50414));
    NOR2X1 U37543 (.A1(n41663), .A2(N3997), .ZN(N50415));
    NOR2X1 U37544 (.A1(n37771), .A2(n26194), .ZN(N50416));
    INVX1 U37545 (.I(n34817), .ZN(N50417));
    NANDX1 U37546 (.A1(N7350), .A2(n18645), .ZN(N50418));
    NANDX1 U37547 (.A1(N5002), .A2(n29363), .ZN(N50419));
    INVX1 U37548 (.I(N12036), .ZN(N50420));
    INVX1 U37549 (.I(n15510), .ZN(N50421));
    NOR2X1 U37550 (.A1(n37676), .A2(n29586), .ZN(N50422));
    NANDX1 U37551 (.A1(n13562), .A2(n18837), .ZN(n50423));
    INVX1 U37552 (.I(n21802), .ZN(N50424));
    NANDX1 U37553 (.A1(n14628), .A2(N521), .ZN(N50425));
    NOR2X1 U37554 (.A1(n33525), .A2(n17622), .ZN(N50426));
    NOR2X1 U37555 (.A1(n37522), .A2(N10738), .ZN(N50427));
    NOR2X1 U37556 (.A1(N9923), .A2(n20761), .ZN(N50428));
    INVX1 U37557 (.I(N6533), .ZN(N50429));
    NOR2X1 U37558 (.A1(N12264), .A2(n42955), .ZN(N50430));
    NOR2X1 U37559 (.A1(n41626), .A2(n26539), .ZN(n50431));
    INVX1 U37560 (.I(n27869), .ZN(N50432));
    NOR2X1 U37561 (.A1(n25369), .A2(n22072), .ZN(N50433));
    INVX1 U37562 (.I(N12135), .ZN(N50434));
    INVX1 U37563 (.I(n26357), .ZN(N50435));
    NOR2X1 U37564 (.A1(n36794), .A2(n30387), .ZN(N50436));
    INVX1 U37565 (.I(n37314), .ZN(N50437));
    INVX1 U37566 (.I(n23627), .ZN(N50438));
    NANDX1 U37567 (.A1(n35638), .A2(n17676), .ZN(N50439));
    INVX1 U37568 (.I(N4761), .ZN(N50440));
    NANDX1 U37569 (.A1(n22321), .A2(n41852), .ZN(N50441));
    NANDX1 U37570 (.A1(n40110), .A2(N10644), .ZN(N50442));
    NOR2X1 U37571 (.A1(n42261), .A2(n41949), .ZN(N50443));
    NOR2X1 U37572 (.A1(n12976), .A2(n26345), .ZN(N50444));
    INVX1 U37573 (.I(n38344), .ZN(N50445));
    NANDX1 U37574 (.A1(n14647), .A2(N7006), .ZN(N50446));
    INVX1 U37575 (.I(n41004), .ZN(N50447));
    INVX1 U37576 (.I(N2938), .ZN(N50448));
    NANDX1 U37577 (.A1(n36694), .A2(n29932), .ZN(N50449));
    NANDX1 U37578 (.A1(n16849), .A2(n31075), .ZN(N50450));
    INVX1 U37579 (.I(n24204), .ZN(N50451));
    NOR2X1 U37580 (.A1(n31864), .A2(n41482), .ZN(N50452));
    NOR2X1 U37581 (.A1(n30244), .A2(N1180), .ZN(N50453));
    NOR2X1 U37582 (.A1(n30567), .A2(n14153), .ZN(N50454));
    INVX1 U37583 (.I(n29043), .ZN(n50455));
    NOR2X1 U37584 (.A1(n42716), .A2(N1596), .ZN(N50456));
    INVX1 U37585 (.I(n37587), .ZN(N50457));
    NOR2X1 U37586 (.A1(N11324), .A2(n34272), .ZN(N50458));
    INVX1 U37587 (.I(N8855), .ZN(N50459));
    NOR2X1 U37588 (.A1(n41925), .A2(n36772), .ZN(n50460));
    NANDX1 U37589 (.A1(n28384), .A2(n28237), .ZN(N50461));
    NOR2X1 U37590 (.A1(n15986), .A2(N11868), .ZN(N50462));
    NOR2X1 U37591 (.A1(n38300), .A2(n33412), .ZN(N50463));
    NOR2X1 U37592 (.A1(n39462), .A2(N9863), .ZN(N50464));
    NOR2X1 U37593 (.A1(n26941), .A2(n40429), .ZN(N50465));
    INVX1 U37594 (.I(n13209), .ZN(N50466));
    NANDX1 U37595 (.A1(n22956), .A2(N12452), .ZN(N50467));
    INVX1 U37596 (.I(n19632), .ZN(N50468));
    NANDX1 U37597 (.A1(N3173), .A2(n30955), .ZN(N50469));
    INVX1 U37598 (.I(n42159), .ZN(N50470));
    NOR2X1 U37599 (.A1(N3796), .A2(n40611), .ZN(N50471));
    INVX1 U37600 (.I(N3448), .ZN(N50472));
    INVX1 U37601 (.I(n40705), .ZN(N50473));
    NOR2X1 U37602 (.A1(n31187), .A2(N9100), .ZN(N50474));
    NOR2X1 U37603 (.A1(n26014), .A2(n32191), .ZN(N50475));
    NANDX1 U37604 (.A1(N11683), .A2(n42053), .ZN(N50476));
    NOR2X1 U37605 (.A1(n38624), .A2(n28689), .ZN(N50477));
    INVX1 U37606 (.I(N8360), .ZN(N50478));
    INVX1 U37607 (.I(n13600), .ZN(N50479));
    NOR2X1 U37608 (.A1(n18169), .A2(n22912), .ZN(N50480));
    INVX1 U37609 (.I(n21341), .ZN(N50481));
    NANDX1 U37610 (.A1(n26934), .A2(n20028), .ZN(N50482));
    NOR2X1 U37611 (.A1(n30729), .A2(N6846), .ZN(N50483));
    INVX1 U37612 (.I(n34176), .ZN(N50484));
    NANDX1 U37613 (.A1(N6110), .A2(N331), .ZN(N50485));
    NOR2X1 U37614 (.A1(N4890), .A2(N7189), .ZN(N50486));
    INVX1 U37615 (.I(n37080), .ZN(N50487));
    NOR2X1 U37616 (.A1(n37138), .A2(n25341), .ZN(N50488));
    NANDX1 U37617 (.A1(n21969), .A2(N10557), .ZN(N50489));
    NOR2X1 U37618 (.A1(n30329), .A2(N11452), .ZN(N50490));
    NANDX1 U37619 (.A1(n40820), .A2(n19301), .ZN(N50491));
    INVX1 U37620 (.I(n37236), .ZN(N50492));
    NOR2X1 U37621 (.A1(N6269), .A2(n20697), .ZN(N50493));
    INVX1 U37622 (.I(N2679), .ZN(N50494));
    NANDX1 U37623 (.A1(n13722), .A2(N1237), .ZN(N50495));
    NOR2X1 U37624 (.A1(N2617), .A2(N7346), .ZN(N50496));
    NOR2X1 U37625 (.A1(N2058), .A2(N1915), .ZN(N50497));
    INVX1 U37626 (.I(n27513), .ZN(N50498));
    NOR2X1 U37627 (.A1(N7335), .A2(N10859), .ZN(N50499));
    NANDX1 U37628 (.A1(n40167), .A2(n32827), .ZN(N50500));
    NANDX1 U37629 (.A1(n20171), .A2(n19683), .ZN(N50501));
    NANDX1 U37630 (.A1(N3455), .A2(N6710), .ZN(N50502));
    INVX1 U37631 (.I(N9650), .ZN(N50503));
    NANDX1 U37632 (.A1(n28379), .A2(n15919), .ZN(N50504));
    NANDX1 U37633 (.A1(n35255), .A2(N8277), .ZN(n50505));
    NANDX1 U37634 (.A1(N5504), .A2(N9513), .ZN(N50506));
    NANDX1 U37635 (.A1(n41272), .A2(n16859), .ZN(N50507));
    NANDX1 U37636 (.A1(n43329), .A2(N8453), .ZN(N50508));
    NANDX1 U37637 (.A1(n17050), .A2(n37127), .ZN(N50509));
    NANDX1 U37638 (.A1(n27908), .A2(N4197), .ZN(N50510));
    NOR2X1 U37639 (.A1(n17262), .A2(N4656), .ZN(n50511));
    NOR2X1 U37640 (.A1(n36945), .A2(n16566), .ZN(N50512));
    INVX1 U37641 (.I(n33334), .ZN(N50513));
    NOR2X1 U37642 (.A1(n23024), .A2(n23487), .ZN(N50514));
    NANDX1 U37643 (.A1(n28622), .A2(n24017), .ZN(N50515));
    NOR2X1 U37644 (.A1(n36899), .A2(n22179), .ZN(N50516));
    INVX1 U37645 (.I(N2939), .ZN(N50517));
    INVX1 U37646 (.I(N7126), .ZN(N50518));
    INVX1 U37647 (.I(N8863), .ZN(N50519));
    NANDX1 U37648 (.A1(N7610), .A2(N4904), .ZN(N50520));
    NOR2X1 U37649 (.A1(N1264), .A2(N8279), .ZN(N50521));
    INVX1 U37650 (.I(n38613), .ZN(N50522));
    NANDX1 U37651 (.A1(n15408), .A2(n43268), .ZN(N50523));
    NOR2X1 U37652 (.A1(n42032), .A2(n16361), .ZN(N50524));
    NOR2X1 U37653 (.A1(n31894), .A2(N10344), .ZN(N50525));
    NOR2X1 U37654 (.A1(N1588), .A2(n43025), .ZN(N50526));
    NOR2X1 U37655 (.A1(n25604), .A2(N3377), .ZN(N50527));
    INVX1 U37656 (.I(n37462), .ZN(N50528));
    NOR2X1 U37657 (.A1(n15539), .A2(n25498), .ZN(N50529));
    NOR2X1 U37658 (.A1(n14696), .A2(n24040), .ZN(N50530));
    INVX1 U37659 (.I(n22305), .ZN(N50531));
    INVX1 U37660 (.I(n30202), .ZN(N50532));
    NOR2X1 U37661 (.A1(n26902), .A2(n28348), .ZN(N50533));
    INVX1 U37662 (.I(n24930), .ZN(n50534));
    INVX1 U37663 (.I(N8183), .ZN(N50535));
    NOR2X1 U37664 (.A1(n31995), .A2(n14223), .ZN(N50536));
    NANDX1 U37665 (.A1(N10096), .A2(n24566), .ZN(N50537));
    INVX1 U37666 (.I(N11683), .ZN(N50538));
    NANDX1 U37667 (.A1(N7940), .A2(n37287), .ZN(N50539));
    NOR2X1 U37668 (.A1(n30860), .A2(n31276), .ZN(N50540));
    NANDX1 U37669 (.A1(n36079), .A2(N2981), .ZN(N50541));
    NANDX1 U37670 (.A1(N7302), .A2(n16701), .ZN(N50542));
    NANDX1 U37671 (.A1(n19286), .A2(N2172), .ZN(N50543));
    NANDX1 U37672 (.A1(n32533), .A2(n18753), .ZN(N50544));
    NANDX1 U37673 (.A1(n40921), .A2(N210), .ZN(N50545));
    NOR2X1 U37674 (.A1(n38783), .A2(n43406), .ZN(N50546));
    INVX1 U37675 (.I(N9534), .ZN(N50547));
    NOR2X1 U37676 (.A1(n28571), .A2(n23779), .ZN(N50548));
    NANDX1 U37677 (.A1(n29933), .A2(n27257), .ZN(N50549));
    NANDX1 U37678 (.A1(n13427), .A2(n34111), .ZN(N50550));
    INVX1 U37679 (.I(n34383), .ZN(N50551));
    NOR2X1 U37680 (.A1(n20510), .A2(n27043), .ZN(N50552));
    INVX1 U37681 (.I(n17491), .ZN(N50553));
    NOR2X1 U37682 (.A1(N8191), .A2(n36776), .ZN(N50554));
    NOR2X1 U37683 (.A1(n30154), .A2(n25836), .ZN(N50555));
    NANDX1 U37684 (.A1(n36993), .A2(n12964), .ZN(N50556));
    INVX1 U37685 (.I(n23474), .ZN(N50557));
    INVX1 U37686 (.I(N11018), .ZN(N50558));
    NOR2X1 U37687 (.A1(N7488), .A2(n21676), .ZN(N50559));
    NANDX1 U37688 (.A1(n20946), .A2(n21100), .ZN(N50560));
    INVX1 U37689 (.I(N4731), .ZN(N50561));
    NOR2X1 U37690 (.A1(N6294), .A2(n28521), .ZN(N50562));
    NOR2X1 U37691 (.A1(n30356), .A2(n38716), .ZN(N50563));
    NOR2X1 U37692 (.A1(n13926), .A2(n34504), .ZN(N50564));
    INVX1 U37693 (.I(n14197), .ZN(N50565));
    INVX1 U37694 (.I(n13237), .ZN(N50566));
    INVX1 U37695 (.I(n29375), .ZN(N50567));
    NANDX1 U37696 (.A1(n17192), .A2(N12575), .ZN(n50568));
    NOR2X1 U37697 (.A1(n28276), .A2(n25728), .ZN(N50569));
    NOR2X1 U37698 (.A1(n28973), .A2(n13884), .ZN(N50570));
    INVX1 U37699 (.I(N7176), .ZN(N50571));
    INVX1 U37700 (.I(n34950), .ZN(N50572));
    INVX1 U37701 (.I(N2837), .ZN(N50573));
    NOR2X1 U37702 (.A1(n36099), .A2(n42282), .ZN(N50574));
    NOR2X1 U37703 (.A1(n38673), .A2(n29165), .ZN(N50575));
    NANDX1 U37704 (.A1(N7964), .A2(n43090), .ZN(N50576));
    NANDX1 U37705 (.A1(n27897), .A2(N3494), .ZN(N50577));
    NOR2X1 U37706 (.A1(n41133), .A2(N9812), .ZN(N50578));
    INVX1 U37707 (.I(n26412), .ZN(N50579));
    NOR2X1 U37708 (.A1(N10893), .A2(n14335), .ZN(N50580));
    NOR2X1 U37709 (.A1(n26301), .A2(n20852), .ZN(N50581));
    NANDX1 U37710 (.A1(n40184), .A2(n24536), .ZN(N50582));
    NOR2X1 U37711 (.A1(N6682), .A2(N5694), .ZN(N50583));
    INVX1 U37712 (.I(N9518), .ZN(N50584));
    NOR2X1 U37713 (.A1(N4743), .A2(N8327), .ZN(N50585));
    NOR2X1 U37714 (.A1(n33095), .A2(n37491), .ZN(N50586));
    NANDX1 U37715 (.A1(n30738), .A2(n26788), .ZN(n50587));
    INVX1 U37716 (.I(n15162), .ZN(N50588));
    INVX1 U37717 (.I(n41251), .ZN(N50589));
    INVX1 U37718 (.I(n19453), .ZN(N50590));
    INVX1 U37719 (.I(n18593), .ZN(n50591));
    NOR2X1 U37720 (.A1(n40141), .A2(n32928), .ZN(N50592));
    INVX1 U37721 (.I(n22969), .ZN(N50593));
    NANDX1 U37722 (.A1(n14286), .A2(n19681), .ZN(n50594));
    NOR2X1 U37723 (.A1(n41599), .A2(n26362), .ZN(n50595));
    NOR2X1 U37724 (.A1(n43395), .A2(n35879), .ZN(N50596));
    NANDX1 U37725 (.A1(n37817), .A2(n33885), .ZN(n50597));
    NOR2X1 U37726 (.A1(n27439), .A2(n17583), .ZN(N50598));
    INVX1 U37727 (.I(n14704), .ZN(N50599));
    NANDX1 U37728 (.A1(n20659), .A2(n19545), .ZN(N50600));
    NANDX1 U37729 (.A1(N8117), .A2(n22046), .ZN(N50601));
    NANDX1 U37730 (.A1(N4213), .A2(n40639), .ZN(n50602));
    NOR2X1 U37731 (.A1(N882), .A2(n19774), .ZN(N50603));
    NOR2X1 U37732 (.A1(n23850), .A2(n19760), .ZN(N50604));
    NANDX1 U37733 (.A1(n33210), .A2(N810), .ZN(N50605));
    INVX1 U37734 (.I(N5779), .ZN(N50606));
    INVX1 U37735 (.I(n41648), .ZN(N50607));
    NOR2X1 U37736 (.A1(n42501), .A2(n35993), .ZN(N50608));
    NOR2X1 U37737 (.A1(N6173), .A2(N9639), .ZN(N50609));
    NOR2X1 U37738 (.A1(n41469), .A2(n14023), .ZN(N50610));
    NANDX1 U37739 (.A1(N8335), .A2(n33567), .ZN(N50611));
    INVX1 U37740 (.I(n16452), .ZN(N50612));
    NOR2X1 U37741 (.A1(N6326), .A2(N10344), .ZN(N50613));
    NOR2X1 U37742 (.A1(n18659), .A2(N905), .ZN(N50614));
    INVX1 U37743 (.I(N4500), .ZN(N50615));
    INVX1 U37744 (.I(n28199), .ZN(N50616));
    INVX1 U37745 (.I(N4172), .ZN(N50617));
    NANDX1 U37746 (.A1(N2879), .A2(N9951), .ZN(N50618));
    NOR2X1 U37747 (.A1(n34207), .A2(n30967), .ZN(N50619));
    NOR2X1 U37748 (.A1(n16407), .A2(N9244), .ZN(N50620));
    NOR2X1 U37749 (.A1(n26045), .A2(n38254), .ZN(N50621));
    NOR2X1 U37750 (.A1(n40067), .A2(n24690), .ZN(N50622));
    NOR2X1 U37751 (.A1(n19842), .A2(N1025), .ZN(N50623));
    INVX1 U37752 (.I(n21662), .ZN(N50624));
    NOR2X1 U37753 (.A1(n13606), .A2(n20648), .ZN(N50625));
    NOR2X1 U37754 (.A1(N4191), .A2(n18767), .ZN(n50626));
    NANDX1 U37755 (.A1(n18625), .A2(N3493), .ZN(N50627));
    NANDX1 U37756 (.A1(n22796), .A2(n22181), .ZN(N50628));
    NOR2X1 U37757 (.A1(n22426), .A2(n28422), .ZN(N50629));
    NANDX1 U37758 (.A1(N9921), .A2(n33690), .ZN(N50630));
    INVX1 U37759 (.I(N8844), .ZN(N50631));
    NOR2X1 U37760 (.A1(N7083), .A2(N3625), .ZN(N50632));
    NOR2X1 U37761 (.A1(n36830), .A2(n17995), .ZN(N50633));
    NANDX1 U37762 (.A1(n13199), .A2(n19019), .ZN(n50634));
    NOR2X1 U37763 (.A1(n34860), .A2(n26368), .ZN(N50635));
    NOR2X1 U37764 (.A1(N1715), .A2(n31735), .ZN(N50636));
    NANDX1 U37765 (.A1(n20481), .A2(N8449), .ZN(N50637));
    NANDX1 U37766 (.A1(n13653), .A2(n33260), .ZN(N50638));
    INVX1 U37767 (.I(n35834), .ZN(N50639));
    INVX1 U37768 (.I(n20889), .ZN(N50640));
    NOR2X1 U37769 (.A1(n15262), .A2(n20489), .ZN(N50641));
    NANDX1 U37770 (.A1(n39772), .A2(n29332), .ZN(N50642));
    INVX1 U37771 (.I(n36535), .ZN(N50643));
    NOR2X1 U37772 (.A1(n38457), .A2(n19572), .ZN(N50644));
    NOR2X1 U37773 (.A1(n38554), .A2(n22450), .ZN(N50645));
    NANDX1 U37774 (.A1(n41914), .A2(N3517), .ZN(N50646));
    INVX1 U37775 (.I(n15407), .ZN(n50647));
    NANDX1 U37776 (.A1(n20485), .A2(n26242), .ZN(N50648));
    NANDX1 U37777 (.A1(n28933), .A2(N12229), .ZN(N50649));
    NANDX1 U37778 (.A1(N8401), .A2(N10691), .ZN(N50650));
    NOR2X1 U37779 (.A1(n15558), .A2(n21259), .ZN(N50651));
    NANDX1 U37780 (.A1(n20500), .A2(n31427), .ZN(N50652));
    INVX1 U37781 (.I(N6479), .ZN(N50653));
    INVX1 U37782 (.I(N3923), .ZN(N50654));
    NOR2X1 U37783 (.A1(n29602), .A2(n42379), .ZN(N50655));
    NANDX1 U37784 (.A1(n26759), .A2(n37461), .ZN(N50656));
    NANDX1 U37785 (.A1(n42935), .A2(n35902), .ZN(N50657));
    NANDX1 U37786 (.A1(n21365), .A2(n40988), .ZN(N50658));
    INVX1 U37787 (.I(n41850), .ZN(N50659));
    INVX1 U37788 (.I(n34737), .ZN(N50660));
    INVX1 U37789 (.I(n15345), .ZN(N50661));
    NANDX1 U37790 (.A1(n15070), .A2(n26035), .ZN(N50662));
    INVX1 U37791 (.I(n20308), .ZN(N50663));
    NANDX1 U37792 (.A1(n42617), .A2(n40807), .ZN(N50664));
    NANDX1 U37793 (.A1(n21370), .A2(n36965), .ZN(N50665));
    INVX1 U37794 (.I(n25292), .ZN(n50666));
    NOR2X1 U37795 (.A1(n18023), .A2(n24199), .ZN(N50667));
    NANDX1 U37796 (.A1(N1309), .A2(N7867), .ZN(N50668));
    INVX1 U37797 (.I(n33923), .ZN(N50669));
    NANDX1 U37798 (.A1(n26542), .A2(N1496), .ZN(N50670));
    INVX1 U37799 (.I(N2417), .ZN(N50671));
    NOR2X1 U37800 (.A1(n34079), .A2(n26833), .ZN(N50672));
    INVX1 U37801 (.I(N5951), .ZN(N50673));
    NOR2X1 U37802 (.A1(N11292), .A2(n21665), .ZN(N50674));
    NANDX1 U37803 (.A1(n31599), .A2(n15166), .ZN(N50675));
    NANDX1 U37804 (.A1(n18613), .A2(n29774), .ZN(N50676));
    INVX1 U37805 (.I(N1785), .ZN(N50677));
    INVX1 U37806 (.I(n39583), .ZN(N50678));
    INVX1 U37807 (.I(n25897), .ZN(N50679));
    NANDX1 U37808 (.A1(n42307), .A2(n16885), .ZN(N50680));
    NANDX1 U37809 (.A1(N940), .A2(N7336), .ZN(N50681));
    NOR2X1 U37810 (.A1(n17161), .A2(N8831), .ZN(N50682));
    INVX1 U37811 (.I(N9257), .ZN(N50683));
    INVX1 U37812 (.I(n19078), .ZN(N50684));
    NANDX1 U37813 (.A1(n38076), .A2(n25028), .ZN(N50685));
    NANDX1 U37814 (.A1(N5895), .A2(N3221), .ZN(n50686));
    NOR2X1 U37815 (.A1(n27173), .A2(N8066), .ZN(N50687));
    NANDX1 U37816 (.A1(n35465), .A2(n37839), .ZN(N50688));
    NANDX1 U37817 (.A1(n37250), .A2(N12561), .ZN(N50689));
    NOR2X1 U37818 (.A1(N11427), .A2(n38457), .ZN(N50690));
    INVX1 U37819 (.I(N10261), .ZN(N50691));
    INVX1 U37820 (.I(N590), .ZN(n50692));
    INVX1 U37821 (.I(N8885), .ZN(N50693));
    NOR2X1 U37822 (.A1(n18041), .A2(N7395), .ZN(N50694));
    NANDX1 U37823 (.A1(n27297), .A2(n38929), .ZN(N50695));
    NOR2X1 U37824 (.A1(n19914), .A2(n23212), .ZN(N50696));
    NOR2X1 U37825 (.A1(n28711), .A2(n18787), .ZN(N50697));
    INVX1 U37826 (.I(n41605), .ZN(N50698));
    NOR2X1 U37827 (.A1(N7529), .A2(n14270), .ZN(N50699));
    NANDX1 U37828 (.A1(N1896), .A2(n34377), .ZN(N50700));
    INVX1 U37829 (.I(n14456), .ZN(N50701));
    NANDX1 U37830 (.A1(n22515), .A2(n42593), .ZN(N50702));
    INVX1 U37831 (.I(n32776), .ZN(N50703));
    INVX1 U37832 (.I(n13279), .ZN(n50704));
    INVX1 U37833 (.I(n42706), .ZN(N50705));
    NOR2X1 U37834 (.A1(N8223), .A2(n39780), .ZN(N50706));
    INVX1 U37835 (.I(n35520), .ZN(N50707));
    NOR2X1 U37836 (.A1(N9163), .A2(N1641), .ZN(N50708));
    NOR2X1 U37837 (.A1(n15726), .A2(n30351), .ZN(N50709));
    INVX1 U37838 (.I(n15189), .ZN(N50710));
    NANDX1 U37839 (.A1(n15608), .A2(n22717), .ZN(N50711));
    NOR2X1 U37840 (.A1(n43239), .A2(n14292), .ZN(N50712));
    NOR2X1 U37841 (.A1(n21175), .A2(n18428), .ZN(N50713));
    NOR2X1 U37842 (.A1(N217), .A2(N7228), .ZN(N50714));
    NOR2X1 U37843 (.A1(n22672), .A2(N7897), .ZN(N50715));
    INVX1 U37844 (.I(N12855), .ZN(N50716));
    INVX1 U37845 (.I(N3691), .ZN(N50717));
    INVX1 U37846 (.I(n36589), .ZN(N50718));
    NANDX1 U37847 (.A1(n35956), .A2(n18032), .ZN(N50719));
    INVX1 U37848 (.I(n37597), .ZN(N50720));
    NOR2X1 U37849 (.A1(n25245), .A2(n14155), .ZN(N50721));
    INVX1 U37850 (.I(n30113), .ZN(N50722));
    NANDX1 U37851 (.A1(N7942), .A2(n42509), .ZN(N50723));
    NANDX1 U37852 (.A1(N7708), .A2(n13329), .ZN(N50724));
    NOR2X1 U37853 (.A1(n18562), .A2(n31756), .ZN(N50725));
    NOR2X1 U37854 (.A1(N8458), .A2(n38983), .ZN(N50726));
    NANDX1 U37855 (.A1(n31130), .A2(n36559), .ZN(n50727));
    NOR2X1 U37856 (.A1(n33664), .A2(n23048), .ZN(N50728));
    NANDX1 U37857 (.A1(N948), .A2(N5844), .ZN(N50729));
    INVX1 U37858 (.I(n36904), .ZN(N50730));
    INVX1 U37859 (.I(N8390), .ZN(N50731));
    NOR2X1 U37860 (.A1(n36240), .A2(n33634), .ZN(N50732));
    NOR2X1 U37861 (.A1(n18254), .A2(n20274), .ZN(N50733));
    NOR2X1 U37862 (.A1(n26195), .A2(n19311), .ZN(N50734));
    INVX1 U37863 (.I(n33902), .ZN(N50735));
    NANDX1 U37864 (.A1(n17359), .A2(n42143), .ZN(N50736));
    INVX1 U37865 (.I(n30512), .ZN(N50737));
    NANDX1 U37866 (.A1(N6112), .A2(n22701), .ZN(N50738));
    NANDX1 U37867 (.A1(n42670), .A2(N7204), .ZN(N50739));
    INVX1 U37868 (.I(n22245), .ZN(n50740));
    INVX1 U37869 (.I(N8756), .ZN(N50741));
    NOR2X1 U37870 (.A1(n27420), .A2(n35339), .ZN(N50742));
    INVX1 U37871 (.I(n35810), .ZN(N50743));
    NANDX1 U37872 (.A1(n24089), .A2(n15651), .ZN(N50744));
    NANDX1 U37873 (.A1(n32023), .A2(n35925), .ZN(N50745));
    INVX1 U37874 (.I(n14745), .ZN(N50746));
    NANDX1 U37875 (.A1(n33567), .A2(n38327), .ZN(N50747));
    INVX1 U37876 (.I(n40606), .ZN(N50748));
    NOR2X1 U37877 (.A1(N1210), .A2(n27645), .ZN(N50749));
    NANDX1 U37878 (.A1(N7321), .A2(N6874), .ZN(N50750));
    INVX1 U37879 (.I(n39670), .ZN(N50751));
    NOR2X1 U37880 (.A1(n15758), .A2(N8122), .ZN(N50752));
    NOR2X1 U37881 (.A1(n14194), .A2(n25889), .ZN(N50753));
    NANDX1 U37882 (.A1(N6060), .A2(n13738), .ZN(N50754));
    NANDX1 U37883 (.A1(N8314), .A2(n27506), .ZN(N50755));
    INVX1 U37884 (.I(n24789), .ZN(N50756));
    NOR2X1 U37885 (.A1(n29205), .A2(N859), .ZN(N50757));
    INVX1 U37886 (.I(n40967), .ZN(N50758));
    NOR2X1 U37887 (.A1(n15335), .A2(n21255), .ZN(N50759));
    NOR2X1 U37888 (.A1(N8859), .A2(n22464), .ZN(N50760));
    INVX1 U37889 (.I(n32344), .ZN(N50761));
    NOR2X1 U37890 (.A1(n35116), .A2(n40293), .ZN(N50762));
    NANDX1 U37891 (.A1(n38872), .A2(N12579), .ZN(N50763));
    INVX1 U37892 (.I(n17386), .ZN(N50764));
    NANDX1 U37893 (.A1(n39350), .A2(n23319), .ZN(N50765));
    INVX1 U37894 (.I(n42767), .ZN(N50766));
    NOR2X1 U37895 (.A1(n20504), .A2(n26801), .ZN(N50767));
    NOR2X1 U37896 (.A1(n34972), .A2(n42856), .ZN(N50768));
    INVX1 U37897 (.I(n35830), .ZN(N50769));
    NOR2X1 U37898 (.A1(n20928), .A2(N6143), .ZN(N50770));
    INVX1 U37899 (.I(n31863), .ZN(N50771));
    NOR2X1 U37900 (.A1(n33737), .A2(N10854), .ZN(N50772));
    NOR2X1 U37901 (.A1(n22608), .A2(n30318), .ZN(N50773));
    NANDX1 U37902 (.A1(N9108), .A2(n35658), .ZN(N50774));
    NANDX1 U37903 (.A1(N11366), .A2(n38800), .ZN(N50775));
    INVX1 U37904 (.I(n27817), .ZN(N50776));
    INVX1 U37905 (.I(n19256), .ZN(N50777));
    NOR2X1 U37906 (.A1(n23652), .A2(n20204), .ZN(N50778));
    NANDX1 U37907 (.A1(n40132), .A2(n14432), .ZN(N50779));
    INVX1 U37908 (.I(n39515), .ZN(N50780));
    NANDX1 U37909 (.A1(n34048), .A2(N5587), .ZN(N50781));
    NOR2X1 U37910 (.A1(n40190), .A2(n30464), .ZN(N50782));
    NOR2X1 U37911 (.A1(N3458), .A2(n20728), .ZN(N50783));
    NOR2X1 U37912 (.A1(n15607), .A2(n33015), .ZN(N50784));
    INVX1 U37913 (.I(N9080), .ZN(N50785));
    NOR2X1 U37914 (.A1(N6107), .A2(n31104), .ZN(N50786));
    NANDX1 U37915 (.A1(N1434), .A2(n37361), .ZN(N50787));
    INVX1 U37916 (.I(n25790), .ZN(N50788));
    NOR2X1 U37917 (.A1(n34368), .A2(n39121), .ZN(N50789));
    NOR2X1 U37918 (.A1(N7934), .A2(n35780), .ZN(N50790));
    INVX1 U37919 (.I(N6152), .ZN(N50791));
    INVX1 U37920 (.I(n21531), .ZN(N50792));
    NOR2X1 U37921 (.A1(n27089), .A2(n16211), .ZN(N50793));
    NANDX1 U37922 (.A1(n14080), .A2(N9601), .ZN(N50794));
    INVX1 U37923 (.I(n24488), .ZN(N50795));
    NANDX1 U37924 (.A1(n35341), .A2(n14030), .ZN(N50796));
    INVX1 U37925 (.I(N948), .ZN(N50797));
    NANDX1 U37926 (.A1(n23551), .A2(n21731), .ZN(N50798));
    INVX1 U37927 (.I(n14664), .ZN(N50799));
    NOR2X1 U37928 (.A1(n39888), .A2(n40453), .ZN(N50800));
    NOR2X1 U37929 (.A1(n20463), .A2(n25782), .ZN(N50801));
    NOR2X1 U37930 (.A1(n18076), .A2(n18089), .ZN(N50802));
    NOR2X1 U37931 (.A1(n24228), .A2(n29271), .ZN(N50803));
    NOR2X1 U37932 (.A1(N10635), .A2(n12887), .ZN(N50804));
    NANDX1 U37933 (.A1(n26911), .A2(n16647), .ZN(N50805));
    INVX1 U37934 (.I(n13493), .ZN(N50806));
    INVX1 U37935 (.I(n34717), .ZN(N50807));
    NOR2X1 U37936 (.A1(N1371), .A2(n41841), .ZN(N50808));
    NANDX1 U37937 (.A1(N3731), .A2(n21919), .ZN(N50809));
    INVX1 U37938 (.I(N5786), .ZN(N50810));
    INVX1 U37939 (.I(n23016), .ZN(N50811));
    NANDX1 U37940 (.A1(n12922), .A2(n20817), .ZN(N50812));
    INVX1 U37941 (.I(n38703), .ZN(N50813));
    NANDX1 U37942 (.A1(n20098), .A2(N3000), .ZN(N50814));
    INVX1 U37943 (.I(N853), .ZN(N50815));
    INVX1 U37944 (.I(N8047), .ZN(N50816));
    NOR2X1 U37945 (.A1(N1685), .A2(n29639), .ZN(N50817));
    INVX1 U37946 (.I(N8011), .ZN(N50818));
    NANDX1 U37947 (.A1(n31250), .A2(n38824), .ZN(N50819));
    NANDX1 U37948 (.A1(n26290), .A2(n40194), .ZN(N50820));
    NANDX1 U37949 (.A1(N11957), .A2(n33604), .ZN(N50821));
    INVX1 U37950 (.I(n19354), .ZN(N50822));
    NANDX1 U37951 (.A1(n34511), .A2(n32049), .ZN(n50823));
    NOR2X1 U37952 (.A1(N3960), .A2(N9393), .ZN(N50824));
    INVX1 U37953 (.I(n42663), .ZN(N50825));
    NOR2X1 U37954 (.A1(N9917), .A2(N2190), .ZN(N50826));
    INVX1 U37955 (.I(N449), .ZN(N50827));
    NANDX1 U37956 (.A1(N7953), .A2(n34768), .ZN(N50828));
    NANDX1 U37957 (.A1(n27272), .A2(n19373), .ZN(N50829));
    NOR2X1 U37958 (.A1(N1159), .A2(N7150), .ZN(N50830));
    INVX1 U37959 (.I(n32594), .ZN(N50831));
    NOR2X1 U37960 (.A1(n15586), .A2(n18925), .ZN(N50832));
    NOR2X1 U37961 (.A1(N5717), .A2(n27174), .ZN(N50833));
    NANDX1 U37962 (.A1(n34786), .A2(N7892), .ZN(N50834));
    NANDX1 U37963 (.A1(n22582), .A2(N11851), .ZN(N50835));
    NOR2X1 U37964 (.A1(N2081), .A2(N721), .ZN(N50836));
    NOR2X1 U37965 (.A1(N1677), .A2(n36062), .ZN(N50837));
    INVX1 U37966 (.I(n35277), .ZN(N50838));
    NOR2X1 U37967 (.A1(n26538), .A2(n26572), .ZN(N50839));
    INVX1 U37968 (.I(N10337), .ZN(N50840));
    NOR2X1 U37969 (.A1(n22592), .A2(N1175), .ZN(N50841));
    NANDX1 U37970 (.A1(n31135), .A2(n33768), .ZN(N50842));
    INVX1 U37971 (.I(N3248), .ZN(N50843));
    NANDX1 U37972 (.A1(n14021), .A2(n42117), .ZN(N50844));
    NANDX1 U37973 (.A1(n24976), .A2(n33430), .ZN(N50845));
    NANDX1 U37974 (.A1(N3867), .A2(N2219), .ZN(N50846));
    NOR2X1 U37975 (.A1(N2470), .A2(n37451), .ZN(N50847));
    NANDX1 U37976 (.A1(n31468), .A2(n39127), .ZN(N50848));
    INVX1 U37977 (.I(N6581), .ZN(N50849));
    NANDX1 U37978 (.A1(N2060), .A2(n33118), .ZN(N50850));
    NANDX1 U37979 (.A1(n34291), .A2(n33134), .ZN(N50851));
    NOR2X1 U37980 (.A1(N3090), .A2(n34308), .ZN(N50852));
    INVX1 U37981 (.I(n34224), .ZN(N50853));
    INVX1 U37982 (.I(n27902), .ZN(n50854));
    NANDX1 U37983 (.A1(n23502), .A2(n41922), .ZN(N50855));
    NOR2X1 U37984 (.A1(N6102), .A2(n13106), .ZN(N50856));
    NANDX1 U37985 (.A1(n29745), .A2(n16972), .ZN(N50857));
    INVX1 U37986 (.I(n21766), .ZN(N50858));
    INVX1 U37987 (.I(n34782), .ZN(N50859));
    INVX1 U37988 (.I(n30269), .ZN(N50860));
    NANDX1 U37989 (.A1(n32992), .A2(n36849), .ZN(n50861));
    INVX1 U37990 (.I(n35051), .ZN(N50862));
    NOR2X1 U37991 (.A1(N966), .A2(n15549), .ZN(n50863));
    NANDX1 U37992 (.A1(N7148), .A2(n18638), .ZN(N50864));
    INVX1 U37993 (.I(N2310), .ZN(N50865));
    NANDX1 U37994 (.A1(n21272), .A2(n30211), .ZN(N50866));
    NOR2X1 U37995 (.A1(n34453), .A2(n18341), .ZN(N50867));
    NANDX1 U37996 (.A1(n30234), .A2(n31446), .ZN(N50868));
    INVX1 U37997 (.I(n16506), .ZN(N50869));
    NOR2X1 U37998 (.A1(n34138), .A2(n38272), .ZN(N50870));
    NOR2X1 U37999 (.A1(n25447), .A2(N9307), .ZN(N50871));
    INVX1 U38000 (.I(n35243), .ZN(N50872));
    INVX1 U38001 (.I(n27391), .ZN(N50873));
    NOR2X1 U38002 (.A1(n23557), .A2(N93), .ZN(N50874));
    NOR2X1 U38003 (.A1(n28785), .A2(N5927), .ZN(N50875));
    NOR2X1 U38004 (.A1(N3951), .A2(N2597), .ZN(N50876));
    INVX1 U38005 (.I(N3020), .ZN(n50877));
    INVX1 U38006 (.I(N9017), .ZN(N50878));
    NANDX1 U38007 (.A1(n37681), .A2(n17037), .ZN(N50879));
    NOR2X1 U38008 (.A1(n24442), .A2(n38162), .ZN(N50880));
    INVX1 U38009 (.I(n40948), .ZN(N50881));
    NANDX1 U38010 (.A1(N11463), .A2(n25427), .ZN(N50882));
    NANDX1 U38011 (.A1(n26590), .A2(n24413), .ZN(N50883));
    NANDX1 U38012 (.A1(n18360), .A2(n12919), .ZN(N50884));
    NANDX1 U38013 (.A1(n40536), .A2(n26155), .ZN(N50885));
    NANDX1 U38014 (.A1(n30526), .A2(N11467), .ZN(N50886));
    NOR2X1 U38015 (.A1(N7022), .A2(N5097), .ZN(N50887));
    NOR2X1 U38016 (.A1(n39620), .A2(n41268), .ZN(N50888));
    INVX1 U38017 (.I(n38317), .ZN(n50889));
    NOR2X1 U38018 (.A1(n29555), .A2(N11881), .ZN(n50890));
    NOR2X1 U38019 (.A1(N204), .A2(n39723), .ZN(N50891));
    NOR2X1 U38020 (.A1(n30831), .A2(n29037), .ZN(N50892));
    NOR2X1 U38021 (.A1(N12785), .A2(N11776), .ZN(N50893));
    NANDX1 U38022 (.A1(n26878), .A2(n18210), .ZN(N50894));
    INVX1 U38023 (.I(n39796), .ZN(N50895));
    NOR2X1 U38024 (.A1(N544), .A2(N12158), .ZN(N50896));
    INVX1 U38025 (.I(n20749), .ZN(n50897));
    NANDX1 U38026 (.A1(n41040), .A2(n27771), .ZN(N50898));
    NANDX1 U38027 (.A1(n19367), .A2(n13598), .ZN(N50899));
    NOR2X1 U38028 (.A1(N921), .A2(n41594), .ZN(N50900));
    NOR2X1 U38029 (.A1(n20155), .A2(n43155), .ZN(N50901));
    NANDX1 U38030 (.A1(n20358), .A2(n39405), .ZN(N50902));
    NOR2X1 U38031 (.A1(N7717), .A2(n14649), .ZN(N50903));
    NANDX1 U38032 (.A1(n20501), .A2(n26424), .ZN(N50904));
    INVX1 U38033 (.I(n37058), .ZN(N50905));
    NANDX1 U38034 (.A1(n25082), .A2(n33381), .ZN(N50906));
    INVX1 U38035 (.I(n25625), .ZN(n50907));
    NANDX1 U38036 (.A1(N10919), .A2(n36054), .ZN(N50908));
    NANDX1 U38037 (.A1(N8487), .A2(n20352), .ZN(n50909));
    INVX1 U38038 (.I(n17533), .ZN(N50910));
    NOR2X1 U38039 (.A1(N6493), .A2(n18453), .ZN(N50911));
    NOR2X1 U38040 (.A1(N6251), .A2(n38607), .ZN(N50912));
    NOR2X1 U38041 (.A1(n29546), .A2(n15492), .ZN(N50913));
    NOR2X1 U38042 (.A1(N10230), .A2(n12888), .ZN(N50914));
    NOR2X1 U38043 (.A1(N3238), .A2(n23069), .ZN(N50915));
    INVX1 U38044 (.I(n24839), .ZN(N50916));
    NOR2X1 U38045 (.A1(n28637), .A2(N6448), .ZN(n50917));
    NOR2X1 U38046 (.A1(n17718), .A2(n21752), .ZN(N50918));
    INVX1 U38047 (.I(n18317), .ZN(N50919));
    NANDX1 U38048 (.A1(N3357), .A2(n16483), .ZN(N50920));
    NOR2X1 U38049 (.A1(n37126), .A2(n34015), .ZN(N50921));
    NOR2X1 U38050 (.A1(N147), .A2(n42147), .ZN(N50922));
    NOR2X1 U38051 (.A1(n39549), .A2(n37281), .ZN(N50923));
    NANDX1 U38052 (.A1(n15302), .A2(n42452), .ZN(N50924));
    NANDX1 U38053 (.A1(n25531), .A2(N1548), .ZN(N50925));
    NANDX1 U38054 (.A1(n18448), .A2(n24616), .ZN(N50926));
    NANDX1 U38055 (.A1(n43286), .A2(n41269), .ZN(N50927));
    NANDX1 U38056 (.A1(N6261), .A2(n37511), .ZN(N50928));
    NOR2X1 U38057 (.A1(n28013), .A2(n25499), .ZN(N50929));
    INVX1 U38058 (.I(n32025), .ZN(N50930));
    NOR2X1 U38059 (.A1(N3050), .A2(n12917), .ZN(n50931));
    INVX1 U38060 (.I(n37064), .ZN(N50932));
    NOR2X1 U38061 (.A1(N2015), .A2(n35738), .ZN(N50933));
    NOR2X1 U38062 (.A1(n41563), .A2(n19226), .ZN(N50934));
    NANDX1 U38063 (.A1(n13393), .A2(N7885), .ZN(n50935));
    NOR2X1 U38064 (.A1(n28603), .A2(N9432), .ZN(N50936));
    NANDX1 U38065 (.A1(n36731), .A2(n23727), .ZN(N50937));
    NOR2X1 U38066 (.A1(n36544), .A2(n21524), .ZN(n50938));
    NOR2X1 U38067 (.A1(n32485), .A2(N5242), .ZN(N50939));
    NANDX1 U38068 (.A1(N6705), .A2(n30740), .ZN(n50940));
    NANDX1 U38069 (.A1(n38729), .A2(N5803), .ZN(N50941));
    NOR2X1 U38070 (.A1(N8173), .A2(N7671), .ZN(N50942));
    NANDX1 U38071 (.A1(n15289), .A2(N9685), .ZN(n50943));
    NANDX1 U38072 (.A1(n38355), .A2(n40927), .ZN(N50944));
    INVX1 U38073 (.I(n34691), .ZN(N50945));
    NOR2X1 U38074 (.A1(n41472), .A2(N1021), .ZN(N50946));
    INVX1 U38075 (.I(n40584), .ZN(n50947));
    NANDX1 U38076 (.A1(N12068), .A2(n20838), .ZN(n50948));
    NOR2X1 U38077 (.A1(N5139), .A2(n42361), .ZN(N50949));
    NANDX1 U38078 (.A1(n27303), .A2(n37283), .ZN(N50950));
    INVX1 U38079 (.I(n34007), .ZN(n50951));
    INVX1 U38080 (.I(N513), .ZN(N50952));
    INVX1 U38081 (.I(n20032), .ZN(N50953));
    NANDX1 U38082 (.A1(n27116), .A2(n27702), .ZN(N50954));
    NOR2X1 U38083 (.A1(n32085), .A2(n27066), .ZN(N50955));
    NANDX1 U38084 (.A1(n16647), .A2(n24521), .ZN(N50956));
    NOR2X1 U38085 (.A1(N7866), .A2(n25047), .ZN(N50957));
    INVX1 U38086 (.I(n42038), .ZN(N50958));
    NANDX1 U38087 (.A1(n35999), .A2(n34227), .ZN(N50959));
    NANDX1 U38088 (.A1(n13365), .A2(n13913), .ZN(N50960));
    NOR2X1 U38089 (.A1(N1933), .A2(N8254), .ZN(N50961));
    INVX1 U38090 (.I(n39215), .ZN(N50962));
    INVX1 U38091 (.I(n25107), .ZN(N50963));
    INVX1 U38092 (.I(n29485), .ZN(N50964));
    INVX1 U38093 (.I(n19684), .ZN(N50965));
    INVX1 U38094 (.I(n17373), .ZN(N50966));
    INVX1 U38095 (.I(n18290), .ZN(n50967));
    INVX1 U38096 (.I(n20659), .ZN(N50968));
    NANDX1 U38097 (.A1(N12312), .A2(n34859), .ZN(N50969));
    NANDX1 U38098 (.A1(N9857), .A2(n16434), .ZN(N50970));
    NANDX1 U38099 (.A1(N8422), .A2(n16817), .ZN(N50971));
    NANDX1 U38100 (.A1(n42648), .A2(n18948), .ZN(N50972));
    NANDX1 U38101 (.A1(N2768), .A2(n26217), .ZN(N50973));
    NANDX1 U38102 (.A1(N701), .A2(n17316), .ZN(n50974));
    NANDX1 U38103 (.A1(n29673), .A2(n32102), .ZN(N50975));
    NANDX1 U38104 (.A1(n15685), .A2(n22359), .ZN(N50976));
    NOR2X1 U38105 (.A1(N7883), .A2(n29412), .ZN(n50977));
    NOR2X1 U38106 (.A1(n26172), .A2(n25076), .ZN(N50978));
    INVX1 U38107 (.I(n41442), .ZN(N50979));
    INVX1 U38108 (.I(n38833), .ZN(N50980));
    NANDX1 U38109 (.A1(N3771), .A2(N11794), .ZN(N50981));
    NANDX1 U38110 (.A1(N1873), .A2(n18291), .ZN(N50982));
    INVX1 U38111 (.I(n34200), .ZN(N50983));
    NANDX1 U38112 (.A1(n25250), .A2(n36968), .ZN(N50984));
    INVX1 U38113 (.I(n43366), .ZN(N50985));
    NANDX1 U38114 (.A1(n26977), .A2(n13753), .ZN(N50986));
    INVX1 U38115 (.I(n15607), .ZN(n50987));
    NOR2X1 U38116 (.A1(n18913), .A2(n27645), .ZN(N50988));
    INVX1 U38117 (.I(n16476), .ZN(N50989));
    NOR2X1 U38118 (.A1(N10622), .A2(n42647), .ZN(N50990));
    INVX1 U38119 (.I(n14596), .ZN(N50991));
    NANDX1 U38120 (.A1(n32574), .A2(n43109), .ZN(N50992));
    INVX1 U38121 (.I(n26025), .ZN(N50993));
    NANDX1 U38122 (.A1(n28749), .A2(n27897), .ZN(N50994));
    NANDX1 U38123 (.A1(n17174), .A2(n18624), .ZN(N50995));
    NOR2X1 U38124 (.A1(n32103), .A2(N1799), .ZN(N50996));
    NOR2X1 U38125 (.A1(n31997), .A2(n29147), .ZN(N50997));
    NOR2X1 U38126 (.A1(N2277), .A2(n32375), .ZN(N50998));
    INVX1 U38127 (.I(n29541), .ZN(N50999));
    NANDX1 U38128 (.A1(n18621), .A2(n13375), .ZN(N51000));
    NOR2X1 U38129 (.A1(n32205), .A2(n23996), .ZN(N51001));
    INVX1 U38130 (.I(n17072), .ZN(N51002));
    INVX1 U38131 (.I(n33121), .ZN(N51003));
    INVX1 U38132 (.I(n27908), .ZN(N51004));
    NOR2X1 U38133 (.A1(n21877), .A2(n18697), .ZN(N51005));
    NOR2X1 U38134 (.A1(N6301), .A2(n27777), .ZN(N51006));
    NOR2X1 U38135 (.A1(n14605), .A2(n20301), .ZN(N51007));
    NANDX1 U38136 (.A1(N6083), .A2(n22487), .ZN(N51008));
    INVX1 U38137 (.I(n35229), .ZN(N51009));
    INVX1 U38138 (.I(n14673), .ZN(N51010));
    NOR2X1 U38139 (.A1(n42625), .A2(N741), .ZN(N51011));
    NANDX1 U38140 (.A1(N7453), .A2(n14115), .ZN(N51012));
    NANDX1 U38141 (.A1(n39657), .A2(n27791), .ZN(N51013));
    NANDX1 U38142 (.A1(n13256), .A2(N2270), .ZN(N51014));
    INVX1 U38143 (.I(N9109), .ZN(N51015));
    NANDX1 U38144 (.A1(N7067), .A2(n30985), .ZN(N51016));
    NOR2X1 U38145 (.A1(n35455), .A2(n26966), .ZN(N51017));
    NOR2X1 U38146 (.A1(n37544), .A2(n31250), .ZN(N51018));
    INVX1 U38147 (.I(n28264), .ZN(N51019));
    NANDX1 U38148 (.A1(N11852), .A2(n40660), .ZN(N51020));
    NOR2X1 U38149 (.A1(n20028), .A2(N11861), .ZN(N51021));
    NOR2X1 U38150 (.A1(N8860), .A2(N2281), .ZN(N51022));
    NANDX1 U38151 (.A1(n16312), .A2(N6076), .ZN(N51023));
    INVX1 U38152 (.I(N12497), .ZN(n51024));
    INVX1 U38153 (.I(N2185), .ZN(n51025));
    INVX1 U38154 (.I(n25815), .ZN(N51026));
    INVX1 U38155 (.I(n14220), .ZN(N51027));
    INVX1 U38156 (.I(n39510), .ZN(N51028));
    INVX1 U38157 (.I(n20111), .ZN(N51029));
    NOR2X1 U38158 (.A1(n18378), .A2(n32648), .ZN(N51030));
    NANDX1 U38159 (.A1(n39307), .A2(n22013), .ZN(N51031));
    INVX1 U38160 (.I(n33166), .ZN(N51032));
    NANDX1 U38161 (.A1(n20054), .A2(n41614), .ZN(N51033));
    INVX1 U38162 (.I(n21594), .ZN(N51034));
    INVX1 U38163 (.I(n19278), .ZN(n51035));
    NANDX1 U38164 (.A1(N172), .A2(n25269), .ZN(N51036));
    NANDX1 U38165 (.A1(n28050), .A2(n27445), .ZN(N51037));
    NANDX1 U38166 (.A1(n30235), .A2(n42877), .ZN(n51038));
    INVX1 U38167 (.I(n19206), .ZN(N51039));
    NOR2X1 U38168 (.A1(N7075), .A2(N4923), .ZN(N51040));
    INVX1 U38169 (.I(n27185), .ZN(N51041));
    NANDX1 U38170 (.A1(n13093), .A2(n16360), .ZN(n51042));
    INVX1 U38171 (.I(n42079), .ZN(N51043));
    INVX1 U38172 (.I(N10410), .ZN(N51044));
    INVX1 U38173 (.I(n28763), .ZN(N51045));
    NANDX1 U38174 (.A1(n19594), .A2(n28861), .ZN(n51046));
    NOR2X1 U38175 (.A1(n29674), .A2(n37818), .ZN(N51047));
    NANDX1 U38176 (.A1(n19526), .A2(n19615), .ZN(N51048));
    NOR2X1 U38177 (.A1(n37255), .A2(N3587), .ZN(N51049));
    INVX1 U38178 (.I(n13697), .ZN(N51050));
    NOR2X1 U38179 (.A1(N2874), .A2(n32902), .ZN(n51051));
    INVX1 U38180 (.I(n43100), .ZN(N51052));
    NANDX1 U38181 (.A1(n34162), .A2(n26813), .ZN(N51053));
    INVX1 U38182 (.I(n36935), .ZN(N51054));
    NANDX1 U38183 (.A1(n30821), .A2(n35541), .ZN(N51055));
    INVX1 U38184 (.I(n30910), .ZN(N51056));
    NOR2X1 U38185 (.A1(n35874), .A2(N7581), .ZN(N51057));
    INVX1 U38186 (.I(n21263), .ZN(N51058));
    NOR2X1 U38187 (.A1(n42148), .A2(n15608), .ZN(N51059));
    NANDX1 U38188 (.A1(N7881), .A2(n24902), .ZN(N51060));
    NANDX1 U38189 (.A1(N1664), .A2(n18169), .ZN(N51061));
    NANDX1 U38190 (.A1(n15360), .A2(N10839), .ZN(N51062));
    INVX1 U38191 (.I(n37942), .ZN(n51063));
    NOR2X1 U38192 (.A1(n18650), .A2(n21973), .ZN(N51064));
    INVX1 U38193 (.I(n35142), .ZN(N51065));
    INVX1 U38194 (.I(n13797), .ZN(N51066));
    NANDX1 U38195 (.A1(n42278), .A2(N5865), .ZN(N51067));
    NANDX1 U38196 (.A1(n19395), .A2(N9066), .ZN(N51068));
    INVX1 U38197 (.I(n26976), .ZN(N51069));
    INVX1 U38198 (.I(n34976), .ZN(N51070));
    INVX1 U38199 (.I(N9895), .ZN(N51071));
    NANDX1 U38200 (.A1(n29844), .A2(n17776), .ZN(N51072));
    INVX1 U38201 (.I(n14843), .ZN(N51073));
    INVX1 U38202 (.I(n39861), .ZN(N51074));
    INVX1 U38203 (.I(n24478), .ZN(N51075));
    NOR2X1 U38204 (.A1(N6542), .A2(n18947), .ZN(N51076));
    NANDX1 U38205 (.A1(n14871), .A2(n30600), .ZN(N51077));
    NOR2X1 U38206 (.A1(n39693), .A2(n42057), .ZN(N51078));
    INVX1 U38207 (.I(N10422), .ZN(N51079));
    INVX1 U38208 (.I(n23075), .ZN(N51080));
    NOR2X1 U38209 (.A1(N6464), .A2(n21820), .ZN(N51081));
    NOR2X1 U38210 (.A1(n33439), .A2(n33039), .ZN(N51082));
    NANDX1 U38211 (.A1(N2147), .A2(n42933), .ZN(N51083));
    NOR2X1 U38212 (.A1(n21671), .A2(N6916), .ZN(N51084));
    INVX1 U38213 (.I(n36513), .ZN(N51085));
    NOR2X1 U38214 (.A1(n31183), .A2(n24032), .ZN(N51086));
    NANDX1 U38215 (.A1(n28090), .A2(n20253), .ZN(N51087));
    NANDX1 U38216 (.A1(N11169), .A2(n35124), .ZN(n51088));
    NANDX1 U38217 (.A1(n14583), .A2(n31344), .ZN(N51089));
    NOR2X1 U38218 (.A1(n42112), .A2(n31445), .ZN(N51090));
    INVX1 U38219 (.I(N11394), .ZN(N51091));
    NOR2X1 U38220 (.A1(n28382), .A2(n33213), .ZN(n51092));
    NANDX1 U38221 (.A1(N8028), .A2(N12459), .ZN(N51093));
    NOR2X1 U38222 (.A1(n43327), .A2(N11920), .ZN(N51094));
    NOR2X1 U38223 (.A1(n21525), .A2(n18835), .ZN(N51095));
    INVX1 U38224 (.I(N4245), .ZN(N51096));
    INVX1 U38225 (.I(n38251), .ZN(N51097));
    NANDX1 U38226 (.A1(n21588), .A2(n22868), .ZN(N51098));
    NANDX1 U38227 (.A1(n16933), .A2(n23716), .ZN(n51099));
    NOR2X1 U38228 (.A1(n42878), .A2(n38298), .ZN(n51100));
    NANDX1 U38229 (.A1(n23934), .A2(n26618), .ZN(N51101));
    NANDX1 U38230 (.A1(N2380), .A2(n27691), .ZN(N51102));
    INVX1 U38231 (.I(n20441), .ZN(N51103));
    NOR2X1 U38232 (.A1(N3616), .A2(n18148), .ZN(n51104));
    NOR2X1 U38233 (.A1(n18773), .A2(n18002), .ZN(N51105));
    INVX1 U38234 (.I(n24200), .ZN(N51106));
    INVX1 U38235 (.I(n40004), .ZN(N51107));
    INVX1 U38236 (.I(N299), .ZN(N51108));
    NANDX1 U38237 (.A1(n15726), .A2(n18255), .ZN(n51109));
    INVX1 U38238 (.I(n38593), .ZN(N51110));
    INVX1 U38239 (.I(n38959), .ZN(N51111));
    NOR2X1 U38240 (.A1(n42851), .A2(n38364), .ZN(N51112));
    NOR2X1 U38241 (.A1(N6789), .A2(n18826), .ZN(N51113));
    INVX1 U38242 (.I(N12492), .ZN(N51114));
    INVX1 U38243 (.I(n37009), .ZN(N51115));
    NOR2X1 U38244 (.A1(n21005), .A2(N648), .ZN(N51116));
    INVX1 U38245 (.I(n39152), .ZN(N51117));
    INVX1 U38246 (.I(n29327), .ZN(N51118));
    NOR2X1 U38247 (.A1(n31066), .A2(N10054), .ZN(N51119));
    INVX1 U38248 (.I(n17277), .ZN(N51120));
    INVX1 U38249 (.I(n32865), .ZN(N51121));
    NOR2X1 U38250 (.A1(N3254), .A2(N7647), .ZN(N51122));
    NOR2X1 U38251 (.A1(n31526), .A2(N10318), .ZN(N51123));
    INVX1 U38252 (.I(n29721), .ZN(N51124));
    INVX1 U38253 (.I(n30120), .ZN(N51125));
    NOR2X1 U38254 (.A1(n16484), .A2(n38625), .ZN(N51126));
    NOR2X1 U38255 (.A1(n18655), .A2(n39189), .ZN(N51127));
    NANDX1 U38256 (.A1(N2762), .A2(n16721), .ZN(N51128));
    NANDX1 U38257 (.A1(n13315), .A2(N12401), .ZN(N51129));
    NANDX1 U38258 (.A1(n42641), .A2(n15762), .ZN(N51130));
    NOR2X1 U38259 (.A1(n42374), .A2(n15176), .ZN(N51131));
    INVX1 U38260 (.I(n29902), .ZN(N51132));
    NOR2X1 U38261 (.A1(N4935), .A2(n22835), .ZN(N51133));
    NANDX1 U38262 (.A1(N11524), .A2(N568), .ZN(N51134));
    NANDX1 U38263 (.A1(N3280), .A2(n30289), .ZN(N51135));
    NANDX1 U38264 (.A1(n23080), .A2(N9558), .ZN(N51136));
    NANDX1 U38265 (.A1(N7912), .A2(n31298), .ZN(N51137));
    NOR2X1 U38266 (.A1(N3629), .A2(n36254), .ZN(n51138));
    NANDX1 U38267 (.A1(N10029), .A2(n41857), .ZN(N51139));
    NOR2X1 U38268 (.A1(n22429), .A2(n13886), .ZN(N51140));
    INVX1 U38269 (.I(n27870), .ZN(N51141));
    NANDX1 U38270 (.A1(n29911), .A2(n43046), .ZN(N51142));
    NANDX1 U38271 (.A1(N6020), .A2(n26974), .ZN(N51143));
    NANDX1 U38272 (.A1(n28855), .A2(n18548), .ZN(N51144));
    NOR2X1 U38273 (.A1(n29422), .A2(n20440), .ZN(N51145));
    INVX1 U38274 (.I(N5918), .ZN(N51146));
    NOR2X1 U38275 (.A1(N5734), .A2(n15476), .ZN(N51147));
    INVX1 U38276 (.I(n13646), .ZN(N51148));
    NOR2X1 U38277 (.A1(n42709), .A2(N6954), .ZN(n51149));
    NANDX1 U38278 (.A1(n28082), .A2(n16982), .ZN(N51150));
    NANDX1 U38279 (.A1(n26770), .A2(n29091), .ZN(N51151));
    NANDX1 U38280 (.A1(n14307), .A2(n13488), .ZN(N51152));
    NOR2X1 U38281 (.A1(N745), .A2(N2741), .ZN(N51153));
    NOR2X1 U38282 (.A1(N6764), .A2(n29714), .ZN(N51154));
    INVX1 U38283 (.I(n25298), .ZN(N51155));
    NOR2X1 U38284 (.A1(n20226), .A2(N928), .ZN(N51156));
    NOR2X1 U38285 (.A1(N2881), .A2(N6845), .ZN(N51157));
    NANDX1 U38286 (.A1(N8614), .A2(N12000), .ZN(n51158));
    INVX1 U38287 (.I(n22259), .ZN(N51159));
    INVX1 U38288 (.I(n21514), .ZN(N51160));
    NANDX1 U38289 (.A1(n23893), .A2(N6123), .ZN(N51161));
    NANDX1 U38290 (.A1(n41191), .A2(n22573), .ZN(N51162));
    NANDX1 U38291 (.A1(n28901), .A2(n26559), .ZN(N51163));
    NOR2X1 U38292 (.A1(n33591), .A2(n16983), .ZN(N51164));
    NOR2X1 U38293 (.A1(n21838), .A2(n13426), .ZN(N51165));
    NOR2X1 U38294 (.A1(n42048), .A2(n38724), .ZN(N51166));
    NANDX1 U38295 (.A1(N8482), .A2(n39651), .ZN(N51167));
    NANDX1 U38296 (.A1(N11362), .A2(N3023), .ZN(N51168));
    NANDX1 U38297 (.A1(n19975), .A2(n15023), .ZN(N51169));
    NANDX1 U38298 (.A1(n31914), .A2(N9682), .ZN(N51170));
    NANDX1 U38299 (.A1(n17653), .A2(n23255), .ZN(N51171));
    NANDX1 U38300 (.A1(N10054), .A2(n20973), .ZN(N51172));
    NANDX1 U38301 (.A1(n31545), .A2(N6401), .ZN(N51173));
    NANDX1 U38302 (.A1(N12732), .A2(n29671), .ZN(N51174));
    NOR2X1 U38303 (.A1(n40131), .A2(n41188), .ZN(N51175));
    NOR2X1 U38304 (.A1(N10299), .A2(n39764), .ZN(N51176));
    NOR2X1 U38305 (.A1(N8089), .A2(n37925), .ZN(N51177));
    NOR2X1 U38306 (.A1(n20786), .A2(N5814), .ZN(N51178));
    NOR2X1 U38307 (.A1(n16305), .A2(n15468), .ZN(N51179));
    NANDX1 U38308 (.A1(n34101), .A2(N3909), .ZN(N51180));
    NOR2X1 U38309 (.A1(n29938), .A2(N11242), .ZN(N51181));
    NOR2X1 U38310 (.A1(n21578), .A2(n21295), .ZN(N51182));
    NANDX1 U38311 (.A1(n25469), .A2(n42520), .ZN(N51183));
    INVX1 U38312 (.I(N12447), .ZN(N51184));
    INVX1 U38313 (.I(n21766), .ZN(N51185));
    INVX1 U38314 (.I(N8437), .ZN(N51186));
    NOR2X1 U38315 (.A1(n23471), .A2(N8415), .ZN(N51187));
    NANDX1 U38316 (.A1(n15467), .A2(n16503), .ZN(N51188));
    NOR2X1 U38317 (.A1(n13961), .A2(n26969), .ZN(N51189));
    NOR2X1 U38318 (.A1(n38310), .A2(n43273), .ZN(N51190));
    NANDX1 U38319 (.A1(n23888), .A2(n23582), .ZN(N51191));
    NOR2X1 U38320 (.A1(n19148), .A2(n43199), .ZN(n51192));
    NANDX1 U38321 (.A1(n37662), .A2(N10984), .ZN(N51193));
    INVX1 U38322 (.I(n33676), .ZN(N51194));
    NANDX1 U38323 (.A1(n25716), .A2(n25771), .ZN(N51195));
    NOR2X1 U38324 (.A1(n27174), .A2(N4064), .ZN(n51196));
    NOR2X1 U38325 (.A1(n35610), .A2(n13224), .ZN(N51197));
    INVX1 U38326 (.I(n33704), .ZN(N51198));
    INVX1 U38327 (.I(n19489), .ZN(n51199));
    NANDX1 U38328 (.A1(n18579), .A2(n23130), .ZN(N51200));
    NANDX1 U38329 (.A1(n13976), .A2(n17967), .ZN(N51201));
    NOR2X1 U38330 (.A1(n14520), .A2(n41854), .ZN(N51202));
    INVX1 U38331 (.I(n18972), .ZN(N51203));
    NANDX1 U38332 (.A1(n36171), .A2(n34666), .ZN(N51204));
    INVX1 U38333 (.I(N3682), .ZN(N51205));
    INVX1 U38334 (.I(n35075), .ZN(N51206));
    NANDX1 U38335 (.A1(N105), .A2(n17373), .ZN(N51207));
    NANDX1 U38336 (.A1(n27278), .A2(N11116), .ZN(N51208));
    NOR2X1 U38337 (.A1(N9095), .A2(n24339), .ZN(N51209));
    INVX1 U38338 (.I(n42798), .ZN(N51210));
    NOR2X1 U38339 (.A1(n39302), .A2(N6060), .ZN(N51211));
    NOR2X1 U38340 (.A1(n18959), .A2(n29442), .ZN(N51212));
    NOR2X1 U38341 (.A1(n26605), .A2(N9153), .ZN(N51213));
    INVX1 U38342 (.I(n24987), .ZN(N51214));
    NOR2X1 U38343 (.A1(N1474), .A2(n32196), .ZN(N51215));
    INVX1 U38344 (.I(n25819), .ZN(N51216));
    NANDX1 U38345 (.A1(n41976), .A2(N208), .ZN(N51217));
    INVX1 U38346 (.I(n28317), .ZN(n51218));
    INVX1 U38347 (.I(n32248), .ZN(N51219));
    INVX1 U38348 (.I(n27589), .ZN(N51220));
    INVX1 U38349 (.I(n15236), .ZN(N51221));
    INVX1 U38350 (.I(N3590), .ZN(N51222));
    INVX1 U38351 (.I(n36009), .ZN(N51223));
    NOR2X1 U38352 (.A1(n20558), .A2(n31748), .ZN(N51224));
    NANDX1 U38353 (.A1(n29197), .A2(n17718), .ZN(N51225));
    NANDX1 U38354 (.A1(N12329), .A2(n16550), .ZN(N51226));
    NOR2X1 U38355 (.A1(n26995), .A2(n18673), .ZN(n51227));
    NOR2X1 U38356 (.A1(N5398), .A2(n13495), .ZN(N51228));
    NANDX1 U38357 (.A1(n38992), .A2(N1678), .ZN(N51229));
    NOR2X1 U38358 (.A1(N10395), .A2(n19674), .ZN(N51230));
    NOR2X1 U38359 (.A1(n32323), .A2(n19118), .ZN(N51231));
    NANDX1 U38360 (.A1(n21893), .A2(n34353), .ZN(N51232));
    NOR2X1 U38361 (.A1(n25482), .A2(N5289), .ZN(N51233));
    NOR2X1 U38362 (.A1(n18293), .A2(n25847), .ZN(N51234));
    NOR2X1 U38363 (.A1(N8583), .A2(N1251), .ZN(N51235));
    NANDX1 U38364 (.A1(N9), .A2(n13579), .ZN(N51236));
    NANDX1 U38365 (.A1(n17408), .A2(n30254), .ZN(N51237));
    NANDX1 U38366 (.A1(n15641), .A2(n35651), .ZN(N51238));
    NOR2X1 U38367 (.A1(N6541), .A2(n20850), .ZN(N51239));
    NANDX1 U38368 (.A1(n30800), .A2(n31245), .ZN(N51240));
    NOR2X1 U38369 (.A1(N11898), .A2(N9775), .ZN(n51241));
    INVX1 U38370 (.I(n20585), .ZN(N51242));
    NOR2X1 U38371 (.A1(n18571), .A2(N12163), .ZN(n51243));
    NANDX1 U38372 (.A1(n23859), .A2(n29428), .ZN(N51244));
    NOR2X1 U38373 (.A1(n39385), .A2(n24649), .ZN(N51245));
    NOR2X1 U38374 (.A1(n40635), .A2(n27267), .ZN(N51246));
    NANDX1 U38375 (.A1(N422), .A2(n13282), .ZN(n51247));
    NANDX1 U38376 (.A1(n20355), .A2(n40802), .ZN(N51248));
    NOR2X1 U38377 (.A1(N12533), .A2(n38343), .ZN(N51249));
    INVX1 U38378 (.I(n33383), .ZN(N51250));
    NOR2X1 U38379 (.A1(n15874), .A2(N10835), .ZN(N51251));
    NOR2X1 U38380 (.A1(n27772), .A2(n20609), .ZN(N51252));
    NOR2X1 U38381 (.A1(n38036), .A2(n41955), .ZN(N51253));
    NOR2X1 U38382 (.A1(n39878), .A2(n34991), .ZN(N51254));
    NANDX1 U38383 (.A1(n15514), .A2(N2847), .ZN(N51255));
    NANDX1 U38384 (.A1(n40162), .A2(N12438), .ZN(N51256));
    INVX1 U38385 (.I(n23957), .ZN(N51257));
    NANDX1 U38386 (.A1(n24996), .A2(n26918), .ZN(N51258));
    INVX1 U38387 (.I(N1878), .ZN(N51259));
    NOR2X1 U38388 (.A1(n17257), .A2(N4090), .ZN(N51260));
    INVX1 U38389 (.I(n35483), .ZN(N51261));
    NANDX1 U38390 (.A1(n36039), .A2(N7885), .ZN(N51262));
    NOR2X1 U38391 (.A1(n28380), .A2(n25336), .ZN(N51263));
    NOR2X1 U38392 (.A1(N4938), .A2(n19899), .ZN(n51264));
    NOR2X1 U38393 (.A1(n33219), .A2(n16305), .ZN(N51265));
    INVX1 U38394 (.I(n41886), .ZN(N51266));
    NOR2X1 U38395 (.A1(n20482), .A2(n25825), .ZN(N51267));
    NANDX1 U38396 (.A1(n32919), .A2(N6927), .ZN(N51268));
    INVX1 U38397 (.I(N1162), .ZN(N51269));
    NANDX1 U38398 (.A1(N4949), .A2(n29564), .ZN(N51270));
    INVX1 U38399 (.I(n29195), .ZN(N51271));
    NOR2X1 U38400 (.A1(n17249), .A2(n37992), .ZN(N51272));
    NANDX1 U38401 (.A1(n34080), .A2(n20238), .ZN(N51273));
    INVX1 U38402 (.I(n18274), .ZN(N51274));
    NANDX1 U38403 (.A1(N7937), .A2(N12755), .ZN(n51275));
    NOR2X1 U38404 (.A1(n17516), .A2(n38871), .ZN(N51276));
    INVX1 U38405 (.I(n23500), .ZN(N51277));
    NANDX1 U38406 (.A1(n31394), .A2(N1525), .ZN(N51278));
    INVX1 U38407 (.I(n13746), .ZN(N51279));
    NOR2X1 U38408 (.A1(n22961), .A2(n20673), .ZN(N51280));
    NANDX1 U38409 (.A1(n24122), .A2(n42274), .ZN(N51281));
    NOR2X1 U38410 (.A1(N10213), .A2(N11961), .ZN(N51282));
    INVX1 U38411 (.I(N3240), .ZN(N51283));
    NOR2X1 U38412 (.A1(N5764), .A2(n31750), .ZN(N51284));
    NOR2X1 U38413 (.A1(n26001), .A2(n14351), .ZN(N51285));
    INVX1 U38414 (.I(n31146), .ZN(N51286));
    INVX1 U38415 (.I(n30204), .ZN(N51287));
    NANDX1 U38416 (.A1(n29483), .A2(n25602), .ZN(N51288));
    NOR2X1 U38417 (.A1(N9510), .A2(n38635), .ZN(N51289));
    NOR2X1 U38418 (.A1(N11034), .A2(n28677), .ZN(N51290));
    NANDX1 U38419 (.A1(n20424), .A2(n41317), .ZN(N51291));
    NOR2X1 U38420 (.A1(N7845), .A2(n21967), .ZN(N51292));
    NOR2X1 U38421 (.A1(N10534), .A2(n21859), .ZN(n51293));
    INVX1 U38422 (.I(n21778), .ZN(N51294));
    NANDX1 U38423 (.A1(n31124), .A2(n27541), .ZN(N51295));
    INVX1 U38424 (.I(n30299), .ZN(N51296));
    INVX1 U38425 (.I(N7086), .ZN(N51297));
    INVX1 U38426 (.I(n20574), .ZN(N51298));
    INVX1 U38427 (.I(n34479), .ZN(N51299));
    INVX1 U38428 (.I(N5063), .ZN(N51300));
    INVX1 U38429 (.I(n18104), .ZN(N51301));
    INVX1 U38430 (.I(n34603), .ZN(N51302));
    NOR2X1 U38431 (.A1(N4965), .A2(N9487), .ZN(N51303));
    NOR2X1 U38432 (.A1(n15069), .A2(N7332), .ZN(N51304));
    NANDX1 U38433 (.A1(n22913), .A2(n18978), .ZN(N51305));
    INVX1 U38434 (.I(n23127), .ZN(N51306));
    NANDX1 U38435 (.A1(n29353), .A2(N1432), .ZN(n51307));
    INVX1 U38436 (.I(N6684), .ZN(N51308));
    NOR2X1 U38437 (.A1(n15197), .A2(n36983), .ZN(N51309));
    INVX1 U38438 (.I(N11963), .ZN(N51310));
    NANDX1 U38439 (.A1(n28654), .A2(n31015), .ZN(N51311));
    NOR2X1 U38440 (.A1(n26342), .A2(n25758), .ZN(N51312));
    NOR2X1 U38441 (.A1(N974), .A2(n19689), .ZN(N51313));
    NOR2X1 U38442 (.A1(n17093), .A2(n24654), .ZN(N51314));
    INVX1 U38443 (.I(N1502), .ZN(N51315));
    INVX1 U38444 (.I(N5219), .ZN(N51316));
    INVX1 U38445 (.I(N8842), .ZN(N51317));
    NOR2X1 U38446 (.A1(n14822), .A2(n31968), .ZN(N51318));
    NANDX1 U38447 (.A1(n33855), .A2(n23079), .ZN(N51319));
    NOR2X1 U38448 (.A1(n40538), .A2(n41730), .ZN(N51320));
    INVX1 U38449 (.I(n23728), .ZN(N51321));
    INVX1 U38450 (.I(n40219), .ZN(N51322));
    NOR2X1 U38451 (.A1(n24671), .A2(n17442), .ZN(n51323));
    NANDX1 U38452 (.A1(n40692), .A2(n43199), .ZN(N51324));
    NOR2X1 U38453 (.A1(n31345), .A2(n19415), .ZN(N51325));
    NOR2X1 U38454 (.A1(N4966), .A2(n33748), .ZN(N51326));
    INVX1 U38455 (.I(n39619), .ZN(N51327));
    NANDX1 U38456 (.A1(n21912), .A2(n37323), .ZN(N51328));
    NOR2X1 U38457 (.A1(n35787), .A2(n41825), .ZN(N51329));
    INVX1 U38458 (.I(N3554), .ZN(n51330));
    NOR2X1 U38459 (.A1(n29773), .A2(n16614), .ZN(N51331));
    INVX1 U38460 (.I(n17710), .ZN(N51332));
    NANDX1 U38461 (.A1(n42680), .A2(n13727), .ZN(N51333));
    NOR2X1 U38462 (.A1(N80), .A2(n28077), .ZN(N51334));
    NOR2X1 U38463 (.A1(n22896), .A2(n14977), .ZN(N51335));
    INVX1 U38464 (.I(n42982), .ZN(N51336));
    INVX1 U38465 (.I(N3766), .ZN(n51337));
    INVX1 U38466 (.I(n40966), .ZN(N51338));
    INVX1 U38467 (.I(n35010), .ZN(n51339));
    INVX1 U38468 (.I(N3398), .ZN(N51340));
    NANDX1 U38469 (.A1(n20643), .A2(n21596), .ZN(N51341));
    NANDX1 U38470 (.A1(n18995), .A2(n28290), .ZN(N51342));
    INVX1 U38471 (.I(n40881), .ZN(N51343));
    INVX1 U38472 (.I(n38442), .ZN(N51344));
    NOR2X1 U38473 (.A1(n21979), .A2(n29519), .ZN(N51345));
    NANDX1 U38474 (.A1(n35706), .A2(n17343), .ZN(N51346));
    INVX1 U38475 (.I(N9990), .ZN(N51347));
    INVX1 U38476 (.I(n28222), .ZN(N51348));
    NOR2X1 U38477 (.A1(N6959), .A2(n17411), .ZN(N51349));
    INVX1 U38478 (.I(N10725), .ZN(N51350));
    INVX1 U38479 (.I(n14988), .ZN(N51351));
    NANDX1 U38480 (.A1(N6624), .A2(n41780), .ZN(N51352));
    NANDX1 U38481 (.A1(N9752), .A2(N8631), .ZN(N51353));
    NANDX1 U38482 (.A1(n38347), .A2(n27625), .ZN(n51354));
    NANDX1 U38483 (.A1(n16703), .A2(n14714), .ZN(N51355));
    NOR2X1 U38484 (.A1(N11672), .A2(n31074), .ZN(n51356));
    NOR2X1 U38485 (.A1(n41191), .A2(n36321), .ZN(N51357));
    INVX1 U38486 (.I(N4741), .ZN(N51358));
    NOR2X1 U38487 (.A1(N12086), .A2(n17029), .ZN(N51359));
    NOR2X1 U38488 (.A1(n37051), .A2(n23987), .ZN(N51360));
    NANDX1 U38489 (.A1(N11073), .A2(n24391), .ZN(N51361));
    NANDX1 U38490 (.A1(n26061), .A2(N8516), .ZN(N51362));
    INVX1 U38491 (.I(n14048), .ZN(N51363));
    NOR2X1 U38492 (.A1(n21476), .A2(n22678), .ZN(N51364));
    NANDX1 U38493 (.A1(N6030), .A2(n39983), .ZN(N51365));
    INVX1 U38494 (.I(n22733), .ZN(N51366));
    NANDX1 U38495 (.A1(n20128), .A2(n34404), .ZN(N51367));
    INVX1 U38496 (.I(n29990), .ZN(N51368));
    NANDX1 U38497 (.A1(n24825), .A2(n32086), .ZN(N51369));
    NANDX1 U38498 (.A1(n22999), .A2(N699), .ZN(n51370));
    NANDX1 U38499 (.A1(n39075), .A2(n27429), .ZN(N51371));
    NOR2X1 U38500 (.A1(n29090), .A2(n38502), .ZN(N51372));
    NANDX1 U38501 (.A1(n34190), .A2(N10770), .ZN(n51373));
    NOR2X1 U38502 (.A1(N2442), .A2(n24817), .ZN(N51374));
    NANDX1 U38503 (.A1(n23917), .A2(n37175), .ZN(N51375));
    INVX1 U38504 (.I(n19626), .ZN(N51376));
    NOR2X1 U38505 (.A1(n38828), .A2(n42358), .ZN(N51377));
    INVX1 U38506 (.I(n15483), .ZN(N51378));
    NANDX1 U38507 (.A1(n33412), .A2(N2001), .ZN(N51379));
    NOR2X1 U38508 (.A1(n14764), .A2(n23766), .ZN(n51380));
    INVX1 U38509 (.I(n37762), .ZN(N51381));
    NOR2X1 U38510 (.A1(n27939), .A2(n23045), .ZN(N51382));
    NANDX1 U38511 (.A1(n41704), .A2(N8662), .ZN(N51383));
    INVX1 U38512 (.I(n26067), .ZN(N51384));
    NANDX1 U38513 (.A1(n37050), .A2(n18945), .ZN(N51385));
    NOR2X1 U38514 (.A1(N8075), .A2(n41014), .ZN(N51386));
    INVX1 U38515 (.I(N1777), .ZN(N51387));
    NOR2X1 U38516 (.A1(n24722), .A2(n25141), .ZN(N51388));
    INVX1 U38517 (.I(n13287), .ZN(N51389));
    INVX1 U38518 (.I(n14964), .ZN(N51390));
    INVX1 U38519 (.I(N6195), .ZN(n51391));
    INVX1 U38520 (.I(n37555), .ZN(N51392));
    INVX1 U38521 (.I(n30409), .ZN(n51393));
    INVX1 U38522 (.I(n38079), .ZN(N51394));
    INVX1 U38523 (.I(n39542), .ZN(N51395));
    INVX1 U38524 (.I(n42652), .ZN(N51396));
    NOR2X1 U38525 (.A1(n15992), .A2(n25460), .ZN(N51397));
    INVX1 U38526 (.I(N5051), .ZN(N51398));
    NANDX1 U38527 (.A1(N8351), .A2(n29702), .ZN(N51399));
    NANDX1 U38528 (.A1(N5892), .A2(n34798), .ZN(N51400));
    NANDX1 U38529 (.A1(N10018), .A2(N5727), .ZN(N51401));
    NANDX1 U38530 (.A1(N9499), .A2(n19013), .ZN(N51402));
    NOR2X1 U38531 (.A1(n24462), .A2(N11797), .ZN(N51403));
    NOR2X1 U38532 (.A1(n31106), .A2(N5879), .ZN(n51404));
    NOR2X1 U38533 (.A1(N7722), .A2(n17481), .ZN(N51405));
    NANDX1 U38534 (.A1(N8802), .A2(N3230), .ZN(N51406));
    INVX1 U38535 (.I(n41133), .ZN(N51407));
    INVX1 U38536 (.I(n30610), .ZN(N51408));
    NANDX1 U38537 (.A1(n20088), .A2(n35660), .ZN(N51409));
    INVX1 U38538 (.I(n28439), .ZN(N51410));
    INVX1 U38539 (.I(n17668), .ZN(N51411));
    NANDX1 U38540 (.A1(N2895), .A2(n15595), .ZN(N51412));
    NOR2X1 U38541 (.A1(n41773), .A2(N5510), .ZN(N51413));
    INVX1 U38542 (.I(n17313), .ZN(N51414));
    NANDX1 U38543 (.A1(N3875), .A2(n18789), .ZN(N51415));
    INVX1 U38544 (.I(n24660), .ZN(N51416));
    NOR2X1 U38545 (.A1(N5765), .A2(n32381), .ZN(N51417));
    INVX1 U38546 (.I(N2733), .ZN(N51418));
    NOR2X1 U38547 (.A1(n24737), .A2(n17351), .ZN(N51419));
    NANDX1 U38548 (.A1(N1627), .A2(n37640), .ZN(N51420));
    INVX1 U38549 (.I(N11394), .ZN(N51421));
    NOR2X1 U38550 (.A1(n31878), .A2(n29512), .ZN(N51422));
    NOR2X1 U38551 (.A1(N6074), .A2(N10050), .ZN(N51423));
    NANDX1 U38552 (.A1(n21668), .A2(n33756), .ZN(N51424));
    INVX1 U38553 (.I(n16858), .ZN(N51425));
    NANDX1 U38554 (.A1(n39263), .A2(N7897), .ZN(N51426));
    NANDX1 U38555 (.A1(N4260), .A2(N11301), .ZN(N51427));
    NANDX1 U38556 (.A1(n18606), .A2(N6745), .ZN(N51428));
    NOR2X1 U38557 (.A1(n40113), .A2(N9477), .ZN(n51429));
    NOR2X1 U38558 (.A1(N11058), .A2(n26827), .ZN(N51430));
    NANDX1 U38559 (.A1(N12684), .A2(N10675), .ZN(N51431));
    NANDX1 U38560 (.A1(n13757), .A2(n30182), .ZN(N51432));
    NANDX1 U38561 (.A1(n43269), .A2(n17786), .ZN(N51433));
    NANDX1 U38562 (.A1(n42998), .A2(n41436), .ZN(N51434));
    NOR2X1 U38563 (.A1(n33281), .A2(n19914), .ZN(N51435));
    NOR2X1 U38564 (.A1(n36129), .A2(N5384), .ZN(N51436));
    NOR2X1 U38565 (.A1(n42851), .A2(N9643), .ZN(N51437));
    INVX1 U38566 (.I(n30760), .ZN(N51438));
    INVX1 U38567 (.I(n31074), .ZN(N51439));
    NANDX1 U38568 (.A1(n14569), .A2(n30231), .ZN(N51440));
    NANDX1 U38569 (.A1(n25626), .A2(N3265), .ZN(N51441));
    NOR2X1 U38570 (.A1(n27989), .A2(n13939), .ZN(N51442));
    NOR2X1 U38571 (.A1(n41746), .A2(N648), .ZN(N51443));
    INVX1 U38572 (.I(n31222), .ZN(N51444));
    INVX1 U38573 (.I(n14842), .ZN(N51445));
    NANDX1 U38574 (.A1(n16396), .A2(n13437), .ZN(N51446));
    INVX1 U38575 (.I(n25989), .ZN(N51447));
    NOR2X1 U38576 (.A1(N2892), .A2(n31373), .ZN(N51448));
    NOR2X1 U38577 (.A1(N2270), .A2(n30695), .ZN(N51449));
    INVX1 U38578 (.I(n33030), .ZN(N51450));
    NANDX1 U38579 (.A1(n22889), .A2(n30287), .ZN(n51451));
    NOR2X1 U38580 (.A1(N9647), .A2(n35223), .ZN(N51452));
    INVX1 U38581 (.I(n12912), .ZN(N51453));
    NOR2X1 U38582 (.A1(n42374), .A2(n26850), .ZN(N51454));
    NOR2X1 U38583 (.A1(n30327), .A2(n27498), .ZN(N51455));
    NOR2X1 U38584 (.A1(n18076), .A2(n35610), .ZN(N51456));
    NOR2X1 U38585 (.A1(N5350), .A2(n41686), .ZN(N51457));
    NANDX1 U38586 (.A1(n15584), .A2(n13882), .ZN(N51458));
    NANDX1 U38587 (.A1(N8155), .A2(N1782), .ZN(N51459));
    INVX1 U38588 (.I(N10425), .ZN(N51460));
    NANDX1 U38589 (.A1(N5462), .A2(n33134), .ZN(N51461));
    INVX1 U38590 (.I(n28350), .ZN(n51462));
    NOR2X1 U38591 (.A1(n16066), .A2(n37997), .ZN(N51463));
    NOR2X1 U38592 (.A1(n30451), .A2(N7436), .ZN(N51464));
    NANDX1 U38593 (.A1(n29352), .A2(n23965), .ZN(N51465));
    NANDX1 U38594 (.A1(n16206), .A2(n41142), .ZN(N51466));
    NANDX1 U38595 (.A1(n23961), .A2(n22960), .ZN(N51467));
    NANDX1 U38596 (.A1(n29310), .A2(n21173), .ZN(N51468));
    INVX1 U38597 (.I(n34573), .ZN(N51469));
    NOR2X1 U38598 (.A1(n23156), .A2(n42728), .ZN(N51470));
    NOR2X1 U38599 (.A1(n26482), .A2(n42832), .ZN(N51471));
    NANDX1 U38600 (.A1(n31943), .A2(n32493), .ZN(n51472));
    NANDX1 U38601 (.A1(n16820), .A2(n42120), .ZN(N51473));
    INVX1 U38602 (.I(N1024), .ZN(N51474));
    NANDX1 U38603 (.A1(N4590), .A2(n41611), .ZN(N51475));
    INVX1 U38604 (.I(n33941), .ZN(N51476));
    NANDX1 U38605 (.A1(N3376), .A2(n39826), .ZN(N51477));
    NOR2X1 U38606 (.A1(n33698), .A2(N9994), .ZN(N51478));
    INVX1 U38607 (.I(n24382), .ZN(N51479));
    NOR2X1 U38608 (.A1(n43264), .A2(n22017), .ZN(N51480));
    NANDX1 U38609 (.A1(n34846), .A2(n34852), .ZN(N51481));
    NANDX1 U38610 (.A1(N7569), .A2(n17861), .ZN(N51482));
    NANDX1 U38611 (.A1(N2448), .A2(n39483), .ZN(N51483));
    NANDX1 U38612 (.A1(N3993), .A2(N12830), .ZN(N51484));
    NANDX1 U38613 (.A1(n21604), .A2(N3534), .ZN(N51485));
    INVX1 U38614 (.I(n15873), .ZN(N51486));
    NANDX1 U38615 (.A1(n34740), .A2(n39493), .ZN(N51487));
    INVX1 U38616 (.I(n27795), .ZN(N51488));
    INVX1 U38617 (.I(n22908), .ZN(N51489));
    NOR2X1 U38618 (.A1(N2367), .A2(N1527), .ZN(N51490));
    NOR2X1 U38619 (.A1(n31349), .A2(N1319), .ZN(N51491));
    NOR2X1 U38620 (.A1(N7960), .A2(n25844), .ZN(N51492));
    INVX1 U38621 (.I(n27297), .ZN(N51493));
    INVX1 U38622 (.I(n42696), .ZN(N51494));
    NANDX1 U38623 (.A1(n25539), .A2(n38706), .ZN(N51495));
    INVX1 U38624 (.I(n29531), .ZN(N51496));
    NOR2X1 U38625 (.A1(n39434), .A2(n40815), .ZN(N51497));
    NANDX1 U38626 (.A1(N4541), .A2(n13215), .ZN(n51498));
    INVX1 U38627 (.I(n28960), .ZN(N51499));
    INVX1 U38628 (.I(n39235), .ZN(N51500));
    NANDX1 U38629 (.A1(n34761), .A2(N8350), .ZN(n51501));
    INVX1 U38630 (.I(n26808), .ZN(N51502));
    NANDX1 U38631 (.A1(n19911), .A2(N4364), .ZN(n51503));
    NANDX1 U38632 (.A1(N9895), .A2(N2003), .ZN(N51504));
    NANDX1 U38633 (.A1(N1579), .A2(n29300), .ZN(N51505));
    NOR2X1 U38634 (.A1(n33954), .A2(n21501), .ZN(N51506));
    NOR2X1 U38635 (.A1(n29188), .A2(n21418), .ZN(N51507));
    INVX1 U38636 (.I(n16611), .ZN(N51508));
    NANDX1 U38637 (.A1(n38107), .A2(N7567), .ZN(N51509));
    NOR2X1 U38638 (.A1(n41001), .A2(N194), .ZN(N51510));
    NANDX1 U38639 (.A1(n39916), .A2(n39428), .ZN(N51511));
    INVX1 U38640 (.I(n20885), .ZN(N51512));
    NOR2X1 U38641 (.A1(n31351), .A2(n37372), .ZN(N51513));
    NANDX1 U38642 (.A1(n40941), .A2(n41735), .ZN(N51514));
    INVX1 U38643 (.I(n40515), .ZN(N51515));
    INVX1 U38644 (.I(n21131), .ZN(n51516));
    NANDX1 U38645 (.A1(n19245), .A2(n17146), .ZN(N51517));
    INVX1 U38646 (.I(n40745), .ZN(N51518));
    NOR2X1 U38647 (.A1(N7970), .A2(n18690), .ZN(N51519));
    NOR2X1 U38648 (.A1(n14260), .A2(n15429), .ZN(N51520));
    NANDX1 U38649 (.A1(n21826), .A2(n27028), .ZN(n51521));
    NANDX1 U38650 (.A1(N11699), .A2(n13794), .ZN(N51522));
    NANDX1 U38651 (.A1(N7655), .A2(n13843), .ZN(N51523));
    NOR2X1 U38652 (.A1(n34791), .A2(n34873), .ZN(N51524));
    NOR2X1 U38653 (.A1(n38651), .A2(n22021), .ZN(N51525));
    INVX1 U38654 (.I(n33065), .ZN(N51526));
    INVX1 U38655 (.I(n40100), .ZN(N51527));
    NANDX1 U38656 (.A1(n17684), .A2(n15872), .ZN(N51528));
    INVX1 U38657 (.I(n29618), .ZN(N51529));
    NOR2X1 U38658 (.A1(N2455), .A2(n27267), .ZN(N51530));
    INVX1 U38659 (.I(n28126), .ZN(N51531));
    NOR2X1 U38660 (.A1(n36942), .A2(N4959), .ZN(n51532));
    NOR2X1 U38661 (.A1(N10177), .A2(N12473), .ZN(N51533));
    NOR2X1 U38662 (.A1(n23970), .A2(n16430), .ZN(N51534));
    NOR2X1 U38663 (.A1(n27492), .A2(n30951), .ZN(n51535));
    NOR2X1 U38664 (.A1(n18892), .A2(n39371), .ZN(n51536));
    INVX1 U38665 (.I(n40912), .ZN(N51537));
    NOR2X1 U38666 (.A1(n27832), .A2(n16503), .ZN(N51538));
    NOR2X1 U38667 (.A1(n28234), .A2(n23866), .ZN(N51539));
    INVX1 U38668 (.I(n35462), .ZN(n51540));
    NANDX1 U38669 (.A1(N7584), .A2(n27596), .ZN(N51541));
    NOR2X1 U38670 (.A1(n29097), .A2(N12250), .ZN(N51542));
    NANDX1 U38671 (.A1(N12246), .A2(n17208), .ZN(N51543));
    NANDX1 U38672 (.A1(n22422), .A2(n19360), .ZN(N51544));
    NANDX1 U38673 (.A1(n36071), .A2(n35789), .ZN(N51545));
    NANDX1 U38674 (.A1(n20091), .A2(n12947), .ZN(N51546));
    NANDX1 U38675 (.A1(n38982), .A2(n41997), .ZN(N51547));
    NANDX1 U38676 (.A1(n26102), .A2(n34258), .ZN(N51548));
    NANDX1 U38677 (.A1(n42604), .A2(n23146), .ZN(n51549));
    NOR2X1 U38678 (.A1(N12677), .A2(n27905), .ZN(N51550));
    NOR2X1 U38679 (.A1(N12367), .A2(n25168), .ZN(N51551));
    INVX1 U38680 (.I(N6171), .ZN(N51552));
    INVX1 U38681 (.I(n36574), .ZN(N51553));
    NANDX1 U38682 (.A1(N12717), .A2(N10309), .ZN(N51554));
    INVX1 U38683 (.I(n24818), .ZN(N51555));
    NANDX1 U38684 (.A1(N1474), .A2(n17417), .ZN(N51556));
    NOR2X1 U38685 (.A1(n42736), .A2(n37507), .ZN(N51557));
    INVX1 U38686 (.I(n17283), .ZN(N51558));
    INVX1 U38687 (.I(N12816), .ZN(N51559));
    NANDX1 U38688 (.A1(n38477), .A2(N3601), .ZN(N51560));
    INVX1 U38689 (.I(n27288), .ZN(N51561));
    NANDX1 U38690 (.A1(N9123), .A2(n39964), .ZN(N51562));
    INVX1 U38691 (.I(N5852), .ZN(N51563));
    INVX1 U38692 (.I(n26026), .ZN(N51564));
    NANDX1 U38693 (.A1(N4708), .A2(n26498), .ZN(N51565));
    INVX1 U38694 (.I(n25567), .ZN(N51566));
    NANDX1 U38695 (.A1(n23265), .A2(N4369), .ZN(N51567));
    NANDX1 U38696 (.A1(n42613), .A2(n38995), .ZN(N51568));
    NOR2X1 U38697 (.A1(N486), .A2(n38258), .ZN(N51569));
    INVX1 U38698 (.I(N4457), .ZN(N51570));
    NANDX1 U38699 (.A1(n23745), .A2(n17272), .ZN(n51571));
    NOR2X1 U38700 (.A1(n18750), .A2(N10553), .ZN(N51572));
    INVX1 U38701 (.I(n35717), .ZN(N51573));
    INVX1 U38702 (.I(n24683), .ZN(N51574));
    INVX1 U38703 (.I(n27836), .ZN(N51575));
    INVX1 U38704 (.I(n30746), .ZN(N51576));
    NANDX1 U38705 (.A1(N6917), .A2(n25134), .ZN(N51577));
    NOR2X1 U38706 (.A1(n19873), .A2(n40380), .ZN(N51578));
    INVX1 U38707 (.I(n43138), .ZN(N51579));
    NOR2X1 U38708 (.A1(N11907), .A2(n31958), .ZN(N51580));
    NOR2X1 U38709 (.A1(n39562), .A2(n32443), .ZN(N51581));
    NANDX1 U38710 (.A1(n40611), .A2(n26579), .ZN(N51582));
    NOR2X1 U38711 (.A1(n20884), .A2(N379), .ZN(N51583));
    NOR2X1 U38712 (.A1(n29313), .A2(N611), .ZN(N51584));
    NOR2X1 U38713 (.A1(n21557), .A2(n27588), .ZN(n51585));
    INVX1 U38714 (.I(n43445), .ZN(N51586));
    NANDX1 U38715 (.A1(n21493), .A2(n20399), .ZN(N51587));
    INVX1 U38716 (.I(n28410), .ZN(N51588));
    INVX1 U38717 (.I(n17074), .ZN(N51589));
    NOR2X1 U38718 (.A1(n20558), .A2(n25531), .ZN(N51590));
    NOR2X1 U38719 (.A1(n45401), .A2(N1793), .ZN(N51591));
    NANDX1 U38720 (.A1(N7542), .A2(N4083), .ZN(N51592));
    INVX1 U38721 (.I(n24693), .ZN(N51593));
    NOR2X1 U38722 (.A1(n48976), .A2(n21944), .ZN(N51594));
    NANDX1 U38723 (.A1(N1661), .A2(n23292), .ZN(N51595));
    NANDX1 U38724 (.A1(n40901), .A2(n17680), .ZN(N51596));
    NANDX1 U38725 (.A1(n37484), .A2(N11173), .ZN(N51597));
    INVX1 U38726 (.I(n43561), .ZN(N51598));
    INVX1 U38727 (.I(n34936), .ZN(N51599));
    NANDX1 U38728 (.A1(N4274), .A2(N8614), .ZN(N51600));
    NANDX1 U38729 (.A1(n26812), .A2(n29172), .ZN(N51601));
    INVX1 U38730 (.I(n35195), .ZN(N51602));
    INVX1 U38731 (.I(N7814), .ZN(N51603));
    NOR2X1 U38732 (.A1(N553), .A2(n33512), .ZN(N51604));
    INVX1 U38733 (.I(n46861), .ZN(N51605));
    INVX1 U38734 (.I(N11583), .ZN(N51606));
    NANDX1 U38735 (.A1(n20984), .A2(n13243), .ZN(N51607));
    INVX1 U38736 (.I(n39597), .ZN(N51608));
    NANDX1 U38737 (.A1(n28215), .A2(N8154), .ZN(N51609));
    NANDX1 U38738 (.A1(n39387), .A2(n47637), .ZN(N51610));
    NOR2X1 U38739 (.A1(n22945), .A2(n30985), .ZN(n51611));
    INVX1 U38740 (.I(n48834), .ZN(N51612));
    INVX1 U38741 (.I(n49122), .ZN(N51613));
    NOR2X1 U38742 (.A1(n38797), .A2(N3555), .ZN(N51614));
    NANDX1 U38743 (.A1(N10192), .A2(n32984), .ZN(N51615));
    NOR2X1 U38744 (.A1(N10745), .A2(n14908), .ZN(N51616));
    NOR2X1 U38745 (.A1(N6017), .A2(N5860), .ZN(N51617));
    NANDX1 U38746 (.A1(n44849), .A2(n48460), .ZN(N51618));
    NOR2X1 U38747 (.A1(N3795), .A2(N6496), .ZN(N51619));
    NANDX1 U38748 (.A1(n32009), .A2(n14649), .ZN(N51620));
    NOR2X1 U38749 (.A1(n41423), .A2(N10698), .ZN(N51621));
    NANDX1 U38750 (.A1(n34395), .A2(N11710), .ZN(N51622));
    NOR2X1 U38751 (.A1(n31640), .A2(n51307), .ZN(N51623));
    NOR2X1 U38752 (.A1(n25725), .A2(n38516), .ZN(N51624));
    INVX1 U38753 (.I(N3415), .ZN(N51625));
    NOR2X1 U38754 (.A1(n33989), .A2(N912), .ZN(N51626));
    INVX1 U38755 (.I(n48896), .ZN(N51627));
    INVX1 U38756 (.I(N5524), .ZN(N51628));
    INVX1 U38757 (.I(n35877), .ZN(N51629));
    NOR2X1 U38758 (.A1(n43271), .A2(n20805), .ZN(N51630));
    NANDX1 U38759 (.A1(n49766), .A2(n29903), .ZN(N51631));
    NANDX1 U38760 (.A1(n34443), .A2(n49067), .ZN(N51632));
    NOR2X1 U38761 (.A1(n45140), .A2(n40297), .ZN(N51633));
    INVX1 U38762 (.I(N5261), .ZN(N51634));
    NOR2X1 U38763 (.A1(n22155), .A2(n26595), .ZN(N51635));
    NOR2X1 U38764 (.A1(n47879), .A2(n35138), .ZN(N51636));
    NOR2X1 U38765 (.A1(n21322), .A2(N2285), .ZN(N51637));
    NANDX1 U38766 (.A1(n22233), .A2(N1791), .ZN(N51638));
    INVX1 U38767 (.I(N4864), .ZN(N51639));
    INVX1 U38768 (.I(n43160), .ZN(N51640));
    INVX1 U38769 (.I(n49329), .ZN(N51641));
    INVX1 U38770 (.I(N9957), .ZN(N51642));
    NANDX1 U38771 (.A1(N3048), .A2(n39859), .ZN(N51643));
    NOR2X1 U38772 (.A1(N7518), .A2(n37337), .ZN(N51644));
    NOR2X1 U38773 (.A1(n22685), .A2(n47661), .ZN(N51645));
    INVX1 U38774 (.I(n49561), .ZN(N51646));
    NANDX1 U38775 (.A1(n46927), .A2(n24567), .ZN(N51647));
    NANDX1 U38776 (.A1(n43217), .A2(n29733), .ZN(N51648));
    NANDX1 U38777 (.A1(n12950), .A2(N2045), .ZN(N51649));
    INVX1 U38778 (.I(N5211), .ZN(N51650));
    INVX1 U38779 (.I(N751), .ZN(N51651));
    NOR2X1 U38780 (.A1(N2793), .A2(n13939), .ZN(N51652));
    INVX1 U38781 (.I(N533), .ZN(N51653));
    INVX1 U38782 (.I(n30798), .ZN(N51654));
    INVX1 U38783 (.I(n43471), .ZN(N51655));
    INVX1 U38784 (.I(N10687), .ZN(N51656));
    NOR2X1 U38785 (.A1(n48048), .A2(n44944), .ZN(N51657));
    INVX1 U38786 (.I(n44120), .ZN(N51658));
    NANDX1 U38787 (.A1(n20056), .A2(N7201), .ZN(N51659));
    NANDX1 U38788 (.A1(n14651), .A2(n16302), .ZN(N51660));
    NANDX1 U38789 (.A1(n44383), .A2(n20839), .ZN(N51661));
    INVX1 U38790 (.I(n16455), .ZN(N51662));
    INVX1 U38791 (.I(N6541), .ZN(N51663));
    NOR2X1 U38792 (.A1(n47195), .A2(n38231), .ZN(N51664));
    NANDX1 U38793 (.A1(n31161), .A2(N7484), .ZN(N51665));
    NANDX1 U38794 (.A1(n19997), .A2(n38282), .ZN(N51666));
    NANDX1 U38795 (.A1(N11879), .A2(n48993), .ZN(N51667));
    NOR2X1 U38796 (.A1(n32895), .A2(n45453), .ZN(N51668));
    INVX1 U38797 (.I(N3390), .ZN(N51669));
    NANDX1 U38798 (.A1(n51536), .A2(n45062), .ZN(N51670));
    NOR2X1 U38799 (.A1(N5057), .A2(n29740), .ZN(N51671));
    NANDX1 U38800 (.A1(n23410), .A2(n22534), .ZN(N51672));
    NOR2X1 U38801 (.A1(N3124), .A2(n38988), .ZN(N51673));
    INVX1 U38802 (.I(n31281), .ZN(N51674));
    NOR2X1 U38803 (.A1(N12842), .A2(n17923), .ZN(N51675));
    NOR2X1 U38804 (.A1(n14031), .A2(n25406), .ZN(N51676));
    NANDX1 U38805 (.A1(n34027), .A2(n33715), .ZN(N51677));
    NOR2X1 U38806 (.A1(n15933), .A2(n31120), .ZN(N51678));
    NANDX1 U38807 (.A1(n48827), .A2(n46600), .ZN(N51679));
    NOR2X1 U38808 (.A1(n22245), .A2(N3023), .ZN(N51680));
    NANDX1 U38809 (.A1(n15718), .A2(n18235), .ZN(N51681));
    INVX1 U38810 (.I(n45457), .ZN(N51682));
    NOR2X1 U38811 (.A1(N889), .A2(n38018), .ZN(N51683));
    NANDX1 U38812 (.A1(N4012), .A2(n47033), .ZN(N51684));
    NANDX1 U38813 (.A1(n35292), .A2(n46364), .ZN(N51685));
    NANDX1 U38814 (.A1(n23242), .A2(n38804), .ZN(N51686));
    INVX1 U38815 (.I(n48648), .ZN(N51687));
    NOR2X1 U38816 (.A1(N8756), .A2(N802), .ZN(N51688));
    NOR2X1 U38817 (.A1(n24688), .A2(n31921), .ZN(N51689));
    NANDX1 U38818 (.A1(n43543), .A2(n48548), .ZN(N51690));
    NANDX1 U38819 (.A1(n14199), .A2(n51571), .ZN(N51691));
    INVX1 U38820 (.I(n51532), .ZN(N51692));
    NANDX1 U38821 (.A1(n43282), .A2(n45400), .ZN(N51693));
    NANDX1 U38822 (.A1(n44170), .A2(N1857), .ZN(N51694));
    INVX1 U38823 (.I(n18209), .ZN(N51695));
    NANDX1 U38824 (.A1(n49621), .A2(n23529), .ZN(N51696));
    NOR2X1 U38825 (.A1(n40292), .A2(n46770), .ZN(N51697));
    NANDX1 U38826 (.A1(n15021), .A2(n13857), .ZN(N51698));
    NANDX1 U38827 (.A1(n45392), .A2(n14659), .ZN(N51699));
    NANDX1 U38828 (.A1(n18491), .A2(n16607), .ZN(N51700));
    INVX1 U38829 (.I(N10445), .ZN(N51701));
    INVX1 U38830 (.I(n14112), .ZN(N51702));
    NANDX1 U38831 (.A1(n35165), .A2(n28326), .ZN(N51703));
    NANDX1 U38832 (.A1(n23409), .A2(n41635), .ZN(N51704));
    NOR2X1 U38833 (.A1(N1457), .A2(N4244), .ZN(N51705));
    NANDX1 U38834 (.A1(n43276), .A2(n44068), .ZN(N51706));
    INVX1 U38835 (.I(n41308), .ZN(N51707));
    NOR2X1 U38836 (.A1(n14533), .A2(N39), .ZN(N51708));
    INVX1 U38837 (.I(n37056), .ZN(N51709));
    NANDX1 U38838 (.A1(n16690), .A2(N2903), .ZN(N51710));
    INVX1 U38839 (.I(n31348), .ZN(N51711));
    INVX1 U38840 (.I(n48968), .ZN(N51712));
    INVX1 U38841 (.I(n19732), .ZN(N51713));
    NANDX1 U38842 (.A1(n31549), .A2(N3871), .ZN(N51714));
    NOR2X1 U38843 (.A1(n15125), .A2(n32196), .ZN(N51715));
    NOR2X1 U38844 (.A1(N8561), .A2(n43858), .ZN(N51716));
    NANDX1 U38845 (.A1(n31634), .A2(n48101), .ZN(N51717));
    NANDX1 U38846 (.A1(n44937), .A2(n40580), .ZN(N51718));
    NANDX1 U38847 (.A1(n34656), .A2(n26616), .ZN(N51719));
    NOR2X1 U38848 (.A1(N4722), .A2(n29449), .ZN(N51720));
    NOR2X1 U38849 (.A1(n41396), .A2(n46138), .ZN(N51721));
    NANDX1 U38850 (.A1(n20285), .A2(n47514), .ZN(N51722));
    NANDX1 U38851 (.A1(n39280), .A2(n13908), .ZN(N51723));
    NOR2X1 U38852 (.A1(n17132), .A2(n15484), .ZN(N51724));
    NOR2X1 U38853 (.A1(N11271), .A2(N636), .ZN(N51725));
    NOR2X1 U38854 (.A1(n21639), .A2(n30812), .ZN(N51726));
    INVX1 U38855 (.I(n20431), .ZN(N51727));
    NOR2X1 U38856 (.A1(n51380), .A2(N1148), .ZN(N51728));
    NOR2X1 U38857 (.A1(N10399), .A2(N4322), .ZN(N51729));
    NANDX1 U38858 (.A1(N7042), .A2(n22027), .ZN(N51730));
    NANDX1 U38859 (.A1(N6518), .A2(n16844), .ZN(N51731));
    NOR2X1 U38860 (.A1(N1068), .A2(n44535), .ZN(N51732));
    INVX1 U38861 (.I(n18609), .ZN(N51733));
    NANDX1 U38862 (.A1(n33008), .A2(n32516), .ZN(n51734));
    INVX1 U38863 (.I(n20167), .ZN(N51735));
    NOR2X1 U38864 (.A1(N193), .A2(n31437), .ZN(N51736));
    NANDX1 U38865 (.A1(n41175), .A2(N1487), .ZN(N51737));
    NOR2X1 U38866 (.A1(n44454), .A2(n43534), .ZN(N51738));
    INVX1 U38867 (.I(n14273), .ZN(N51739));
    NOR2X1 U38868 (.A1(N4590), .A2(n46287), .ZN(N51740));
    INVX1 U38869 (.I(n35094), .ZN(N51741));
    INVX1 U38870 (.I(N11085), .ZN(N51742));
    INVX1 U38871 (.I(N8258), .ZN(N51743));
    NANDX1 U38872 (.A1(n43762), .A2(n30941), .ZN(n51744));
    INVX1 U38873 (.I(n37489), .ZN(N51745));
    INVX1 U38874 (.I(n50594), .ZN(N51746));
    NANDX1 U38875 (.A1(N504), .A2(N12027), .ZN(N51747));
    NOR2X1 U38876 (.A1(n18530), .A2(N12219), .ZN(N51748));
    NOR2X1 U38877 (.A1(n37191), .A2(n23421), .ZN(N51749));
    NOR2X1 U38878 (.A1(N5104), .A2(n37902), .ZN(N51750));
    NOR2X1 U38879 (.A1(n35461), .A2(N586), .ZN(N51751));
    NOR2X1 U38880 (.A1(n40050), .A2(n16900), .ZN(N51752));
    NANDX1 U38881 (.A1(n23555), .A2(n40256), .ZN(n51753));
    NANDX1 U38882 (.A1(n42285), .A2(n48514), .ZN(N51754));
    NOR2X1 U38883 (.A1(N4486), .A2(n49482), .ZN(N51755));
    NOR2X1 U38884 (.A1(n41974), .A2(n17471), .ZN(N51756));
    NANDX1 U38885 (.A1(n30910), .A2(n39590), .ZN(N51757));
    INVX1 U38886 (.I(n18396), .ZN(N51758));
    NANDX1 U38887 (.A1(n14242), .A2(n28962), .ZN(N51759));
    NANDX1 U38888 (.A1(n37662), .A2(n41015), .ZN(N51760));
    NANDX1 U38889 (.A1(n45591), .A2(n15041), .ZN(N51761));
    NANDX1 U38890 (.A1(n16204), .A2(N3776), .ZN(N51762));
    NOR2X1 U38891 (.A1(n33103), .A2(N3184), .ZN(N51763));
    INVX1 U38892 (.I(n21771), .ZN(N51764));
    NANDX1 U38893 (.A1(n18697), .A2(n40312), .ZN(N51765));
    INVX1 U38894 (.I(n23182), .ZN(N51766));
    INVX1 U38895 (.I(n43087), .ZN(N51767));
    NOR2X1 U38896 (.A1(n25703), .A2(N11468), .ZN(N51768));
    NOR2X1 U38897 (.A1(n13705), .A2(n13491), .ZN(N51769));
    NOR2X1 U38898 (.A1(N11880), .A2(n27732), .ZN(N51770));
    NANDX1 U38899 (.A1(n47245), .A2(n35421), .ZN(N51771));
    NANDX1 U38900 (.A1(n36126), .A2(n29423), .ZN(N51772));
    NOR2X1 U38901 (.A1(n30494), .A2(n45626), .ZN(N51773));
    NANDX1 U38902 (.A1(n13324), .A2(n27140), .ZN(N51774));
    NANDX1 U38903 (.A1(n19709), .A2(n18938), .ZN(N51775));
    INVX1 U38904 (.I(N8433), .ZN(N51776));
    NANDX1 U38905 (.A1(n40783), .A2(N1643), .ZN(N51777));
    INVX1 U38906 (.I(n32281), .ZN(N51778));
    INVX1 U38907 (.I(N11624), .ZN(N51779));
    NOR2X1 U38908 (.A1(n51330), .A2(n46944), .ZN(N51780));
    NANDX1 U38909 (.A1(n24285), .A2(N7235), .ZN(N51781));
    NANDX1 U38910 (.A1(N4585), .A2(N2892), .ZN(N51782));
    INVX1 U38911 (.I(n47516), .ZN(N51783));
    NOR2X1 U38912 (.A1(N8307), .A2(n23928), .ZN(N51784));
    INVX1 U38913 (.I(N2344), .ZN(N51785));
    NANDX1 U38914 (.A1(N1274), .A2(n51100), .ZN(N51786));
    NANDX1 U38915 (.A1(n42598), .A2(n40065), .ZN(N51787));
    NANDX1 U38916 (.A1(n21058), .A2(n17754), .ZN(N51788));
    INVX1 U38917 (.I(n22700), .ZN(N51789));
    NOR2X1 U38918 (.A1(N10907), .A2(N7937), .ZN(N51790));
    INVX1 U38919 (.I(n24683), .ZN(N51791));
    NANDX1 U38920 (.A1(n32270), .A2(n21976), .ZN(N51792));
    INVX1 U38921 (.I(n39504), .ZN(N51793));
    NOR2X1 U38922 (.A1(n28191), .A2(N12423), .ZN(N51794));
    INVX1 U38923 (.I(n45734), .ZN(N51795));
    NANDX1 U38924 (.A1(n34192), .A2(n18073), .ZN(N51796));
    NOR2X1 U38925 (.A1(N6563), .A2(n43803), .ZN(N51797));
    NANDX1 U38926 (.A1(N6074), .A2(n44546), .ZN(N51798));
    NANDX1 U38927 (.A1(n16167), .A2(n42333), .ZN(N51799));
    NANDX1 U38928 (.A1(n33920), .A2(n50931), .ZN(N51800));
    NANDX1 U38929 (.A1(n37594), .A2(n31866), .ZN(N51801));
    INVX1 U38930 (.I(n22919), .ZN(N51802));
    INVX1 U38931 (.I(n44358), .ZN(N51803));
    NOR2X1 U38932 (.A1(n26935), .A2(n16375), .ZN(N51804));
    NOR2X1 U38933 (.A1(n43963), .A2(n44565), .ZN(N51805));
    NOR2X1 U38934 (.A1(n18260), .A2(N8739), .ZN(N51806));
    NANDX1 U38935 (.A1(n22479), .A2(n26811), .ZN(N51807));
    NANDX1 U38936 (.A1(n29041), .A2(n40641), .ZN(N51808));
    NOR2X1 U38937 (.A1(N5143), .A2(n33598), .ZN(N51809));
    NANDX1 U38938 (.A1(n21309), .A2(n45959), .ZN(N51810));
    INVX1 U38939 (.I(N3640), .ZN(N51811));
    NANDX1 U38940 (.A1(n22050), .A2(n41233), .ZN(N51812));
    INVX1 U38941 (.I(n37114), .ZN(N51813));
    NANDX1 U38942 (.A1(N565), .A2(n29883), .ZN(N51814));
    NANDX1 U38943 (.A1(n49116), .A2(n16285), .ZN(N51815));
    NANDX1 U38944 (.A1(N11518), .A2(n30878), .ZN(N51816));
    INVX1 U38945 (.I(n51393), .ZN(N51817));
    INVX1 U38946 (.I(n20307), .ZN(N51818));
    NANDX1 U38947 (.A1(n36454), .A2(n46771), .ZN(N51819));
    NOR2X1 U38948 (.A1(n25507), .A2(n23980), .ZN(N51820));
    NOR2X1 U38949 (.A1(n29132), .A2(n46119), .ZN(N51821));
    NANDX1 U38950 (.A1(n23502), .A2(n31070), .ZN(N51822));
    NOR2X1 U38951 (.A1(n38831), .A2(N1531), .ZN(N51823));
    NOR2X1 U38952 (.A1(N4464), .A2(n38644), .ZN(N51824));
    NANDX1 U38953 (.A1(n26645), .A2(n38554), .ZN(N51825));
    INVX1 U38954 (.I(n45788), .ZN(N51826));
    NANDX1 U38955 (.A1(n39158), .A2(N5717), .ZN(N51827));
    INVX1 U38956 (.I(N12445), .ZN(N51828));
    NANDX1 U38957 (.A1(n43771), .A2(n32751), .ZN(N51829));
    NOR2X1 U38958 (.A1(n28636), .A2(n27934), .ZN(N51830));
    NOR2X1 U38959 (.A1(n24170), .A2(n21941), .ZN(N51831));
    NANDX1 U38960 (.A1(n23330), .A2(n16472), .ZN(N51832));
    INVX1 U38961 (.I(n46831), .ZN(N51833));
    NOR2X1 U38962 (.A1(n50097), .A2(N4101), .ZN(N51834));
    INVX1 U38963 (.I(N9621), .ZN(N51835));
    INVX1 U38964 (.I(N6155), .ZN(N51836));
    NANDX1 U38965 (.A1(N5237), .A2(n44708), .ZN(N51837));
    NANDX1 U38966 (.A1(n51024), .A2(n17986), .ZN(N51838));
    NANDX1 U38967 (.A1(N5152), .A2(n22141), .ZN(N51839));
    NANDX1 U38968 (.A1(n32289), .A2(n35939), .ZN(N51840));
    NANDX1 U38969 (.A1(N8505), .A2(n12987), .ZN(N51841));
    NANDX1 U38970 (.A1(n27687), .A2(N7184), .ZN(N51842));
    NANDX1 U38971 (.A1(N159), .A2(n30513), .ZN(n51843));
    INVX1 U38972 (.I(n20431), .ZN(N51844));
    NANDX1 U38973 (.A1(n18333), .A2(n18940), .ZN(N51845));
    NANDX1 U38974 (.A1(N7459), .A2(n50176), .ZN(N51846));
    NANDX1 U38975 (.A1(n13613), .A2(N1911), .ZN(N51847));
    NOR2X1 U38976 (.A1(n28349), .A2(n15099), .ZN(N51848));
    NOR2X1 U38977 (.A1(n46334), .A2(n15856), .ZN(N51849));
    INVX1 U38978 (.I(n16887), .ZN(N51850));
    NOR2X1 U38979 (.A1(n33847), .A2(n22853), .ZN(N51851));
    INVX1 U38980 (.I(N12379), .ZN(N51852));
    INVX1 U38981 (.I(n29005), .ZN(N51853));
    INVX1 U38982 (.I(n13051), .ZN(N51854));
    NANDX1 U38983 (.A1(n40224), .A2(n13591), .ZN(N51855));
    NANDX1 U38984 (.A1(N9066), .A2(n30990), .ZN(N51856));
    NANDX1 U38985 (.A1(n49621), .A2(n22518), .ZN(N51857));
    NANDX1 U38986 (.A1(n48209), .A2(n22609), .ZN(N51858));
    NANDX1 U38987 (.A1(n20147), .A2(n49553), .ZN(N51859));
    NOR2X1 U38988 (.A1(n35245), .A2(n45959), .ZN(N51860));
    NANDX1 U38989 (.A1(n51100), .A2(n25901), .ZN(N51861));
    NANDX1 U38990 (.A1(n50184), .A2(N8160), .ZN(N51862));
    INVX1 U38991 (.I(n35276), .ZN(N51863));
    NOR2X1 U38992 (.A1(N2275), .A2(N12692), .ZN(N51864));
    INVX1 U38993 (.I(n36941), .ZN(N51865));
    INVX1 U38994 (.I(n40882), .ZN(n51866));
    INVX1 U38995 (.I(N1722), .ZN(N51867));
    INVX1 U38996 (.I(n51549), .ZN(N51868));
    INVX1 U38997 (.I(n18008), .ZN(N51869));
    NANDX1 U38998 (.A1(n27282), .A2(n36244), .ZN(N51870));
    INVX1 U38999 (.I(N12446), .ZN(N51871));
    NOR2X1 U39000 (.A1(n34695), .A2(N4342), .ZN(N51872));
    NOR2X1 U39001 (.A1(n29065), .A2(N12600), .ZN(N51873));
    NANDX1 U39002 (.A1(n24994), .A2(N7771), .ZN(N51874));
    NANDX1 U39003 (.A1(N3181), .A2(n25795), .ZN(N51875));
    NOR2X1 U39004 (.A1(n45334), .A2(n49686), .ZN(N51876));
    NANDX1 U39005 (.A1(n24377), .A2(N5066), .ZN(N51877));
    NOR2X1 U39006 (.A1(n13670), .A2(n25625), .ZN(N51878));
    NANDX1 U39007 (.A1(n33645), .A2(n25586), .ZN(N51879));
    NOR2X1 U39008 (.A1(N65), .A2(n18091), .ZN(N51880));
    INVX1 U39009 (.I(N6336), .ZN(N51881));
    NANDX1 U39010 (.A1(n21098), .A2(N11138), .ZN(N51882));
    INVX1 U39011 (.I(n25440), .ZN(N51883));
    NOR2X1 U39012 (.A1(n15404), .A2(N8067), .ZN(N51884));
    INVX1 U39013 (.I(N10425), .ZN(N51885));
    NOR2X1 U39014 (.A1(n30624), .A2(n13605), .ZN(N51886));
    NANDX1 U39015 (.A1(n14137), .A2(n28966), .ZN(N51887));
    NANDX1 U39016 (.A1(N10340), .A2(N1754), .ZN(N51888));
    NOR2X1 U39017 (.A1(n24176), .A2(n37040), .ZN(N51889));
    NANDX1 U39018 (.A1(N9760), .A2(n19096), .ZN(N51890));
    INVX1 U39019 (.I(n21103), .ZN(N51891));
    NOR2X1 U39020 (.A1(n45794), .A2(n29755), .ZN(N51892));
    INVX1 U39021 (.I(n49027), .ZN(N51893));
    NOR2X1 U39022 (.A1(n49893), .A2(n35365), .ZN(N51894));
    NANDX1 U39023 (.A1(n19517), .A2(n20796), .ZN(n51895));
    NANDX1 U39024 (.A1(n20343), .A2(N1248), .ZN(N51896));
    NOR2X1 U39025 (.A1(n50967), .A2(n14852), .ZN(N51897));
    INVX1 U39026 (.I(n13515), .ZN(N51898));
    NOR2X1 U39027 (.A1(N1721), .A2(n45470), .ZN(N51899));
    NANDX1 U39028 (.A1(n38158), .A2(n39673), .ZN(N51900));
    INVX1 U39029 (.I(n18660), .ZN(N51901));
    NANDX1 U39030 (.A1(n41762), .A2(n46363), .ZN(N51902));
    NOR2X1 U39031 (.A1(N977), .A2(n40569), .ZN(N51903));
    INVX1 U39032 (.I(n39732), .ZN(N51904));
    NOR2X1 U39033 (.A1(N9636), .A2(n38037), .ZN(N51905));
    INVX1 U39034 (.I(n25983), .ZN(N51906));
    NANDX1 U39035 (.A1(N12607), .A2(n50395), .ZN(N51907));
    NANDX1 U39036 (.A1(n13854), .A2(n30700), .ZN(N51908));
    NANDX1 U39037 (.A1(n50322), .A2(N1048), .ZN(N51909));
    NANDX1 U39038 (.A1(N12579), .A2(n24384), .ZN(N51910));
    INVX1 U39039 (.I(n49793), .ZN(N51911));
    NANDX1 U39040 (.A1(N4454), .A2(n20871), .ZN(N51912));
    NANDX1 U39041 (.A1(n23914), .A2(n32660), .ZN(N51913));
    NOR2X1 U39042 (.A1(n12888), .A2(n33636), .ZN(N51914));
    NANDX1 U39043 (.A1(n23260), .A2(n43396), .ZN(N51915));
    INVX1 U39044 (.I(n32895), .ZN(N51916));
    NOR2X1 U39045 (.A1(n34828), .A2(n28905), .ZN(N51917));
    INVX1 U39046 (.I(n17462), .ZN(N51918));
    NANDX1 U39047 (.A1(n23787), .A2(N1344), .ZN(N51919));
    NANDX1 U39048 (.A1(n41116), .A2(n21693), .ZN(N51920));
    INVX1 U39049 (.I(N12015), .ZN(N51921));
    NANDX1 U39050 (.A1(n23898), .A2(n28384), .ZN(N51922));
    NOR2X1 U39051 (.A1(n26495), .A2(N2865), .ZN(N51923));
    NOR2X1 U39052 (.A1(n47752), .A2(n26778), .ZN(N51924));
    INVX1 U39053 (.I(N12195), .ZN(n51925));
    NOR2X1 U39054 (.A1(N8108), .A2(n17206), .ZN(N51926));
    NOR2X1 U39055 (.A1(n51503), .A2(n30251), .ZN(N51927));
    NOR2X1 U39056 (.A1(n29758), .A2(n35106), .ZN(N51928));
    INVX1 U39057 (.I(N5621), .ZN(N51929));
    NOR2X1 U39058 (.A1(n32546), .A2(n29408), .ZN(N51930));
    NANDX1 U39059 (.A1(n31012), .A2(n18935), .ZN(N51931));
    NANDX1 U39060 (.A1(n30526), .A2(N978), .ZN(N51932));
    INVX1 U39061 (.I(n24452), .ZN(N51933));
    NOR2X1 U39062 (.A1(n22459), .A2(n20974), .ZN(N51934));
    NOR2X1 U39063 (.A1(n45832), .A2(n17137), .ZN(N51935));
    NANDX1 U39064 (.A1(n50275), .A2(n50947), .ZN(n51936));
    NANDX1 U39065 (.A1(N6794), .A2(n38180), .ZN(N51937));
    NANDX1 U39066 (.A1(N6708), .A2(n16842), .ZN(N51938));
    INVX1 U39067 (.I(N6493), .ZN(N51939));
    INVX1 U39068 (.I(N848), .ZN(N51940));
    NOR2X1 U39069 (.A1(n44571), .A2(n33393), .ZN(N51941));
    INVX1 U39070 (.I(n38537), .ZN(N51942));
    NANDX1 U39071 (.A1(n30483), .A2(n24223), .ZN(N51943));
    NANDX1 U39072 (.A1(n31460), .A2(n44179), .ZN(N51944));
    INVX1 U39073 (.I(n30848), .ZN(N51945));
    INVX1 U39074 (.I(n28823), .ZN(N51946));
    INVX1 U39075 (.I(N9292), .ZN(N51947));
    NOR2X1 U39076 (.A1(n32157), .A2(N7979), .ZN(N51948));
    INVX1 U39077 (.I(N10934), .ZN(N51949));
    INVX1 U39078 (.I(N1937), .ZN(N51950));
    NOR2X1 U39079 (.A1(n43096), .A2(n40395), .ZN(N51951));
    NANDX1 U39080 (.A1(n49588), .A2(n32398), .ZN(N51952));
    NOR2X1 U39081 (.A1(n31729), .A2(n46996), .ZN(N51953));
    INVX1 U39082 (.I(n21661), .ZN(N51954));
    NOR2X1 U39083 (.A1(n27404), .A2(N556), .ZN(N51955));
    NOR2X1 U39084 (.A1(N10801), .A2(N2043), .ZN(N51956));
    NOR2X1 U39085 (.A1(n40266), .A2(n32891), .ZN(N51957));
    NOR2X1 U39086 (.A1(n39116), .A2(n36018), .ZN(N51958));
    NANDX1 U39087 (.A1(N3514), .A2(n16587), .ZN(N51959));
    INVX1 U39088 (.I(n40475), .ZN(N51960));
    INVX1 U39089 (.I(n29545), .ZN(N51961));
    NANDX1 U39090 (.A1(n20210), .A2(n42668), .ZN(N51962));
    INVX1 U39091 (.I(N8913), .ZN(N51963));
    INVX1 U39092 (.I(N3671), .ZN(N51964));
    NOR2X1 U39093 (.A1(n42424), .A2(n50666), .ZN(N51965));
    NOR2X1 U39094 (.A1(N12497), .A2(N3049), .ZN(N51966));
    NANDX1 U39095 (.A1(n34668), .A2(n31242), .ZN(N51967));
    INVX1 U39096 (.I(n36710), .ZN(N51968));
    NANDX1 U39097 (.A1(N1603), .A2(n18012), .ZN(N51969));
    NANDX1 U39098 (.A1(n40718), .A2(n24058), .ZN(N51970));
    INVX1 U39099 (.I(n44231), .ZN(N51971));
    NOR2X1 U39100 (.A1(n36220), .A2(N3146), .ZN(n51972));
    INVX1 U39101 (.I(n14177), .ZN(N51973));
    NOR2X1 U39102 (.A1(N6812), .A2(n26872), .ZN(N51974));
    NOR2X1 U39103 (.A1(n37340), .A2(n37567), .ZN(N51975));
    NANDX1 U39104 (.A1(N5831), .A2(n28403), .ZN(N51976));
    NOR2X1 U39105 (.A1(n40496), .A2(N10927), .ZN(N51977));
    NOR2X1 U39106 (.A1(n50977), .A2(n45594), .ZN(N51978));
    NOR2X1 U39107 (.A1(N12314), .A2(n30715), .ZN(N51979));
    NANDX1 U39108 (.A1(n13916), .A2(n18755), .ZN(N51980));
    INVX1 U39109 (.I(N3045), .ZN(N51981));
    NANDX1 U39110 (.A1(n35360), .A2(n17303), .ZN(N51982));
    NANDX1 U39111 (.A1(n19991), .A2(n20448), .ZN(N51983));
    NOR2X1 U39112 (.A1(N4195), .A2(n36032), .ZN(N51984));
    NOR2X1 U39113 (.A1(n31067), .A2(n22889), .ZN(N51985));
    INVX1 U39114 (.I(n17045), .ZN(N51986));
    NOR2X1 U39115 (.A1(n30122), .A2(n15475), .ZN(N51987));
    NOR2X1 U39116 (.A1(n40646), .A2(n26401), .ZN(N51988));
    NANDX1 U39117 (.A1(n40034), .A2(n20406), .ZN(N51989));
    NANDX1 U39118 (.A1(n22375), .A2(n21149), .ZN(N51990));
    NOR2X1 U39119 (.A1(n36290), .A2(n39903), .ZN(N51991));
    INVX1 U39120 (.I(N9362), .ZN(N51992));
    NANDX1 U39121 (.A1(n46482), .A2(n26664), .ZN(N51993));
    INVX1 U39122 (.I(n14884), .ZN(N51994));
    INVX1 U39123 (.I(n34776), .ZN(N51995));
    NOR2X1 U39124 (.A1(N1583), .A2(n21728), .ZN(N51996));
    NANDX1 U39125 (.A1(n46088), .A2(n16048), .ZN(N51997));
    INVX1 U39126 (.I(N7915), .ZN(N51998));
    NOR2X1 U39127 (.A1(n44336), .A2(N2579), .ZN(N51999));
    INVX1 U39128 (.I(n19148), .ZN(N52000));
    INVX1 U39129 (.I(n15315), .ZN(N52001));
    NOR2X1 U39130 (.A1(n22719), .A2(n37689), .ZN(N52002));
    INVX1 U39131 (.I(n19928), .ZN(N52003));
    INVX1 U39132 (.I(n40660), .ZN(N52004));
    NOR2X1 U39133 (.A1(n31751), .A2(N11841), .ZN(N52005));
    NANDX1 U39134 (.A1(n28443), .A2(n36504), .ZN(N52006));
    INVX1 U39135 (.I(n45582), .ZN(N52007));
    NOR2X1 U39136 (.A1(n21577), .A2(n17192), .ZN(N52008));
    NANDX1 U39137 (.A1(N11777), .A2(N11691), .ZN(N52009));
    NANDX1 U39138 (.A1(N10665), .A2(n41222), .ZN(n52010));
    INVX1 U39139 (.I(N3412), .ZN(N52011));
    NOR2X1 U39140 (.A1(n18972), .A2(n44176), .ZN(N52012));
    NOR2X1 U39141 (.A1(n34286), .A2(N2169), .ZN(N52013));
    NANDX1 U39142 (.A1(n20387), .A2(n32898), .ZN(N52014));
    NANDX1 U39143 (.A1(N12804), .A2(n43585), .ZN(N52015));
    NANDX1 U39144 (.A1(n14583), .A2(N3837), .ZN(N52016));
    NANDX1 U39145 (.A1(n43025), .A2(n40340), .ZN(N52017));
    NANDX1 U39146 (.A1(N7046), .A2(n30058), .ZN(N52018));
    NOR2X1 U39147 (.A1(n24237), .A2(N11532), .ZN(N52019));
    NANDX1 U39148 (.A1(n35928), .A2(N9053), .ZN(N52020));
    INVX1 U39149 (.I(n25561), .ZN(N52021));
    INVX1 U39150 (.I(N11781), .ZN(N52022));
    INVX1 U39151 (.I(n41742), .ZN(N52023));
    NOR2X1 U39152 (.A1(n21492), .A2(n24439), .ZN(n52024));
    NANDX1 U39153 (.A1(n26315), .A2(n14853), .ZN(N52025));
    NANDX1 U39154 (.A1(n42709), .A2(n27657), .ZN(N52026));
    NANDX1 U39155 (.A1(n38564), .A2(n42239), .ZN(N52027));
    NANDX1 U39156 (.A1(n30390), .A2(N3703), .ZN(N52028));
    INVX1 U39157 (.I(N3098), .ZN(N52029));
    NANDX1 U39158 (.A1(n37361), .A2(n48970), .ZN(N52030));
    INVX1 U39159 (.I(n48893), .ZN(N52031));
    NOR2X1 U39160 (.A1(n19323), .A2(n27973), .ZN(N52032));
    INVX1 U39161 (.I(n14911), .ZN(N52033));
    NANDX1 U39162 (.A1(n45207), .A2(N2710), .ZN(N52034));
    INVX1 U39163 (.I(n19602), .ZN(N52035));
    INVX1 U39164 (.I(N5391), .ZN(N52036));
    INVX1 U39165 (.I(n20544), .ZN(N52037));
    NOR2X1 U39166 (.A1(N5625), .A2(n33280), .ZN(N52038));
    NANDX1 U39167 (.A1(n28697), .A2(n20255), .ZN(N52039));
    INVX1 U39168 (.I(N4017), .ZN(N52040));
    NOR2X1 U39169 (.A1(n33895), .A2(n41292), .ZN(N52041));
    NANDX1 U39170 (.A1(n44642), .A2(n27064), .ZN(N52042));
    INVX1 U39171 (.I(n49654), .ZN(N52043));
    NOR2X1 U39172 (.A1(N7881), .A2(n39004), .ZN(N52044));
    NANDX1 U39173 (.A1(n41307), .A2(N2327), .ZN(N52045));
    NOR2X1 U39174 (.A1(N4953), .A2(n26652), .ZN(N52046));
    NANDX1 U39175 (.A1(n24554), .A2(n20881), .ZN(N52047));
    NANDX1 U39176 (.A1(n20718), .A2(N11452), .ZN(N52048));
    INVX1 U39177 (.I(n26342), .ZN(N52049));
    INVX1 U39178 (.I(n50938), .ZN(N52050));
    NOR2X1 U39179 (.A1(n35014), .A2(n51158), .ZN(N52051));
    NOR2X1 U39180 (.A1(N4098), .A2(n33465), .ZN(N52052));
    NOR2X1 U39181 (.A1(n19511), .A2(n48134), .ZN(N52053));
    NANDX1 U39182 (.A1(n32306), .A2(n46199), .ZN(N52054));
    INVX1 U39183 (.I(n40187), .ZN(N52055));
    NOR2X1 U39184 (.A1(n45900), .A2(n51521), .ZN(N52056));
    NANDX1 U39185 (.A1(N7479), .A2(n26502), .ZN(N52057));
    INVX1 U39186 (.I(n23213), .ZN(N52058));
    INVX1 U39187 (.I(N1913), .ZN(N52059));
    INVX1 U39188 (.I(n41801), .ZN(N52060));
    NANDX1 U39189 (.A1(n47375), .A2(n38170), .ZN(N52061));
    INVX1 U39190 (.I(n46724), .ZN(N52062));
    NANDX1 U39191 (.A1(N11548), .A2(n46294), .ZN(N52063));
    INVX1 U39192 (.I(n37261), .ZN(N52064));
    INVX1 U39193 (.I(n29542), .ZN(N52065));
    NANDX1 U39194 (.A1(n16359), .A2(n15446), .ZN(N52066));
    INVX1 U39195 (.I(N10970), .ZN(N52067));
    NOR2X1 U39196 (.A1(n26087), .A2(n14612), .ZN(n52068));
    NOR2X1 U39197 (.A1(n47635), .A2(n42196), .ZN(N52069));
    NOR2X1 U39198 (.A1(n22548), .A2(n23227), .ZN(N52070));
    NANDX1 U39199 (.A1(n43631), .A2(n46755), .ZN(N52071));
    NANDX1 U39200 (.A1(n33843), .A2(n30147), .ZN(N52072));
    NOR2X1 U39201 (.A1(n20424), .A2(N6681), .ZN(N52073));
    NOR2X1 U39202 (.A1(n32071), .A2(n39844), .ZN(N52074));
    INVX1 U39203 (.I(n42828), .ZN(N52075));
    INVX1 U39204 (.I(n23839), .ZN(N52076));
    NOR2X1 U39205 (.A1(n30698), .A2(n40197), .ZN(N52077));
    NANDX1 U39206 (.A1(n38214), .A2(n21194), .ZN(N52078));
    INVX1 U39207 (.I(n34328), .ZN(N52079));
    INVX1 U39208 (.I(N5314), .ZN(N52080));
    NOR2X1 U39209 (.A1(n48028), .A2(n16108), .ZN(N52081));
    NANDX1 U39210 (.A1(n19667), .A2(n50114), .ZN(N52082));
    INVX1 U39211 (.I(n36449), .ZN(N52083));
    INVX1 U39212 (.I(n48834), .ZN(n52084));
    INVX1 U39213 (.I(n31109), .ZN(N52085));
    INVX1 U39214 (.I(n43303), .ZN(N52086));
    INVX1 U39215 (.I(n19768), .ZN(N52087));
    INVX1 U39216 (.I(n14482), .ZN(n52088));
    NOR2X1 U39217 (.A1(n27101), .A2(N8348), .ZN(N52089));
    NOR2X1 U39218 (.A1(n27827), .A2(n48544), .ZN(N52090));
    INVX1 U39219 (.I(n14452), .ZN(N52091));
    INVX1 U39220 (.I(N1710), .ZN(N52092));
    NOR2X1 U39221 (.A1(n45598), .A2(n28639), .ZN(n52093));
    NANDX1 U39222 (.A1(n42038), .A2(n44747), .ZN(N52094));
    INVX1 U39223 (.I(n31732), .ZN(N52095));
    INVX1 U39224 (.I(n13919), .ZN(N52096));
    NANDX1 U39225 (.A1(N252), .A2(n32780), .ZN(N52097));
    INVX1 U39226 (.I(n31360), .ZN(N52098));
    NANDX1 U39227 (.A1(n14957), .A2(n41816), .ZN(N52099));
    INVX1 U39228 (.I(n16543), .ZN(N52100));
    NOR2X1 U39229 (.A1(n42895), .A2(n43643), .ZN(N52101));
    INVX1 U39230 (.I(n44710), .ZN(N52102));
    NOR2X1 U39231 (.A1(N1655), .A2(n22805), .ZN(N52103));
    INVX1 U39232 (.I(n41420), .ZN(n52104));
    NANDX1 U39233 (.A1(N1552), .A2(n35430), .ZN(N52105));
    NOR2X1 U39234 (.A1(n29117), .A2(n47495), .ZN(N52106));
    NANDX1 U39235 (.A1(n49659), .A2(n27638), .ZN(N52107));
    NANDX1 U39236 (.A1(n33605), .A2(n14257), .ZN(N52108));
    NANDX1 U39237 (.A1(n14797), .A2(n37499), .ZN(N52109));
    NANDX1 U39238 (.A1(n35273), .A2(N868), .ZN(N52110));
    INVX1 U39239 (.I(n15573), .ZN(N52111));
    NANDX1 U39240 (.A1(n39471), .A2(N6880), .ZN(N52112));
    NOR2X1 U39241 (.A1(n22554), .A2(N1), .ZN(N52113));
    INVX1 U39242 (.I(n24209), .ZN(N52114));
    NOR2X1 U39243 (.A1(n25349), .A2(n35656), .ZN(N52115));
    NANDX1 U39244 (.A1(n26900), .A2(n41113), .ZN(N52116));
    INVX1 U39245 (.I(n26044), .ZN(N52117));
    NANDX1 U39246 (.A1(n48509), .A2(n24114), .ZN(N52118));
    INVX1 U39247 (.I(n18202), .ZN(N52119));
    NANDX1 U39248 (.A1(n18969), .A2(n39735), .ZN(N52120));
    NANDX1 U39249 (.A1(N4879), .A2(N11066), .ZN(N52121));
    INVX1 U39250 (.I(n27362), .ZN(N52122));
    NOR2X1 U39251 (.A1(N11828), .A2(n14799), .ZN(N52123));
    NOR2X1 U39252 (.A1(n18707), .A2(n15907), .ZN(N52124));
    NOR2X1 U39253 (.A1(n40323), .A2(n36895), .ZN(N52125));
    NANDX1 U39254 (.A1(n33155), .A2(n32271), .ZN(N52126));
    NOR2X1 U39255 (.A1(n20529), .A2(N7582), .ZN(N52127));
    INVX1 U39256 (.I(N1111), .ZN(N52128));
    INVX1 U39257 (.I(N1167), .ZN(N52129));
    NANDX1 U39258 (.A1(n27766), .A2(N5879), .ZN(N52130));
    INVX1 U39259 (.I(N3924), .ZN(N52131));
    INVX1 U39260 (.I(n47611), .ZN(N52132));
    NANDX1 U39261 (.A1(n29725), .A2(N7088), .ZN(N52133));
    INVX1 U39262 (.I(n27115), .ZN(N52134));
    NANDX1 U39263 (.A1(N2960), .A2(n41913), .ZN(N52135));
    NANDX1 U39264 (.A1(n21666), .A2(N6231), .ZN(N52136));
    NANDX1 U39265 (.A1(N10400), .A2(n13153), .ZN(N52137));
    INVX1 U39266 (.I(n43554), .ZN(N52138));
    NOR2X1 U39267 (.A1(n34866), .A2(n34111), .ZN(N52139));
    INVX1 U39268 (.I(n50602), .ZN(N52140));
    INVX1 U39269 (.I(n26684), .ZN(N52141));
    INVX1 U39270 (.I(N3280), .ZN(N52142));
    INVX1 U39271 (.I(N6059), .ZN(N52143));
    NANDX1 U39272 (.A1(n28401), .A2(N933), .ZN(N52144));
    NANDX1 U39273 (.A1(n23279), .A2(n30657), .ZN(N52145));
    INVX1 U39274 (.I(n14411), .ZN(N52146));
    INVX1 U39275 (.I(N7237), .ZN(N52147));
    NOR2X1 U39276 (.A1(n18124), .A2(n42275), .ZN(N52148));
    NANDX1 U39277 (.A1(n45970), .A2(n22045), .ZN(N52149));
    INVX1 U39278 (.I(n29151), .ZN(N52150));
    INVX1 U39279 (.I(n33043), .ZN(N52151));
    NOR2X1 U39280 (.A1(N5620), .A2(n15565), .ZN(N52152));
    INVX1 U39281 (.I(N4634), .ZN(N52153));
    NOR2X1 U39282 (.A1(N12756), .A2(n26430), .ZN(N52154));
    INVX1 U39283 (.I(n37233), .ZN(N52155));
    INVX1 U39284 (.I(n26892), .ZN(N52156));
    NOR2X1 U39285 (.A1(n33420), .A2(n34069), .ZN(N52157));
    NANDX1 U39286 (.A1(n34104), .A2(n18361), .ZN(N52158));
    INVX1 U39287 (.I(n31931), .ZN(N52159));
    INVX1 U39288 (.I(N9159), .ZN(N52160));
    NANDX1 U39289 (.A1(n37899), .A2(n18221), .ZN(N52161));
    NOR2X1 U39290 (.A1(n29971), .A2(N7710), .ZN(N52162));
    NANDX1 U39291 (.A1(N725), .A2(n40752), .ZN(N52163));
    NANDX1 U39292 (.A1(N6345), .A2(n26345), .ZN(N52164));
    NOR2X1 U39293 (.A1(n32594), .A2(n17186), .ZN(N52165));
    NANDX1 U39294 (.A1(N7435), .A2(n32922), .ZN(N52166));
    NOR2X1 U39295 (.A1(N9950), .A2(N8225), .ZN(N52167));
    NANDX1 U39296 (.A1(n13397), .A2(n42293), .ZN(N52168));
    INVX1 U39297 (.I(n17528), .ZN(N52169));
    NOR2X1 U39298 (.A1(n25927), .A2(n49458), .ZN(N52170));
    NANDX1 U39299 (.A1(N5113), .A2(n17951), .ZN(N52171));
    NANDX1 U39300 (.A1(n23333), .A2(n32414), .ZN(N52172));
    NOR2X1 U39301 (.A1(n31042), .A2(n24438), .ZN(N52173));
    NANDX1 U39302 (.A1(n41821), .A2(n31091), .ZN(N52174));
    INVX1 U39303 (.I(n16577), .ZN(N52175));
    INVX1 U39304 (.I(n43920), .ZN(N52176));
    NOR2X1 U39305 (.A1(N7681), .A2(n51354), .ZN(N52177));
    NANDX1 U39306 (.A1(n50394), .A2(n31331), .ZN(N52178));
    NOR2X1 U39307 (.A1(n25592), .A2(n44727), .ZN(N52179));
    NANDX1 U39308 (.A1(n29757), .A2(N10667), .ZN(N52180));
    NOR2X1 U39309 (.A1(N4095), .A2(N8536), .ZN(n52181));
    INVX1 U39310 (.I(N9207), .ZN(N52182));
    NOR2X1 U39311 (.A1(n15324), .A2(N2567), .ZN(N52183));
    NANDX1 U39312 (.A1(n49554), .A2(N3636), .ZN(N52184));
    NANDX1 U39313 (.A1(n32921), .A2(n45456), .ZN(N52185));
    INVX1 U39314 (.I(n44247), .ZN(N52186));
    NANDX1 U39315 (.A1(n26711), .A2(n36579), .ZN(N52187));
    NANDX1 U39316 (.A1(N4419), .A2(N6372), .ZN(N52188));
    INVX1 U39317 (.I(N3224), .ZN(N52189));
    NANDX1 U39318 (.A1(n22675), .A2(n50431), .ZN(N52190));
    INVX1 U39319 (.I(n28342), .ZN(N52191));
    NOR2X1 U39320 (.A1(N11535), .A2(n13101), .ZN(N52192));
    NOR2X1 U39321 (.A1(n20071), .A2(n45781), .ZN(N52193));
    NANDX1 U39322 (.A1(n16585), .A2(n31132), .ZN(N52194));
    INVX1 U39323 (.I(n45512), .ZN(N52195));
    INVX1 U39324 (.I(n39744), .ZN(N52196));
    NOR2X1 U39325 (.A1(N10430), .A2(n33612), .ZN(N52197));
    INVX1 U39326 (.I(n24704), .ZN(N52198));
    INVX1 U39327 (.I(n38566), .ZN(N52199));
    INVX1 U39328 (.I(N6701), .ZN(N52200));
    NOR2X1 U39329 (.A1(n37682), .A2(N6057), .ZN(N52201));
    NOR2X1 U39330 (.A1(n23796), .A2(n50348), .ZN(N52202));
    NOR2X1 U39331 (.A1(n24664), .A2(n48717), .ZN(N52203));
    INVX1 U39332 (.I(n36199), .ZN(N52204));
    NOR2X1 U39333 (.A1(n16425), .A2(n26297), .ZN(N52205));
    NOR2X1 U39334 (.A1(n49968), .A2(n12909), .ZN(n52206));
    NOR2X1 U39335 (.A1(N4516), .A2(n28448), .ZN(N52207));
    INVX1 U39336 (.I(n44260), .ZN(N52208));
    NANDX1 U39337 (.A1(n36750), .A2(n26283), .ZN(N52209));
    NOR2X1 U39338 (.A1(N9866), .A2(n40366), .ZN(N52210));
    NOR2X1 U39339 (.A1(n19559), .A2(n17094), .ZN(N52211));
    NANDX1 U39340 (.A1(n27268), .A2(n44767), .ZN(N52212));
    NANDX1 U39341 (.A1(n51063), .A2(n13554), .ZN(N52213));
    NANDX1 U39342 (.A1(n45755), .A2(N10682), .ZN(N52214));
    NOR2X1 U39343 (.A1(N393), .A2(n42526), .ZN(N52215));
    NOR2X1 U39344 (.A1(n48305), .A2(n38590), .ZN(N52216));
    NOR2X1 U39345 (.A1(N9625), .A2(n14197), .ZN(N52217));
    INVX1 U39346 (.I(n38072), .ZN(N52218));
    NANDX1 U39347 (.A1(n46313), .A2(n23890), .ZN(N52219));
    INVX1 U39348 (.I(n21007), .ZN(N52220));
    NOR2X1 U39349 (.A1(n13928), .A2(n31400), .ZN(N52221));
    NOR2X1 U39350 (.A1(N3515), .A2(n18521), .ZN(N52222));
    NOR2X1 U39351 (.A1(N810), .A2(N11699), .ZN(N52223));
    INVX1 U39352 (.I(n21901), .ZN(N52224));
    NANDX1 U39353 (.A1(n28581), .A2(n16067), .ZN(N52225));
    NOR2X1 U39354 (.A1(n19671), .A2(n16459), .ZN(N52226));
    INVX1 U39355 (.I(n27186), .ZN(N52227));
    NANDX1 U39356 (.A1(N5515), .A2(N3107), .ZN(N52228));
    NOR2X1 U39357 (.A1(n41328), .A2(N5160), .ZN(N52229));
    NANDX1 U39358 (.A1(n30257), .A2(n51472), .ZN(N52230));
    NANDX1 U39359 (.A1(N4347), .A2(n42506), .ZN(N52231));
    NOR2X1 U39360 (.A1(n39891), .A2(n43933), .ZN(N52232));
    NANDX1 U39361 (.A1(n43405), .A2(N10866), .ZN(N52233));
    NANDX1 U39362 (.A1(n44214), .A2(n44180), .ZN(N52234));
    NOR2X1 U39363 (.A1(n36142), .A2(n39460), .ZN(N52235));
    NOR2X1 U39364 (.A1(N620), .A2(n15448), .ZN(N52236));
    NOR2X1 U39365 (.A1(n38694), .A2(n33962), .ZN(N52237));
    NANDX1 U39366 (.A1(n21896), .A2(N9504), .ZN(n52238));
    INVX1 U39367 (.I(n14722), .ZN(N52239));
    NOR2X1 U39368 (.A1(N1721), .A2(n15647), .ZN(N52240));
    INVX1 U39369 (.I(n23220), .ZN(N52241));
    NANDX1 U39370 (.A1(N3874), .A2(n14138), .ZN(N52242));
    INVX1 U39371 (.I(n43764), .ZN(N52243));
    NANDX1 U39372 (.A1(n22992), .A2(N5608), .ZN(N52244));
    NANDX1 U39373 (.A1(N9704), .A2(n19849), .ZN(N52245));
    INVX1 U39374 (.I(n39254), .ZN(N52246));
    NANDX1 U39375 (.A1(n41042), .A2(n15824), .ZN(N52247));
    NOR2X1 U39376 (.A1(N4901), .A2(n42037), .ZN(N52248));
    INVX1 U39377 (.I(N8890), .ZN(N52249));
    NOR2X1 U39378 (.A1(n35639), .A2(n40010), .ZN(N52250));
    NANDX1 U39379 (.A1(n20389), .A2(N9280), .ZN(N52251));
    INVX1 U39380 (.I(N6063), .ZN(N52252));
    NANDX1 U39381 (.A1(N5403), .A2(n16552), .ZN(N52253));
    NOR2X1 U39382 (.A1(n41156), .A2(n21830), .ZN(N52254));
    NANDX1 U39383 (.A1(n17666), .A2(n44822), .ZN(N52255));
    NOR2X1 U39384 (.A1(N5040), .A2(n24553), .ZN(N52256));
    NOR2X1 U39385 (.A1(N6622), .A2(n33834), .ZN(N52257));
    INVX1 U39386 (.I(n47663), .ZN(N52258));
    INVX1 U39387 (.I(N1406), .ZN(N52259));
    NANDX1 U39388 (.A1(N10134), .A2(n15149), .ZN(N52260));
    NANDX1 U39389 (.A1(n45624), .A2(n20815), .ZN(N52261));
    NOR2X1 U39390 (.A1(N4471), .A2(n41203), .ZN(N52262));
    INVX1 U39391 (.I(n38242), .ZN(N52263));
    INVX1 U39392 (.I(N8016), .ZN(N52264));
    INVX1 U39393 (.I(n33845), .ZN(N52265));
    NANDX1 U39394 (.A1(n33212), .A2(N4087), .ZN(N52266));
    INVX1 U39395 (.I(n50877), .ZN(N52267));
    NOR2X1 U39396 (.A1(n40914), .A2(n25945), .ZN(N52268));
    INVX1 U39397 (.I(N11279), .ZN(N52269));
    INVX1 U39398 (.I(n17377), .ZN(N52270));
    INVX1 U39399 (.I(n50257), .ZN(N52271));
    INVX1 U39400 (.I(n30684), .ZN(N52272));
    NANDX1 U39401 (.A1(n47194), .A2(n15860), .ZN(N52273));
    INVX1 U39402 (.I(n41230), .ZN(N52274));
    NANDX1 U39403 (.A1(n42670), .A2(n45700), .ZN(N52275));
    INVX1 U39404 (.I(n41879), .ZN(N52276));
    NOR2X1 U39405 (.A1(n43582), .A2(n19922), .ZN(N52277));
    INVX1 U39406 (.I(n47454), .ZN(N52278));
    NOR2X1 U39407 (.A1(n19293), .A2(n51540), .ZN(N52279));
    NOR2X1 U39408 (.A1(n40198), .A2(n40503), .ZN(N52280));
    NOR2X1 U39409 (.A1(n14554), .A2(N2430), .ZN(N52281));
    INVX1 U39410 (.I(n17147), .ZN(N52282));
    NOR2X1 U39411 (.A1(n49361), .A2(n15815), .ZN(N52283));
    NANDX1 U39412 (.A1(n28456), .A2(N7102), .ZN(N52284));
    NOR2X1 U39413 (.A1(n44315), .A2(n29870), .ZN(N52285));
    NOR2X1 U39414 (.A1(n29401), .A2(n42567), .ZN(N52286));
    NANDX1 U39415 (.A1(n47333), .A2(n32857), .ZN(N52287));
    NANDX1 U39416 (.A1(n39326), .A2(N1190), .ZN(N52288));
    NANDX1 U39417 (.A1(N5219), .A2(n33449), .ZN(N52289));
    NANDX1 U39418 (.A1(N5171), .A2(N1340), .ZN(N52290));
    NANDX1 U39419 (.A1(n15701), .A2(N10144), .ZN(N52291));
    NOR2X1 U39420 (.A1(n39747), .A2(N254), .ZN(N52292));
    NANDX1 U39421 (.A1(N7964), .A2(n49615), .ZN(N52293));
    INVX1 U39422 (.I(n34858), .ZN(N52294));
    INVX1 U39423 (.I(n40520), .ZN(N52295));
    NANDX1 U39424 (.A1(n40825), .A2(n18801), .ZN(N52296));
    INVX1 U39425 (.I(n18637), .ZN(N52297));
    NOR2X1 U39426 (.A1(n37422), .A2(n35997), .ZN(N52298));
    NOR2X1 U39427 (.A1(n37699), .A2(n45350), .ZN(N52299));
    NANDX1 U39428 (.A1(n24057), .A2(n50568), .ZN(N52300));
    INVX1 U39429 (.I(n29708), .ZN(N52301));
    NANDX1 U39430 (.A1(n40283), .A2(n45583), .ZN(N52302));
    INVX1 U39431 (.I(n20454), .ZN(N52303));
    INVX1 U39432 (.I(n29625), .ZN(N52304));
    INVX1 U39433 (.I(n42027), .ZN(N52305));
    NANDX1 U39434 (.A1(n18733), .A2(n23856), .ZN(N52306));
    INVX1 U39435 (.I(n15243), .ZN(N52307));
    NANDX1 U39436 (.A1(n39887), .A2(N4479), .ZN(N52308));
    NANDX1 U39437 (.A1(n49440), .A2(n44731), .ZN(N52309));
    INVX1 U39438 (.I(n35274), .ZN(N52310));
    NOR2X1 U39439 (.A1(n37315), .A2(n43000), .ZN(N52311));
    INVX1 U39440 (.I(n21194), .ZN(N52312));
    INVX1 U39441 (.I(n21879), .ZN(N52313));
    NOR2X1 U39442 (.A1(n15204), .A2(n47645), .ZN(N52314));
    INVX1 U39443 (.I(n30814), .ZN(N52315));
    NOR2X1 U39444 (.A1(n39312), .A2(N3649), .ZN(N52316));
    NANDX1 U39445 (.A1(n30047), .A2(n45675), .ZN(N52317));
    INVX1 U39446 (.I(n18807), .ZN(N52318));
    INVX1 U39447 (.I(n27319), .ZN(N52319));
    NANDX1 U39448 (.A1(n22373), .A2(n15617), .ZN(N52320));
    NANDX1 U39449 (.A1(n45604), .A2(n13469), .ZN(N52321));
    NOR2X1 U39450 (.A1(n48640), .A2(n18770), .ZN(N52322));
    NANDX1 U39451 (.A1(n34367), .A2(N10181), .ZN(N52323));
    NOR2X1 U39452 (.A1(n25588), .A2(n47265), .ZN(N52324));
    INVX1 U39453 (.I(N4165), .ZN(N52325));
    NOR2X1 U39454 (.A1(N3369), .A2(n23023), .ZN(n52326));
    INVX1 U39455 (.I(N10919), .ZN(N52327));
    NANDX1 U39456 (.A1(n15370), .A2(n18121), .ZN(n52328));
    INVX1 U39457 (.I(n31073), .ZN(N52329));
    INVX1 U39458 (.I(n51243), .ZN(N52330));
    NANDX1 U39459 (.A1(N8669), .A2(N3732), .ZN(N52331));
    NOR2X1 U39460 (.A1(n24285), .A2(N12286), .ZN(N52332));
    NOR2X1 U39461 (.A1(N7781), .A2(n35599), .ZN(N52333));
    INVX1 U39462 (.I(n26550), .ZN(N52334));
    NOR2X1 U39463 (.A1(n36876), .A2(N6759), .ZN(N52335));
    NOR2X1 U39464 (.A1(N10875), .A2(N2435), .ZN(N52336));
    INVX1 U39465 (.I(n15039), .ZN(N52337));
    NANDX1 U39466 (.A1(N10959), .A2(N8090), .ZN(N52338));
    NOR2X1 U39467 (.A1(n21877), .A2(N10480), .ZN(N52339));
    NOR2X1 U39468 (.A1(n39997), .A2(n42916), .ZN(N52340));
    NANDX1 U39469 (.A1(n42962), .A2(n42570), .ZN(N52341));
    NOR2X1 U39470 (.A1(N42), .A2(n46301), .ZN(N52342));
    INVX1 U39471 (.I(n45943), .ZN(N52343));
    INVX1 U39472 (.I(n47475), .ZN(N52344));
    NANDX1 U39473 (.A1(n34241), .A2(n49984), .ZN(N52345));
    NOR2X1 U39474 (.A1(N10757), .A2(n35271), .ZN(N52346));
    NANDX1 U39475 (.A1(n32651), .A2(n16174), .ZN(N52347));
    INVX1 U39476 (.I(n40241), .ZN(N52348));
    NOR2X1 U39477 (.A1(n34479), .A2(n51199), .ZN(N52349));
    NANDX1 U39478 (.A1(n51158), .A2(n43103), .ZN(N52350));
    NANDX1 U39479 (.A1(N1647), .A2(N1539), .ZN(N52351));
    NANDX1 U39480 (.A1(N4823), .A2(n44501), .ZN(N52352));
    NOR2X1 U39481 (.A1(N5426), .A2(n44542), .ZN(N52353));
    NANDX1 U39482 (.A1(n17471), .A2(N8924), .ZN(N52354));
    NOR2X1 U39483 (.A1(n34973), .A2(n32675), .ZN(N52355));
    INVX1 U39484 (.I(N3397), .ZN(N52356));
    INVX1 U39485 (.I(n32112), .ZN(N52357));
    NOR2X1 U39486 (.A1(N6885), .A2(n34790), .ZN(N52358));
    INVX1 U39487 (.I(N6433), .ZN(N52359));
    INVX1 U39488 (.I(N4492), .ZN(N52360));
    INVX1 U39489 (.I(n23053), .ZN(N52361));
    NOR2X1 U39490 (.A1(N10509), .A2(n36184), .ZN(N52362));
    NANDX1 U39491 (.A1(n33771), .A2(n37722), .ZN(N52363));
    INVX1 U39492 (.I(n38594), .ZN(N52364));
    INVX1 U39493 (.I(n30166), .ZN(N52365));
    INVX1 U39494 (.I(n45204), .ZN(N52366));
    NOR2X1 U39495 (.A1(N1545), .A2(N2539), .ZN(N52367));
    NANDX1 U39496 (.A1(n36517), .A2(n35213), .ZN(N52368));
    INVX1 U39497 (.I(N9941), .ZN(N52369));
    NOR2X1 U39498 (.A1(n50863), .A2(n48608), .ZN(N52370));
    NANDX1 U39499 (.A1(n34064), .A2(n21887), .ZN(N52371));
    INVX1 U39500 (.I(N5918), .ZN(N52372));
    NOR2X1 U39501 (.A1(n30911), .A2(n50587), .ZN(N52373));
    NOR2X1 U39502 (.A1(N11447), .A2(n35182), .ZN(N52374));
    NANDX1 U39503 (.A1(n45218), .A2(n42931), .ZN(N52375));
    NANDX1 U39504 (.A1(N2251), .A2(n43593), .ZN(N52376));
    NOR2X1 U39505 (.A1(n16297), .A2(n37208), .ZN(N52377));
    NOR2X1 U39506 (.A1(n39457), .A2(n39746), .ZN(N52378));
    NANDX1 U39507 (.A1(n46001), .A2(n44987), .ZN(N52379));
    NANDX1 U39508 (.A1(N4354), .A2(n30025), .ZN(N52380));
    NOR2X1 U39509 (.A1(n22989), .A2(n43564), .ZN(N52381));
    NANDX1 U39510 (.A1(n14903), .A2(N11947), .ZN(N52382));
    INVX1 U39511 (.I(N11309), .ZN(N52383));
    NOR2X1 U39512 (.A1(n33602), .A2(n13178), .ZN(N52384));
    INVX1 U39513 (.I(n38811), .ZN(N52385));
    NOR2X1 U39514 (.A1(n17960), .A2(n30154), .ZN(N52386));
    NANDX1 U39515 (.A1(n41826), .A2(n22158), .ZN(N52387));
    NANDX1 U39516 (.A1(n28150), .A2(N7777), .ZN(N52388));
    INVX1 U39517 (.I(n16018), .ZN(N52389));
    NOR2X1 U39518 (.A1(n15321), .A2(N10431), .ZN(N52390));
    INVX1 U39519 (.I(n19025), .ZN(N52391));
    NOR2X1 U39520 (.A1(N11001), .A2(n22004), .ZN(N52392));
    NOR2X1 U39521 (.A1(N2976), .A2(N7458), .ZN(N52393));
    INVX1 U39522 (.I(n36538), .ZN(N52394));
    INVX1 U39523 (.I(N4038), .ZN(N52395));
    NOR2X1 U39524 (.A1(n24075), .A2(n17215), .ZN(N52396));
    INVX1 U39525 (.I(N11297), .ZN(N52397));
    INVX1 U39526 (.I(N10152), .ZN(N52398));
    NANDX1 U39527 (.A1(N6631), .A2(n22005), .ZN(N52399));
    NANDX1 U39528 (.A1(n27824), .A2(n50155), .ZN(N52400));
    NOR2X1 U39529 (.A1(n28219), .A2(n14584), .ZN(N52401));
    NOR2X1 U39530 (.A1(n13567), .A2(n46630), .ZN(N52402));
    INVX1 U39531 (.I(n32591), .ZN(N52403));
    INVX1 U39532 (.I(n42580), .ZN(N52404));
    NOR2X1 U39533 (.A1(n39240), .A2(n15583), .ZN(N52405));
    NOR2X1 U39534 (.A1(N10354), .A2(N532), .ZN(N52406));
    INVX1 U39535 (.I(n14391), .ZN(N52407));
    INVX1 U39536 (.I(n16654), .ZN(N52408));
    NANDX1 U39537 (.A1(N12173), .A2(n27950), .ZN(N52409));
    NANDX1 U39538 (.A1(n43940), .A2(n39428), .ZN(N52410));
    NOR2X1 U39539 (.A1(n14356), .A2(n21474), .ZN(N52411));
    NOR2X1 U39540 (.A1(n34538), .A2(N2941), .ZN(N52412));
    NOR2X1 U39541 (.A1(n19150), .A2(N1957), .ZN(N52413));
    NOR2X1 U39542 (.A1(n14191), .A2(N11920), .ZN(N52414));
    NANDX1 U39543 (.A1(n45632), .A2(n24528), .ZN(N52415));
    NOR2X1 U39544 (.A1(n33283), .A2(n40110), .ZN(N52416));
    NOR2X1 U39545 (.A1(n13664), .A2(N10670), .ZN(N52417));
    INVX1 U39546 (.I(n28055), .ZN(N52418));
    NANDX1 U39547 (.A1(N10861), .A2(n29688), .ZN(N52419));
    INVX1 U39548 (.I(n38811), .ZN(N52420));
    NANDX1 U39549 (.A1(n26817), .A2(n48266), .ZN(N52421));
    NOR2X1 U39550 (.A1(N11201), .A2(n39767), .ZN(N52422));
    NANDX1 U39551 (.A1(n45738), .A2(n42707), .ZN(N52423));
    NANDX1 U39552 (.A1(n13299), .A2(n44663), .ZN(N52424));
    INVX1 U39553 (.I(n49106), .ZN(N52425));
    INVX1 U39554 (.I(n47535), .ZN(N52426));
    NOR2X1 U39555 (.A1(n51138), .A2(n47057), .ZN(N52427));
    INVX1 U39556 (.I(n39659), .ZN(N52428));
    NANDX1 U39557 (.A1(n30151), .A2(n20356), .ZN(N52429));
    NOR2X1 U39558 (.A1(N6617), .A2(n21034), .ZN(n52430));
    INVX1 U39559 (.I(N6332), .ZN(N52431));
    INVX1 U39560 (.I(n32620), .ZN(N52432));
    INVX1 U39561 (.I(n30728), .ZN(N52433));
    NANDX1 U39562 (.A1(n48381), .A2(n41928), .ZN(N52434));
    INVX1 U39563 (.I(n13637), .ZN(N52435));
    NOR2X1 U39564 (.A1(N238), .A2(n40785), .ZN(N52436));
    NOR2X1 U39565 (.A1(n14928), .A2(N10243), .ZN(N52437));
    NANDX1 U39566 (.A1(n41538), .A2(N6190), .ZN(N52438));
    NANDX1 U39567 (.A1(N11115), .A2(n23274), .ZN(N52439));
    NOR2X1 U39568 (.A1(n20802), .A2(n41987), .ZN(N52440));
    NOR2X1 U39569 (.A1(n41157), .A2(N3320), .ZN(N52441));
    INVX1 U39570 (.I(N10602), .ZN(N52442));
    NANDX1 U39571 (.A1(n29736), .A2(n14513), .ZN(N52443));
    NANDX1 U39572 (.A1(n13387), .A2(n45240), .ZN(N52444));
    INVX1 U39573 (.I(n31795), .ZN(N52445));
    NANDX1 U39574 (.A1(n16574), .A2(n45432), .ZN(N52446));
    INVX1 U39575 (.I(n16811), .ZN(N52447));
    NANDX1 U39576 (.A1(n31114), .A2(n31739), .ZN(N52448));
    NOR2X1 U39577 (.A1(n39678), .A2(n43304), .ZN(N52449));
    INVX1 U39578 (.I(n39802), .ZN(N52450));
    NANDX1 U39579 (.A1(n44361), .A2(N4825), .ZN(N52451));
    NANDX1 U39580 (.A1(n34760), .A2(n51585), .ZN(N52452));
    INVX1 U39581 (.I(N8107), .ZN(N52453));
    INVX1 U39582 (.I(n15446), .ZN(n52454));
    NANDX1 U39583 (.A1(N1549), .A2(n29958), .ZN(N52455));
    INVX1 U39584 (.I(n36551), .ZN(N52456));
    NOR2X1 U39585 (.A1(n42437), .A2(n16758), .ZN(N52457));
    NANDX1 U39586 (.A1(N7422), .A2(n32217), .ZN(N52458));
    NOR2X1 U39587 (.A1(n24233), .A2(n15256), .ZN(N52459));
    INVX1 U39588 (.I(n25999), .ZN(N52460));
    INVX1 U39589 (.I(N184), .ZN(N52461));
    NANDX1 U39590 (.A1(n21269), .A2(n39986), .ZN(N52462));
    INVX1 U39591 (.I(n14042), .ZN(N52463));
    NANDX1 U39592 (.A1(n35819), .A2(n18829), .ZN(N52464));
    INVX1 U39593 (.I(n40663), .ZN(N52465));
    INVX1 U39594 (.I(n16619), .ZN(N52466));
    NOR2X1 U39595 (.A1(n32169), .A2(n39784), .ZN(N52467));
    NANDX1 U39596 (.A1(n45534), .A2(n24746), .ZN(N52468));
    NANDX1 U39597 (.A1(N6410), .A2(n41503), .ZN(N52469));
    NOR2X1 U39598 (.A1(n13831), .A2(n43747), .ZN(N52470));
    NANDX1 U39599 (.A1(N8091), .A2(n29031), .ZN(N52471));
    NOR2X1 U39600 (.A1(n34089), .A2(n29212), .ZN(N52472));
    INVX1 U39601 (.I(n21831), .ZN(N52473));
    NOR2X1 U39602 (.A1(n30626), .A2(N12402), .ZN(N52474));
    INVX1 U39603 (.I(n45463), .ZN(N52475));
    NOR2X1 U39604 (.A1(N1790), .A2(N8708), .ZN(N52476));
    NOR2X1 U39605 (.A1(n28724), .A2(n46943), .ZN(N52477));
    NANDX1 U39606 (.A1(N9304), .A2(n35138), .ZN(N52478));
    INVX1 U39607 (.I(n24865), .ZN(N52479));
    INVX1 U39608 (.I(n49362), .ZN(N52480));
    NANDX1 U39609 (.A1(n41442), .A2(n16772), .ZN(N52481));
    NOR2X1 U39610 (.A1(n33600), .A2(n16750), .ZN(N52482));
    INVX1 U39611 (.I(N11042), .ZN(N52483));
    INVX1 U39612 (.I(n27339), .ZN(N52484));
    NOR2X1 U39613 (.A1(n19463), .A2(n19197), .ZN(N52485));
    NANDX1 U39614 (.A1(n50088), .A2(n31599), .ZN(N52486));
    NOR2X1 U39615 (.A1(n13990), .A2(n19875), .ZN(N52487));
    INVX1 U39616 (.I(n22697), .ZN(N52488));
    NOR2X1 U39617 (.A1(n22647), .A2(n39667), .ZN(N52489));
    NANDX1 U39618 (.A1(N1978), .A2(n23216), .ZN(N52490));
    NOR2X1 U39619 (.A1(n48458), .A2(N1539), .ZN(N52491));
    NANDX1 U39620 (.A1(n28143), .A2(n42980), .ZN(N52492));
    NOR2X1 U39621 (.A1(n13302), .A2(n46607), .ZN(N52493));
    NOR2X1 U39622 (.A1(N6552), .A2(N6061), .ZN(N52494));
    INVX1 U39623 (.I(N3919), .ZN(N52495));
    INVX1 U39624 (.I(N6716), .ZN(N52496));
    NOR2X1 U39625 (.A1(N3899), .A2(n26831), .ZN(N52497));
    NOR2X1 U39626 (.A1(n47621), .A2(n40820), .ZN(N52498));
    NANDX1 U39627 (.A1(n19928), .A2(n33545), .ZN(N52499));
    INVX1 U39628 (.I(N12602), .ZN(N52500));
    NANDX1 U39629 (.A1(N12576), .A2(n14579), .ZN(N52501));
    NANDX1 U39630 (.A1(n42890), .A2(N11448), .ZN(N52502));
    NANDX1 U39631 (.A1(n19389), .A2(N9618), .ZN(N52503));
    INVX1 U39632 (.I(n34275), .ZN(N52504));
    NANDX1 U39633 (.A1(n46046), .A2(n14323), .ZN(N52505));
    NOR2X1 U39634 (.A1(n22134), .A2(N1576), .ZN(N52506));
    NOR2X1 U39635 (.A1(N8503), .A2(n29908), .ZN(N52507));
    NOR2X1 U39636 (.A1(n34017), .A2(N5150), .ZN(N52508));
    INVX1 U39637 (.I(n30049), .ZN(N52509));
    NANDX1 U39638 (.A1(n35942), .A2(n20004), .ZN(N52510));
    NOR2X1 U39639 (.A1(n47809), .A2(n32605), .ZN(N52511));
    NANDX1 U39640 (.A1(N8796), .A2(n47183), .ZN(N52512));
    INVX1 U39641 (.I(n21714), .ZN(N52513));
    NANDX1 U39642 (.A1(n34134), .A2(n41102), .ZN(N52514));
    INVX1 U39643 (.I(N3601), .ZN(N52515));
    NANDX1 U39644 (.A1(n31222), .A2(n19675), .ZN(N52516));
    NOR2X1 U39645 (.A1(n30720), .A2(n41808), .ZN(N52517));
    NOR2X1 U39646 (.A1(N4164), .A2(n50311), .ZN(n52518));
    NOR2X1 U39647 (.A1(n22338), .A2(n32739), .ZN(N52519));
    NOR2X1 U39648 (.A1(n13665), .A2(n32816), .ZN(N52520));
    INVX1 U39649 (.I(n19635), .ZN(N52521));
    INVX1 U39650 (.I(n50365), .ZN(N52522));
    INVX1 U39651 (.I(N3864), .ZN(N52523));
    NOR2X1 U39652 (.A1(n16294), .A2(n51046), .ZN(N52524));
    INVX1 U39653 (.I(n38007), .ZN(N52525));
    INVX1 U39654 (.I(n40243), .ZN(N52526));
    NOR2X1 U39655 (.A1(n36418), .A2(n43844), .ZN(N52527));
    NANDX1 U39656 (.A1(n37667), .A2(N11930), .ZN(N52528));
    INVX1 U39657 (.I(n38414), .ZN(N52529));
    NANDX1 U39658 (.A1(N9216), .A2(N12605), .ZN(N52530));
    NANDX1 U39659 (.A1(n18865), .A2(n34943), .ZN(N52531));
    NOR2X1 U39660 (.A1(N3691), .A2(n18635), .ZN(N52532));
    NANDX1 U39661 (.A1(n34486), .A2(N8297), .ZN(N52533));
    NANDX1 U39662 (.A1(N3290), .A2(n45767), .ZN(N52534));
    INVX1 U39663 (.I(n13285), .ZN(N52535));
    INVX1 U39664 (.I(N2676), .ZN(N52536));
    INVX1 U39665 (.I(n40123), .ZN(N52537));
    INVX1 U39666 (.I(n38021), .ZN(N52538));
    NOR2X1 U39667 (.A1(N7264), .A2(n30276), .ZN(N52539));
    INVX1 U39668 (.I(n14959), .ZN(N52540));
    NANDX1 U39669 (.A1(n28537), .A2(N1784), .ZN(N52541));
    NOR2X1 U39670 (.A1(N7781), .A2(n14389), .ZN(N52542));
    NOR2X1 U39671 (.A1(n48261), .A2(n19359), .ZN(N52543));
    NANDX1 U39672 (.A1(N363), .A2(n37993), .ZN(N52544));
    INVX1 U39673 (.I(N4876), .ZN(n52545));
    NOR2X1 U39674 (.A1(n51243), .A2(N8165), .ZN(N52546));
    NANDX1 U39675 (.A1(n32845), .A2(n21449), .ZN(N52547));
    NANDX1 U39676 (.A1(N5548), .A2(n19227), .ZN(N52548));
    NOR2X1 U39677 (.A1(n27982), .A2(n27275), .ZN(N52549));
    NANDX1 U39678 (.A1(N5273), .A2(n27578), .ZN(N52550));
    INVX1 U39679 (.I(n20231), .ZN(N52551));
    NOR2X1 U39680 (.A1(n44800), .A2(n22015), .ZN(N52552));
    NOR2X1 U39681 (.A1(n22608), .A2(N6431), .ZN(N52553));
    NANDX1 U39682 (.A1(n19280), .A2(n25789), .ZN(N52554));
    INVX1 U39683 (.I(n41258), .ZN(N52555));
    INVX1 U39684 (.I(n46849), .ZN(N52556));
    NANDX1 U39685 (.A1(n28510), .A2(n46504), .ZN(N52557));
    NOR2X1 U39686 (.A1(n39006), .A2(n49376), .ZN(N52558));
    NANDX1 U39687 (.A1(n30001), .A2(n24951), .ZN(N52559));
    NANDX1 U39688 (.A1(n31147), .A2(N1344), .ZN(N52560));
    INVX1 U39689 (.I(n48348), .ZN(N52561));
    NANDX1 U39690 (.A1(n38291), .A2(n34639), .ZN(N52562));
    NANDX1 U39691 (.A1(n48128), .A2(n49466), .ZN(N52563));
    NANDX1 U39692 (.A1(n42373), .A2(n20486), .ZN(N52564));
    INVX1 U39693 (.I(n35158), .ZN(N52565));
    INVX1 U39694 (.I(n42751), .ZN(N52566));
    INVX1 U39695 (.I(n51051), .ZN(N52567));
    INVX1 U39696 (.I(n25379), .ZN(N52568));
    INVX1 U39697 (.I(N1893), .ZN(N52569));
    NOR2X1 U39698 (.A1(n48304), .A2(n40898), .ZN(N52570));
    INVX1 U39699 (.I(n42489), .ZN(N52571));
    NOR2X1 U39700 (.A1(n13059), .A2(N4312), .ZN(N52572));
    INVX1 U39701 (.I(n36018), .ZN(N52573));
    INVX1 U39702 (.I(n38860), .ZN(N52574));
    NANDX1 U39703 (.A1(n23343), .A2(n21910), .ZN(N52575));
    NOR2X1 U39704 (.A1(n41498), .A2(n19787), .ZN(N52576));
    INVX1 U39705 (.I(N2310), .ZN(n52577));
    INVX1 U39706 (.I(n28673), .ZN(N52578));
    NOR2X1 U39707 (.A1(n20093), .A2(n19835), .ZN(N52579));
    INVX1 U39708 (.I(n19555), .ZN(N52580));
    INVX1 U39709 (.I(N11403), .ZN(N52581));
    NANDX1 U39710 (.A1(n46698), .A2(N1724), .ZN(N52582));
    NANDX1 U39711 (.A1(n36007), .A2(N11448), .ZN(N52583));
    INVX1 U39712 (.I(n25344), .ZN(N52584));
    NANDX1 U39713 (.A1(n48719), .A2(n15856), .ZN(N52585));
    NANDX1 U39714 (.A1(N12155), .A2(N3127), .ZN(N52586));
    NOR2X1 U39715 (.A1(N5525), .A2(n46652), .ZN(N52587));
    NOR2X1 U39716 (.A1(n47022), .A2(n14851), .ZN(N52588));
    INVX1 U39717 (.I(n49332), .ZN(N52589));
    INVX1 U39718 (.I(N3213), .ZN(N52590));
    NANDX1 U39719 (.A1(n15270), .A2(n44663), .ZN(N52591));
    NOR2X1 U39720 (.A1(n34824), .A2(n37880), .ZN(N52592));
    NANDX1 U39721 (.A1(n40029), .A2(n32989), .ZN(N52593));
    INVX1 U39722 (.I(n20332), .ZN(N52594));
    NANDX1 U39723 (.A1(n15834), .A2(n13152), .ZN(N52595));
    NOR2X1 U39724 (.A1(N10367), .A2(n31898), .ZN(N52596));
    NOR2X1 U39725 (.A1(N10945), .A2(n14081), .ZN(N52597));
    NANDX1 U39726 (.A1(n24184), .A2(n19605), .ZN(N52598));
    NOR2X1 U39727 (.A1(N8629), .A2(n15039), .ZN(N52599));
    INVX1 U39728 (.I(N4784), .ZN(N52600));
    NOR2X1 U39729 (.A1(n50112), .A2(N7996), .ZN(N52601));
    NANDX1 U39730 (.A1(n13793), .A2(N1071), .ZN(N52602));
    NANDX1 U39731 (.A1(n18645), .A2(N8978), .ZN(N52603));
    INVX1 U39732 (.I(N7085), .ZN(N52604));
    NOR2X1 U39733 (.A1(n37947), .A2(n49032), .ZN(n52605));
    NANDX1 U39734 (.A1(n23808), .A2(n32211), .ZN(N52606));
    NANDX1 U39735 (.A1(n34175), .A2(N12521), .ZN(n52607));
    NOR2X1 U39736 (.A1(n15147), .A2(n26601), .ZN(N52608));
    INVX1 U39737 (.I(N9358), .ZN(N52609));
    NOR2X1 U39738 (.A1(n36028), .A2(n17986), .ZN(N52610));
    NOR2X1 U39739 (.A1(N9402), .A2(n22770), .ZN(N52611));
    NANDX1 U39740 (.A1(n29541), .A2(N793), .ZN(n52612));
    NANDX1 U39741 (.A1(n43333), .A2(n23479), .ZN(N52613));
    NOR2X1 U39742 (.A1(n32005), .A2(n32457), .ZN(N52614));
    INVX1 U39743 (.I(N9117), .ZN(N52615));
    NOR2X1 U39744 (.A1(n44584), .A2(n28177), .ZN(N52616));
    NANDX1 U39745 (.A1(n16804), .A2(N8799), .ZN(N52617));
    INVX1 U39746 (.I(n21006), .ZN(N52618));
    NANDX1 U39747 (.A1(n41886), .A2(n36152), .ZN(N52619));
    NANDX1 U39748 (.A1(N7858), .A2(n45510), .ZN(N52620));
    NANDX1 U39749 (.A1(n13913), .A2(n33523), .ZN(N52621));
    INVX1 U39750 (.I(n23314), .ZN(N52622));
    INVX1 U39751 (.I(N11230), .ZN(N52623));
    INVX1 U39752 (.I(n27113), .ZN(N52624));
    NANDX1 U39753 (.A1(n36243), .A2(n50591), .ZN(N52625));
    NANDX1 U39754 (.A1(n16659), .A2(N1487), .ZN(N52626));
    NOR2X1 U39755 (.A1(n25776), .A2(n45937), .ZN(N52627));
    INVX1 U39756 (.I(n23980), .ZN(N52628));
    INVX1 U39757 (.I(n16130), .ZN(N52629));
    NOR2X1 U39758 (.A1(n47629), .A2(n37135), .ZN(N52630));
    NOR2X1 U39759 (.A1(N7954), .A2(n43314), .ZN(N52631));
    INVX1 U39760 (.I(n15811), .ZN(N52632));
    NOR2X1 U39761 (.A1(N7950), .A2(n51339), .ZN(N52633));
    INVX1 U39762 (.I(n35072), .ZN(N52634));
    NANDX1 U39763 (.A1(n15517), .A2(n46301), .ZN(n52635));
    NANDX1 U39764 (.A1(N12657), .A2(n21328), .ZN(N52636));
    INVX1 U39765 (.I(n33276), .ZN(N52637));
    NOR2X1 U39766 (.A1(n17287), .A2(n34762), .ZN(N52638));
    NANDX1 U39767 (.A1(n13090), .A2(n50727), .ZN(N52639));
    NANDX1 U39768 (.A1(n37069), .A2(n29010), .ZN(N52640));
    INVX1 U39769 (.I(n39874), .ZN(N52641));
    INVX1 U39770 (.I(N6736), .ZN(N52642));
    NOR2X1 U39771 (.A1(N3031), .A2(n20078), .ZN(N52643));
    NANDX1 U39772 (.A1(n18841), .A2(n27340), .ZN(N52644));
    INVX1 U39773 (.I(n18591), .ZN(N52645));
    NANDX1 U39774 (.A1(n29201), .A2(N11683), .ZN(N52646));
    NOR2X1 U39775 (.A1(n45529), .A2(n49273), .ZN(N52647));
    NOR2X1 U39776 (.A1(n36884), .A2(n49900), .ZN(N52648));
    NANDX1 U39777 (.A1(N6316), .A2(n15598), .ZN(N52649));
    INVX1 U39778 (.I(N12051), .ZN(N52650));
    NANDX1 U39779 (.A1(n43585), .A2(n17111), .ZN(N52651));
    NOR2X1 U39780 (.A1(n21006), .A2(n38301), .ZN(N52652));
    INVX1 U39781 (.I(n37699), .ZN(N52653));
    INVX1 U39782 (.I(n49738), .ZN(N52654));
    INVX1 U39783 (.I(n35141), .ZN(N52655));
    NANDX1 U39784 (.A1(n29597), .A2(n32509), .ZN(N52656));
    NOR2X1 U39785 (.A1(n18215), .A2(n19073), .ZN(N52657));
    NANDX1 U39786 (.A1(n29898), .A2(n42770), .ZN(N52658));
    INVX1 U39787 (.I(n27582), .ZN(N52659));
    NANDX1 U39788 (.A1(n30128), .A2(n47509), .ZN(n52660));
    NOR2X1 U39789 (.A1(n36444), .A2(n33135), .ZN(N52661));
    INVX1 U39790 (.I(n18522), .ZN(N52662));
    INVX1 U39791 (.I(n30430), .ZN(N52663));
    NANDX1 U39792 (.A1(N7688), .A2(n21463), .ZN(N52664));
    INVX1 U39793 (.I(n23400), .ZN(N52665));
    INVX1 U39794 (.I(n29052), .ZN(N52666));
    NOR2X1 U39795 (.A1(n48301), .A2(n34220), .ZN(N52667));
    NOR2X1 U39796 (.A1(n26309), .A2(n15140), .ZN(N52668));
    NOR2X1 U39797 (.A1(n44524), .A2(n34213), .ZN(N52669));
    INVX1 U39798 (.I(n44449), .ZN(N52670));
    NANDX1 U39799 (.A1(n20117), .A2(n42058), .ZN(N52671));
    NOR2X1 U39800 (.A1(n50245), .A2(n37978), .ZN(N52672));
    INVX1 U39801 (.I(N5128), .ZN(N52673));
    INVX1 U39802 (.I(N3790), .ZN(N52674));
    NOR2X1 U39803 (.A1(n21401), .A2(N4248), .ZN(N52675));
    INVX1 U39804 (.I(n50704), .ZN(N52676));
    NOR2X1 U39805 (.A1(n43296), .A2(n22515), .ZN(N52677));
    NANDX1 U39806 (.A1(n20759), .A2(n14091), .ZN(N52678));
    NANDX1 U39807 (.A1(N3390), .A2(n41585), .ZN(N52679));
    NANDX1 U39808 (.A1(n18530), .A2(n17566), .ZN(N52680));
    NOR2X1 U39809 (.A1(n22770), .A2(n44439), .ZN(N52681));
    INVX1 U39810 (.I(n48163), .ZN(N52682));
    INVX1 U39811 (.I(n37472), .ZN(N52683));
    INVX1 U39812 (.I(n33239), .ZN(N52684));
    NOR2X1 U39813 (.A1(n36476), .A2(n38366), .ZN(N52685));
    INVX1 U39814 (.I(N10293), .ZN(N52686));
    NANDX1 U39815 (.A1(n26457), .A2(n14540), .ZN(N52687));
    NOR2X1 U39816 (.A1(n25572), .A2(N10278), .ZN(N52688));
    NOR2X1 U39817 (.A1(n48086), .A2(n13588), .ZN(N52689));
    NANDX1 U39818 (.A1(N10588), .A2(n35226), .ZN(N52690));
    NANDX1 U39819 (.A1(n22201), .A2(N1613), .ZN(N52691));
    INVX1 U39820 (.I(N9794), .ZN(N52692));
    INVX1 U39821 (.I(n50202), .ZN(N52693));
    INVX1 U39822 (.I(N7937), .ZN(N52694));
    INVX1 U39823 (.I(n37227), .ZN(N52695));
    INVX1 U39824 (.I(n14720), .ZN(N52696));
    INVX1 U39825 (.I(N9325), .ZN(N52697));
    INVX1 U39826 (.I(n27271), .ZN(N52698));
    NANDX1 U39827 (.A1(n31515), .A2(N7724), .ZN(N52699));
    INVX1 U39828 (.I(n46055), .ZN(N52700));
    NANDX1 U39829 (.A1(n14820), .A2(N4744), .ZN(N52701));
    INVX1 U39830 (.I(n32933), .ZN(N52702));
    INVX1 U39831 (.I(n46083), .ZN(N52703));
    NOR2X1 U39832 (.A1(n23584), .A2(n33371), .ZN(N52704));
    INVX1 U39833 (.I(n25197), .ZN(N52705));
    NANDX1 U39834 (.A1(n15570), .A2(N7747), .ZN(N52706));
    NANDX1 U39835 (.A1(n18213), .A2(n15684), .ZN(N52707));
    NOR2X1 U39836 (.A1(N3851), .A2(n31119), .ZN(N52708));
    NANDX1 U39837 (.A1(n44344), .A2(N10471), .ZN(N52709));
    NANDX1 U39838 (.A1(n20026), .A2(n24851), .ZN(N52710));
    INVX1 U39839 (.I(n49365), .ZN(N52711));
    NANDX1 U39840 (.A1(n26610), .A2(n36878), .ZN(N52712));
    NANDX1 U39841 (.A1(n31353), .A2(n17502), .ZN(N52713));
    INVX1 U39842 (.I(n19711), .ZN(N52714));
    INVX1 U39843 (.I(n15454), .ZN(N52715));
    NANDX1 U39844 (.A1(n15395), .A2(n21229), .ZN(N52716));
    INVX1 U39845 (.I(n46225), .ZN(N52717));
    INVX1 U39846 (.I(n24649), .ZN(N52718));
    NOR2X1 U39847 (.A1(n25039), .A2(N10360), .ZN(N52719));
    NANDX1 U39848 (.A1(n50505), .A2(N11507), .ZN(N52720));
    NOR2X1 U39849 (.A1(n13288), .A2(n21977), .ZN(N52721));
    INVX1 U39850 (.I(N3341), .ZN(N52722));
    INVX1 U39851 (.I(n17661), .ZN(N52723));
    NANDX1 U39852 (.A1(n30954), .A2(n44270), .ZN(N52724));
    INVX1 U39853 (.I(n51516), .ZN(N52725));
    NOR2X1 U39854 (.A1(n47140), .A2(N1833), .ZN(N52726));
    NOR2X1 U39855 (.A1(n29164), .A2(n38902), .ZN(N52727));
    NANDX1 U39856 (.A1(n14586), .A2(n30159), .ZN(N52728));
    NOR2X1 U39857 (.A1(N9223), .A2(n36984), .ZN(N52729));
    INVX1 U39858 (.I(n33303), .ZN(N52730));
    INVX1 U39859 (.I(n19061), .ZN(N52731));
    NOR2X1 U39860 (.A1(n30967), .A2(n30567), .ZN(N52732));
    NOR2X1 U39861 (.A1(n14282), .A2(N956), .ZN(N52733));
    NANDX1 U39862 (.A1(n17623), .A2(n17811), .ZN(N52734));
    INVX1 U39863 (.I(n40356), .ZN(N52735));
    NOR2X1 U39864 (.A1(n16077), .A2(n48378), .ZN(N52736));
    NANDX1 U39865 (.A1(N10139), .A2(n13957), .ZN(N52737));
    NANDX1 U39866 (.A1(n45528), .A2(n13149), .ZN(N52738));
    NANDX1 U39867 (.A1(n21034), .A2(n27734), .ZN(N52739));
    INVX1 U39868 (.I(N5087), .ZN(N52740));
    NOR2X1 U39869 (.A1(n45035), .A2(n43760), .ZN(N52741));
    INVX1 U39870 (.I(n25496), .ZN(N52742));
    INVX1 U39871 (.I(N10770), .ZN(N52743));
    NOR2X1 U39872 (.A1(N11827), .A2(n39344), .ZN(N52744));
    NANDX1 U39873 (.A1(n34398), .A2(n23463), .ZN(N52745));
    NOR2X1 U39874 (.A1(N620), .A2(n46858), .ZN(N52746));
    NANDX1 U39875 (.A1(n19411), .A2(N11347), .ZN(N52747));
    NANDX1 U39876 (.A1(n38130), .A2(n43101), .ZN(N52748));
    NANDX1 U39877 (.A1(n28709), .A2(n37040), .ZN(N52749));
    NANDX1 U39878 (.A1(n36573), .A2(n28102), .ZN(N52750));
    INVX1 U39879 (.I(n44624), .ZN(N52751));
    NANDX1 U39880 (.A1(n37471), .A2(n38070), .ZN(N52752));
    INVX1 U39881 (.I(n17813), .ZN(N52753));
    NANDX1 U39882 (.A1(n28234), .A2(n50198), .ZN(N52754));
    NANDX1 U39883 (.A1(n40060), .A2(n37954), .ZN(N52755));
    NOR2X1 U39884 (.A1(n44485), .A2(n31444), .ZN(N52756));
    NANDX1 U39885 (.A1(n45104), .A2(n48330), .ZN(N52757));
    INVX1 U39886 (.I(n34543), .ZN(N52758));
    INVX1 U39887 (.I(n48908), .ZN(N52759));
    INVX1 U39888 (.I(n21216), .ZN(N52760));
    INVX1 U39889 (.I(n19820), .ZN(N52761));
    NANDX1 U39890 (.A1(n49623), .A2(N4804), .ZN(N52762));
    NOR2X1 U39891 (.A1(n28522), .A2(n19455), .ZN(N52763));
    INVX1 U39892 (.I(n14404), .ZN(N52764));
    NOR2X1 U39893 (.A1(n33370), .A2(N2245), .ZN(N52765));
    NANDX1 U39894 (.A1(n31631), .A2(N854), .ZN(N52766));
    INVX1 U39895 (.I(n41719), .ZN(N52767));
    NOR2X1 U39896 (.A1(n37344), .A2(n34615), .ZN(N52768));
    INVX1 U39897 (.I(n33470), .ZN(N52769));
    INVX1 U39898 (.I(N7048), .ZN(N52770));
    NANDX1 U39899 (.A1(n32701), .A2(n36751), .ZN(N52771));
    INVX1 U39900 (.I(n23812), .ZN(N52772));
    NOR2X1 U39901 (.A1(n31027), .A2(n43631), .ZN(N52773));
    NANDX1 U39902 (.A1(n29061), .A2(n18462), .ZN(N52774));
    INVX1 U39903 (.I(n27610), .ZN(N52775));
    NOR2X1 U39904 (.A1(n25852), .A2(N12042), .ZN(N52776));
    NOR2X1 U39905 (.A1(n29249), .A2(n14286), .ZN(N52777));
    INVX1 U39906 (.I(N9292), .ZN(N52778));
    INVX1 U39907 (.I(n33130), .ZN(N52779));
    NANDX1 U39908 (.A1(n23974), .A2(n40501), .ZN(N52780));
    NANDX1 U39909 (.A1(n34280), .A2(n43998), .ZN(N52781));
    NANDX1 U39910 (.A1(n41327), .A2(N9221), .ZN(N52782));
    NANDX1 U39911 (.A1(n26489), .A2(n44967), .ZN(N52783));
    NOR2X1 U39912 (.A1(N2894), .A2(n24406), .ZN(N52784));
    INVX1 U39913 (.I(n37555), .ZN(N52785));
    INVX1 U39914 (.I(n39265), .ZN(N52786));
    INVX1 U39915 (.I(n51104), .ZN(N52787));
    INVX1 U39916 (.I(n21303), .ZN(N52788));
    INVX1 U39917 (.I(N1144), .ZN(N52789));
    INVX1 U39918 (.I(n25842), .ZN(N52790));
    NOR2X1 U39919 (.A1(n29870), .A2(n40980), .ZN(N52791));
    NOR2X1 U39920 (.A1(n50907), .A2(n34981), .ZN(N52792));
    NANDX1 U39921 (.A1(n24999), .A2(n17672), .ZN(N52793));
    NANDX1 U39922 (.A1(n27220), .A2(N7410), .ZN(N52794));
    NANDX1 U39923 (.A1(n32170), .A2(N3926), .ZN(N52795));
    INVX1 U39924 (.I(N9342), .ZN(N52796));
    INVX1 U39925 (.I(n19351), .ZN(N52797));
    NANDX1 U39926 (.A1(n14402), .A2(n12873), .ZN(N52798));
    NANDX1 U39927 (.A1(n39824), .A2(N12388), .ZN(n52799));
    NOR2X1 U39928 (.A1(N9538), .A2(n45560), .ZN(N52800));
    NOR2X1 U39929 (.A1(n30117), .A2(n41429), .ZN(N52801));
    NANDX1 U39930 (.A1(N8398), .A2(N848), .ZN(N52802));
    NOR2X1 U39931 (.A1(n29333), .A2(n35829), .ZN(N52803));
    NANDX1 U39932 (.A1(N2743), .A2(N1912), .ZN(N52804));
    INVX1 U39933 (.I(n29962), .ZN(N52805));
    NANDX1 U39934 (.A1(n14066), .A2(n32159), .ZN(N52806));
    INVX1 U39935 (.I(N9012), .ZN(N52807));
    NANDX1 U39936 (.A1(n33326), .A2(n49978), .ZN(N52808));
    NOR2X1 U39937 (.A1(n47727), .A2(N11262), .ZN(N52809));
    NANDX1 U39938 (.A1(n35963), .A2(n45265), .ZN(N52810));
    NANDX1 U39939 (.A1(n15528), .A2(N9264), .ZN(N52811));
    NANDX1 U39940 (.A1(n45644), .A2(n50692), .ZN(N52812));
    INVX1 U39941 (.I(n24070), .ZN(n52813));
    NOR2X1 U39942 (.A1(n36814), .A2(N1814), .ZN(N52814));
    NOR2X1 U39943 (.A1(N5378), .A2(N4556), .ZN(N52815));
    NOR2X1 U39944 (.A1(n39492), .A2(N4545), .ZN(N52816));
    NANDX1 U39945 (.A1(N1970), .A2(n36704), .ZN(N52817));
    NOR2X1 U39946 (.A1(N10981), .A2(n48232), .ZN(N52818));
    INVX1 U39947 (.I(N9370), .ZN(N52819));
    INVX1 U39948 (.I(n13067), .ZN(N52820));
    NANDX1 U39949 (.A1(N7892), .A2(n49029), .ZN(N52821));
    NOR2X1 U39950 (.A1(N4168), .A2(n34584), .ZN(N52822));
    NOR2X1 U39951 (.A1(N6671), .A2(n28640), .ZN(N52823));
    NOR2X1 U39952 (.A1(n31625), .A2(N1121), .ZN(N52824));
    NOR2X1 U39953 (.A1(n38466), .A2(n24550), .ZN(N52825));
    NANDX1 U39954 (.A1(n13871), .A2(n29105), .ZN(N52826));
    NOR2X1 U39955 (.A1(N1775), .A2(n33649), .ZN(N52827));
    INVX1 U39956 (.I(N3744), .ZN(N52828));
    NOR2X1 U39957 (.A1(N11725), .A2(n36340), .ZN(N52829));
    NOR2X1 U39958 (.A1(n28653), .A2(n15737), .ZN(N52830));
    NOR2X1 U39959 (.A1(n41719), .A2(N6396), .ZN(N52831));
    NANDX1 U39960 (.A1(n39159), .A2(n33964), .ZN(N52832));
    NANDX1 U39961 (.A1(n43770), .A2(n49179), .ZN(N52833));
    INVX1 U39962 (.I(n20821), .ZN(N52834));
    NOR2X1 U39963 (.A1(n35775), .A2(n43557), .ZN(N52835));
    NOR2X1 U39964 (.A1(n22653), .A2(n16518), .ZN(N52836));
    INVX1 U39965 (.I(N6551), .ZN(n52837));
    INVX1 U39966 (.I(n27366), .ZN(N52838));
    NOR2X1 U39967 (.A1(n49299), .A2(n25517), .ZN(N52839));
    NOR2X1 U39968 (.A1(N8118), .A2(n37241), .ZN(N52840));
    NOR2X1 U39969 (.A1(n45141), .A2(n14305), .ZN(N52841));
    NOR2X1 U39970 (.A1(N8946), .A2(N4435), .ZN(N52842));
    NOR2X1 U39971 (.A1(n32231), .A2(n13621), .ZN(N52843));
    NOR2X1 U39972 (.A1(n29710), .A2(N5803), .ZN(N52844));
    NANDX1 U39973 (.A1(n33860), .A2(n48239), .ZN(N52845));
    NANDX1 U39974 (.A1(n18047), .A2(N10236), .ZN(N52846));
    NANDX1 U39975 (.A1(N10727), .A2(n26753), .ZN(N52847));
    NANDX1 U39976 (.A1(n17277), .A2(n42403), .ZN(N52848));
    NOR2X1 U39977 (.A1(n47218), .A2(N10141), .ZN(N52849));
    INVX1 U39978 (.I(n29313), .ZN(N52850));
    NOR2X1 U39979 (.A1(n20067), .A2(n17776), .ZN(N52851));
    NANDX1 U39980 (.A1(N4400), .A2(n21975), .ZN(N52852));
    NOR2X1 U39981 (.A1(n30450), .A2(N2597), .ZN(N52853));
    NANDX1 U39982 (.A1(n14099), .A2(n38799), .ZN(N52854));
    NANDX1 U39983 (.A1(n41517), .A2(n50974), .ZN(N52855));
    INVX1 U39984 (.I(n38167), .ZN(N52856));
    NOR2X1 U39985 (.A1(n23069), .A2(n48402), .ZN(N52857));
    INVX1 U39986 (.I(N3823), .ZN(N52858));
    NOR2X1 U39987 (.A1(N8581), .A2(n42715), .ZN(N52859));
    NOR2X1 U39988 (.A1(n47451), .A2(n38344), .ZN(N52860));
    NOR2X1 U39989 (.A1(n30277), .A2(n37685), .ZN(N52861));
    NOR2X1 U39990 (.A1(n20371), .A2(n25488), .ZN(N52862));
    NOR2X1 U39991 (.A1(n46386), .A2(n17490), .ZN(N52863));
    NANDX1 U39992 (.A1(n25248), .A2(n41702), .ZN(N52864));
    NOR2X1 U39993 (.A1(n39346), .A2(n28912), .ZN(N52865));
    INVX1 U39994 (.I(n50890), .ZN(N52866));
    NOR2X1 U39995 (.A1(n49472), .A2(n37468), .ZN(N52867));
    NANDX1 U39996 (.A1(n42568), .A2(N4310), .ZN(N52868));
    INVX1 U39997 (.I(n46390), .ZN(N52869));
    INVX1 U39998 (.I(N10739), .ZN(N52870));
    NANDX1 U39999 (.A1(N3928), .A2(n28217), .ZN(N52871));
    NOR2X1 U40000 (.A1(n20092), .A2(n28521), .ZN(N52872));
    NANDX1 U40001 (.A1(N2925), .A2(n48891), .ZN(N52873));
    INVX1 U40002 (.I(n19184), .ZN(N52874));
    NOR2X1 U40003 (.A1(n44988), .A2(n26226), .ZN(N52875));
    NOR2X1 U40004 (.A1(n35102), .A2(n26309), .ZN(N52876));
    INVX1 U40005 (.I(N12425), .ZN(N52877));
    INVX1 U40006 (.I(n47638), .ZN(N52878));
    NANDX1 U40007 (.A1(n17054), .A2(N3545), .ZN(N52879));
    NANDX1 U40008 (.A1(N8034), .A2(N7854), .ZN(N52880));
    NANDX1 U40009 (.A1(n24451), .A2(n27373), .ZN(n52881));
    NOR2X1 U40010 (.A1(n31995), .A2(n31300), .ZN(N52882));
    NANDX1 U40011 (.A1(n26295), .A2(n51391), .ZN(N52883));
    INVX1 U40012 (.I(n49922), .ZN(N52884));
    NANDX1 U40013 (.A1(n31179), .A2(n25833), .ZN(N52885));
    NOR2X1 U40014 (.A1(n44895), .A2(n40848), .ZN(N52886));
    NOR2X1 U40015 (.A1(N2298), .A2(n24361), .ZN(N52887));
    NANDX1 U40016 (.A1(n20662), .A2(N6814), .ZN(N52888));
    NOR2X1 U40017 (.A1(n16711), .A2(n39179), .ZN(N52889));
    NOR2X1 U40018 (.A1(n41872), .A2(N3423), .ZN(N52890));
    NOR2X1 U40019 (.A1(n19753), .A2(n21413), .ZN(N52891));
    NOR2X1 U40020 (.A1(n47126), .A2(n50141), .ZN(N52892));
    NOR2X1 U40021 (.A1(n48453), .A2(N3909), .ZN(N52893));
    NOR2X1 U40022 (.A1(n18284), .A2(n37785), .ZN(N52894));
    INVX1 U40023 (.I(n42627), .ZN(N52895));
    INVX1 U40024 (.I(n15802), .ZN(N52896));
    NANDX1 U40025 (.A1(N2326), .A2(N5062), .ZN(N52897));
    NANDX1 U40026 (.A1(n26240), .A2(n51038), .ZN(N52898));
    NANDX1 U40027 (.A1(n46901), .A2(N6263), .ZN(N52899));
    INVX1 U40028 (.I(N12024), .ZN(N52900));
    NANDX1 U40029 (.A1(N1764), .A2(n23923), .ZN(N52901));
    NANDX1 U40030 (.A1(n22193), .A2(n43675), .ZN(N52902));
    NANDX1 U40031 (.A1(n37101), .A2(n39212), .ZN(N52903));
    NOR2X1 U40032 (.A1(n32415), .A2(N6105), .ZN(N52904));
    INVX1 U40033 (.I(n24051), .ZN(N52905));
    INVX1 U40034 (.I(N12250), .ZN(N52906));
    NOR2X1 U40035 (.A1(n15426), .A2(n51241), .ZN(N52907));
    NANDX1 U40036 (.A1(n49990), .A2(n23595), .ZN(N52908));
    NOR2X1 U40037 (.A1(n21159), .A2(n49834), .ZN(N52909));
    INVX1 U40038 (.I(n28444), .ZN(N52910));
    NANDX1 U40039 (.A1(n32239), .A2(N9455), .ZN(N52911));
    NANDX1 U40040 (.A1(n17736), .A2(n32835), .ZN(N52912));
    NANDX1 U40041 (.A1(N6655), .A2(N3439), .ZN(N52913));
    INVX1 U40042 (.I(n38603), .ZN(N52914));
    INVX1 U40043 (.I(N857), .ZN(N52915));
    NOR2X1 U40044 (.A1(n42981), .A2(N6961), .ZN(N52916));
    NOR2X1 U40045 (.A1(n15443), .A2(N1376), .ZN(N52917));
    INVX1 U40046 (.I(n29463), .ZN(N52918));
    INVX1 U40047 (.I(n25499), .ZN(N52919));
    NANDX1 U40048 (.A1(n15203), .A2(n19121), .ZN(N52920));
    INVX1 U40049 (.I(N6389), .ZN(N52921));
    NANDX1 U40050 (.A1(n38581), .A2(N4860), .ZN(N52922));
    INVX1 U40051 (.I(n40847), .ZN(N52923));
    INVX1 U40052 (.I(N8148), .ZN(N52924));
    INVX1 U40053 (.I(n17176), .ZN(N52925));
    NANDX1 U40054 (.A1(n13649), .A2(n42231), .ZN(N52926));
    NANDX1 U40055 (.A1(n22279), .A2(N1209), .ZN(N52927));
    NANDX1 U40056 (.A1(N9822), .A2(n14218), .ZN(N52928));
    NOR2X1 U40057 (.A1(n23418), .A2(n29660), .ZN(N52929));
    NANDX1 U40058 (.A1(n49264), .A2(n29150), .ZN(N52930));
    NOR2X1 U40059 (.A1(n44790), .A2(N6873), .ZN(N52931));
    INVX1 U40060 (.I(n33938), .ZN(N52932));
    INVX1 U40061 (.I(n21810), .ZN(N52933));
    NOR2X1 U40062 (.A1(n19731), .A2(n48285), .ZN(N52934));
    INVX1 U40063 (.I(N8989), .ZN(N52935));
    NANDX1 U40064 (.A1(n32044), .A2(n37599), .ZN(N52936));
    NANDX1 U40065 (.A1(N9750), .A2(n21275), .ZN(N52937));
    INVX1 U40066 (.I(n22304), .ZN(N52938));
    NANDX1 U40067 (.A1(n41653), .A2(N5743), .ZN(n52939));
    NOR2X1 U40068 (.A1(n25898), .A2(n17759), .ZN(N52940));
    NOR2X1 U40069 (.A1(N3969), .A2(n31150), .ZN(N52941));
    INVX1 U40070 (.I(N3147), .ZN(N52942));
    NOR2X1 U40071 (.A1(n29340), .A2(n31635), .ZN(N52943));
    NANDX1 U40072 (.A1(N11689), .A2(N12785), .ZN(N52944));
    INVX1 U40073 (.I(n33019), .ZN(N52945));
    INVX1 U40074 (.I(n13709), .ZN(N52946));
    NANDX1 U40075 (.A1(N11531), .A2(n46335), .ZN(N52947));
    NOR2X1 U40076 (.A1(n49129), .A2(n14576), .ZN(N52948));
    NANDX1 U40077 (.A1(n18815), .A2(N3432), .ZN(N52949));
    NANDX1 U40078 (.A1(N10780), .A2(n15112), .ZN(N52950));
    NOR2X1 U40079 (.A1(N4210), .A2(n41009), .ZN(N52951));
    INVX1 U40080 (.I(n21057), .ZN(N52952));
    NANDX1 U40081 (.A1(N12541), .A2(N5608), .ZN(N52953));
    NANDX1 U40082 (.A1(n22294), .A2(N4975), .ZN(N52954));
    NANDX1 U40083 (.A1(n17496), .A2(n38280), .ZN(N52955));
    NOR2X1 U40084 (.A1(n34507), .A2(n41326), .ZN(N52956));
    INVX1 U40085 (.I(n48215), .ZN(N52957));
    NOR2X1 U40086 (.A1(n46670), .A2(n42961), .ZN(N52958));
    NOR2X1 U40087 (.A1(n44211), .A2(n27565), .ZN(N52959));
    NANDX1 U40088 (.A1(n33053), .A2(n30996), .ZN(N52960));
    INVX1 U40089 (.I(n13860), .ZN(N52961));
    NOR2X1 U40090 (.A1(n22696), .A2(n18069), .ZN(N52962));
    NANDX1 U40091 (.A1(n25703), .A2(N9154), .ZN(N52963));
    NOR2X1 U40092 (.A1(n38244), .A2(n36377), .ZN(N52964));
    NOR2X1 U40093 (.A1(n30565), .A2(n41351), .ZN(N52965));
    INVX1 U40094 (.I(n48060), .ZN(n52966));
    NANDX1 U40095 (.A1(N1204), .A2(n30978), .ZN(N52967));
    NOR2X1 U40096 (.A1(n36343), .A2(n49221), .ZN(N52968));
    NOR2X1 U40097 (.A1(N1452), .A2(N10621), .ZN(N52969));
    NANDX1 U40098 (.A1(n15690), .A2(n38185), .ZN(N52970));
    INVX1 U40099 (.I(n48743), .ZN(N52971));
    NOR2X1 U40100 (.A1(n42391), .A2(N11014), .ZN(N52972));
    NOR2X1 U40101 (.A1(n35114), .A2(n29083), .ZN(N52973));
    NANDX1 U40102 (.A1(N9229), .A2(n38236), .ZN(N52974));
    NOR2X1 U40103 (.A1(n17500), .A2(n44640), .ZN(N52975));
    NANDX1 U40104 (.A1(n18092), .A2(n34402), .ZN(N52976));
    NOR2X1 U40105 (.A1(n36179), .A2(N2500), .ZN(N52977));
    NOR2X1 U40106 (.A1(n37184), .A2(N11923), .ZN(N52978));
    INVX1 U40107 (.I(n34816), .ZN(N52979));
    NOR2X1 U40108 (.A1(n29494), .A2(n45437), .ZN(N52980));
    NANDX1 U40109 (.A1(n45184), .A2(N2061), .ZN(N52981));
    NOR2X1 U40110 (.A1(n42338), .A2(n41269), .ZN(N52982));
    INVX1 U40111 (.I(N1763), .ZN(N52983));
    NOR2X1 U40112 (.A1(n24250), .A2(N873), .ZN(N52984));
    NOR2X1 U40113 (.A1(n33478), .A2(N9136), .ZN(N52985));
    NANDX1 U40114 (.A1(n21005), .A2(N2187), .ZN(N52986));
    NOR2X1 U40115 (.A1(n39096), .A2(N6617), .ZN(N52987));
    NANDX1 U40116 (.A1(n45302), .A2(N9116), .ZN(N52988));
    NANDX1 U40117 (.A1(n30897), .A2(n42654), .ZN(N52989));
    NOR2X1 U40118 (.A1(n35741), .A2(N7475), .ZN(N52990));
    NOR2X1 U40119 (.A1(n29589), .A2(n30835), .ZN(N52991));
    NOR2X1 U40120 (.A1(N1677), .A2(N7552), .ZN(N52992));
    NANDX1 U40121 (.A1(n42945), .A2(n48276), .ZN(N52993));
    NANDX1 U40122 (.A1(n36379), .A2(n20937), .ZN(N52994));
    INVX1 U40123 (.I(n39120), .ZN(N52995));
    INVX1 U40124 (.I(n17142), .ZN(N52996));
    INVX1 U40125 (.I(n45446), .ZN(N52997));
    NOR2X1 U40126 (.A1(n44665), .A2(N2981), .ZN(N52998));
    INVX1 U40127 (.I(n24812), .ZN(N52999));
    NOR2X1 U40128 (.A1(n26703), .A2(n48247), .ZN(N53000));
    NOR2X1 U40129 (.A1(n17768), .A2(n48136), .ZN(N53001));
    INVX1 U40130 (.I(n25243), .ZN(N53002));
    NOR2X1 U40131 (.A1(n32974), .A2(n26105), .ZN(N53003));
    INVX1 U40132 (.I(n34651), .ZN(N53004));
    NOR2X1 U40133 (.A1(N11046), .A2(n26007), .ZN(N53005));
    NANDX1 U40134 (.A1(n48151), .A2(N10797), .ZN(N53006));
    NANDX1 U40135 (.A1(N4569), .A2(n49916), .ZN(N53007));
    NANDX1 U40136 (.A1(n43326), .A2(N10110), .ZN(N53008));
    INVX1 U40137 (.I(n32681), .ZN(N53009));
    NOR2X1 U40138 (.A1(n34230), .A2(n50269), .ZN(N53010));
    NANDX1 U40139 (.A1(N951), .A2(n25383), .ZN(N53011));
    NANDX1 U40140 (.A1(n50156), .A2(n13179), .ZN(N53012));
    NANDX1 U40141 (.A1(n31926), .A2(N8449), .ZN(N53013));
    NOR2X1 U40142 (.A1(n34927), .A2(n34553), .ZN(N53014));
    INVX1 U40143 (.I(n39605), .ZN(N53015));
    NANDX1 U40144 (.A1(n25524), .A2(n14024), .ZN(N53016));
    INVX1 U40145 (.I(n43703), .ZN(N53017));
    NANDX1 U40146 (.A1(N8327), .A2(n18299), .ZN(N53018));
    NANDX1 U40147 (.A1(n24103), .A2(N10036), .ZN(N53019));
    NANDX1 U40148 (.A1(n33736), .A2(N12744), .ZN(N53020));
    NANDX1 U40149 (.A1(n16377), .A2(N11424), .ZN(N53021));
    NOR2X1 U40150 (.A1(n17327), .A2(N6835), .ZN(N53022));
    NOR2X1 U40151 (.A1(n37511), .A2(n20013), .ZN(n53023));
    NANDX1 U40152 (.A1(n39464), .A2(n28461), .ZN(N53024));
    NANDX1 U40153 (.A1(n22802), .A2(n33041), .ZN(N53025));
    NOR2X1 U40154 (.A1(N10819), .A2(n19690), .ZN(N53026));
    NOR2X1 U40155 (.A1(n46458), .A2(N6709), .ZN(n53027));
    NANDX1 U40156 (.A1(N11333), .A2(n36652), .ZN(N53028));
    NOR2X1 U40157 (.A1(n47740), .A2(N9166), .ZN(N53029));
    INVX1 U40158 (.I(n42669), .ZN(N53030));
    NOR2X1 U40159 (.A1(n47334), .A2(n40783), .ZN(N53031));
    NANDX1 U40160 (.A1(N7170), .A2(N6949), .ZN(N53032));
    NANDX1 U40161 (.A1(n14004), .A2(n41002), .ZN(N53033));
    INVX1 U40162 (.I(N4044), .ZN(N53034));
    NOR2X1 U40163 (.A1(N12074), .A2(n32504), .ZN(N53035));
    NANDX1 U40164 (.A1(n34875), .A2(n35572), .ZN(N53036));
    NANDX1 U40165 (.A1(n15721), .A2(n25289), .ZN(N53037));
    NANDX1 U40166 (.A1(n32206), .A2(N2026), .ZN(N53038));
    NOR2X1 U40167 (.A1(n43539), .A2(n38677), .ZN(N53039));
    NOR2X1 U40168 (.A1(n39690), .A2(n17870), .ZN(N53040));
    INVX1 U40169 (.I(n30770), .ZN(N53041));
    INVX1 U40170 (.I(n47844), .ZN(N53042));
    NOR2X1 U40171 (.A1(n30133), .A2(n25041), .ZN(N53043));
    INVX1 U40172 (.I(n16821), .ZN(N53044));
    NANDX1 U40173 (.A1(n37942), .A2(n41019), .ZN(N53045));
    NANDX1 U40174 (.A1(n22666), .A2(N1504), .ZN(N53046));
    INVX1 U40175 (.I(n19860), .ZN(N53047));
    INVX1 U40176 (.I(n51218), .ZN(N53048));
    INVX1 U40177 (.I(n22127), .ZN(N53049));
    NOR2X1 U40178 (.A1(N725), .A2(N2744), .ZN(N53050));
    NOR2X1 U40179 (.A1(n45266), .A2(n16310), .ZN(N53051));
    INVX1 U40180 (.I(N11186), .ZN(N53052));
    NANDX1 U40181 (.A1(N1929), .A2(N11696), .ZN(N53053));
    INVX1 U40182 (.I(n32727), .ZN(N53054));
    INVX1 U40183 (.I(n46789), .ZN(N53055));
    NOR2X1 U40184 (.A1(n32992), .A2(n43729), .ZN(N53056));
    NANDX1 U40185 (.A1(n42063), .A2(N110), .ZN(N53057));
    NANDX1 U40186 (.A1(n25206), .A2(n22776), .ZN(N53058));
    NANDX1 U40187 (.A1(n40851), .A2(N12663), .ZN(N53059));
    NOR2X1 U40188 (.A1(n40480), .A2(n26691), .ZN(N53060));
    NANDX1 U40189 (.A1(n13810), .A2(n49031), .ZN(N53061));
    INVX1 U40190 (.I(N10780), .ZN(N53062));
    NOR2X1 U40191 (.A1(n49897), .A2(n46427), .ZN(N53063));
    NANDX1 U40192 (.A1(N2720), .A2(n48355), .ZN(N53064));
    NOR2X1 U40193 (.A1(n29544), .A2(n51109), .ZN(n53065));
    INVX1 U40194 (.I(n24744), .ZN(N53066));
    NANDX1 U40195 (.A1(n16613), .A2(n38500), .ZN(N53067));
    INVX1 U40196 (.I(n28704), .ZN(N53068));
    NOR2X1 U40197 (.A1(n18075), .A2(N2321), .ZN(N53069));
    NOR2X1 U40198 (.A1(N7126), .A2(n43171), .ZN(N53070));
    NANDX1 U40199 (.A1(n24199), .A2(n32063), .ZN(N53071));
    NANDX1 U40200 (.A1(n33426), .A2(n15900), .ZN(N53072));
    NOR2X1 U40201 (.A1(n15425), .A2(n26679), .ZN(N53073));
    NOR2X1 U40202 (.A1(n13733), .A2(n43133), .ZN(N53074));
    INVX1 U40203 (.I(n38068), .ZN(N53075));
    NOR2X1 U40204 (.A1(n28945), .A2(n16023), .ZN(n53076));
    INVX1 U40205 (.I(n42538), .ZN(N53077));
    NOR2X1 U40206 (.A1(n41855), .A2(N7563), .ZN(N53078));
    INVX1 U40207 (.I(n42408), .ZN(N53079));
    NANDX1 U40208 (.A1(N6343), .A2(N8894), .ZN(N53080));
    INVX1 U40209 (.I(n37755), .ZN(N53081));
    INVX1 U40210 (.I(N196), .ZN(N53082));
    NANDX1 U40211 (.A1(n31862), .A2(n32258), .ZN(N53083));
    NOR2X1 U40212 (.A1(n35316), .A2(n18185), .ZN(N53084));
    NOR2X1 U40213 (.A1(n50740), .A2(n14892), .ZN(N53085));
    NOR2X1 U40214 (.A1(n12884), .A2(N6436), .ZN(N53086));
    NOR2X1 U40215 (.A1(n50951), .A2(n16363), .ZN(N53087));
    INVX1 U40216 (.I(n15385), .ZN(N53088));
    NANDX1 U40217 (.A1(n31955), .A2(n26179), .ZN(N53089));
    INVX1 U40218 (.I(N9545), .ZN(N53090));
    NANDX1 U40219 (.A1(n50127), .A2(n15838), .ZN(N53091));
    NOR2X1 U40220 (.A1(n29049), .A2(n24451), .ZN(N53092));
    INVX1 U40221 (.I(n36712), .ZN(N53093));
    NANDX1 U40222 (.A1(N8306), .A2(n16985), .ZN(N53094));
    NANDX1 U40223 (.A1(n19395), .A2(N712), .ZN(N53095));
    NOR2X1 U40224 (.A1(n17129), .A2(n51451), .ZN(N53096));
    NANDX1 U40225 (.A1(N5889), .A2(n34362), .ZN(N53097));
    INVX1 U40226 (.I(n47921), .ZN(N53098));
    INVX1 U40227 (.I(n44477), .ZN(N53099));
    INVX1 U40228 (.I(n19137), .ZN(N53100));
    NOR2X1 U40229 (.A1(N9348), .A2(n45315), .ZN(N53101));
    INVX1 U40230 (.I(n40508), .ZN(N53102));
    NANDX1 U40231 (.A1(n38215), .A2(N4757), .ZN(N53103));
    NOR2X1 U40232 (.A1(n15675), .A2(n50823), .ZN(N53104));
    NOR2X1 U40233 (.A1(N798), .A2(n15524), .ZN(N53105));
    NANDX1 U40234 (.A1(n39399), .A2(N12483), .ZN(N53106));
    INVX1 U40235 (.I(n40110), .ZN(N53107));
    NOR2X1 U40236 (.A1(N2431), .A2(N10001), .ZN(N53108));
    NANDX1 U40237 (.A1(N8319), .A2(n44362), .ZN(N53109));
    NANDX1 U40238 (.A1(n26267), .A2(n48114), .ZN(N53110));
    INVX1 U40239 (.I(n33632), .ZN(N53111));
    NANDX1 U40240 (.A1(n37416), .A2(n13007), .ZN(N53112));
    NANDX1 U40241 (.A1(n25504), .A2(N1926), .ZN(N53113));
    NANDX1 U40242 (.A1(N12131), .A2(n28298), .ZN(N53114));
    INVX1 U40243 (.I(n49421), .ZN(N53115));
    NANDX1 U40244 (.A1(n15726), .A2(n50219), .ZN(N53116));
    INVX1 U40245 (.I(N11605), .ZN(N53117));
    INVX1 U40246 (.I(n25566), .ZN(N53118));
    NOR2X1 U40247 (.A1(n48166), .A2(N1604), .ZN(N53119));
    NOR2X1 U40248 (.A1(N6578), .A2(n50909), .ZN(N53120));
    NOR2X1 U40249 (.A1(n50940), .A2(n33507), .ZN(N53121));
    NANDX1 U40250 (.A1(n17493), .A2(N638), .ZN(N53122));
    INVX1 U40251 (.I(n33154), .ZN(N53123));
    INVX1 U40252 (.I(n42231), .ZN(N53124));
    NANDX1 U40253 (.A1(n33585), .A2(n44157), .ZN(N53125));
    INVX1 U40254 (.I(n45715), .ZN(N53126));
    INVX1 U40255 (.I(n21034), .ZN(N53127));
    NANDX1 U40256 (.A1(n18426), .A2(N6787), .ZN(N53128));
    INVX1 U40257 (.I(n31509), .ZN(N53129));
    NANDX1 U40258 (.A1(n50233), .A2(n27102), .ZN(N53130));
    NANDX1 U40259 (.A1(n46811), .A2(n50322), .ZN(N53131));
    NANDX1 U40260 (.A1(n23416), .A2(n49642), .ZN(N53132));
    INVX1 U40261 (.I(n44383), .ZN(N53133));
    INVX1 U40262 (.I(N9524), .ZN(N53134));
    NOR2X1 U40263 (.A1(N2225), .A2(n38748), .ZN(N53135));
    NOR2X1 U40264 (.A1(N10306), .A2(n29391), .ZN(N53136));
    NOR2X1 U40265 (.A1(n43890), .A2(n43575), .ZN(N53137));
    INVX1 U40266 (.I(N8044), .ZN(N53138));
    NOR2X1 U40267 (.A1(n39953), .A2(n21618), .ZN(N53139));
    NOR2X1 U40268 (.A1(n46739), .A2(n33823), .ZN(N53140));
    NOR2X1 U40269 (.A1(n35158), .A2(N2495), .ZN(N53141));
    NOR2X1 U40270 (.A1(n20483), .A2(n19333), .ZN(N53142));
    NANDX1 U40271 (.A1(n48376), .A2(n42749), .ZN(N53143));
    NANDX1 U40272 (.A1(n32335), .A2(n35543), .ZN(N53144));
    NOR2X1 U40273 (.A1(N11887), .A2(n15858), .ZN(N53145));
    NANDX1 U40274 (.A1(n50634), .A2(n29325), .ZN(N53146));
    NANDX1 U40275 (.A1(n50052), .A2(N3773), .ZN(N53147));
    NANDX1 U40276 (.A1(n42038), .A2(n22692), .ZN(N53148));
    NANDX1 U40277 (.A1(n24918), .A2(n32672), .ZN(N53149));
    INVX1 U40278 (.I(n47838), .ZN(N53150));
    INVX1 U40279 (.I(n36685), .ZN(N53151));
    NOR2X1 U40280 (.A1(N3036), .A2(N9208), .ZN(N53152));
    NOR2X1 U40281 (.A1(n45134), .A2(n28540), .ZN(N53153));
    INVX1 U40282 (.I(n41922), .ZN(N53154));
    NOR2X1 U40283 (.A1(n24492), .A2(n22668), .ZN(N53155));
    NOR2X1 U40284 (.A1(n22835), .A2(N4582), .ZN(N53156));
    NANDX1 U40285 (.A1(n45019), .A2(N3628), .ZN(N53157));
    INVX1 U40286 (.I(n25920), .ZN(N53158));
    INVX1 U40287 (.I(n14281), .ZN(N53159));
    INVX1 U40288 (.I(n35773), .ZN(N53160));
    INVX1 U40289 (.I(n31955), .ZN(N53161));
    INVX1 U40290 (.I(n39671), .ZN(N53162));
    INVX1 U40291 (.I(n26967), .ZN(N53163));
    NOR2X1 U40292 (.A1(N11558), .A2(n47673), .ZN(N53164));
    NANDX1 U40293 (.A1(n20765), .A2(n16761), .ZN(N53165));
    INVX1 U40294 (.I(n19333), .ZN(N53166));
    NOR2X1 U40295 (.A1(n46050), .A2(N9060), .ZN(N53167));
    NOR2X1 U40296 (.A1(n38745), .A2(N4358), .ZN(N53168));
    NOR2X1 U40297 (.A1(n43327), .A2(n37129), .ZN(N53169));
    INVX1 U40298 (.I(n16982), .ZN(N53170));
    NANDX1 U40299 (.A1(n21256), .A2(N10716), .ZN(N53171));
    NANDX1 U40300 (.A1(n20377), .A2(n46488), .ZN(N53172));
    NOR2X1 U40301 (.A1(n22360), .A2(n47233), .ZN(N53173));
    NANDX1 U40302 (.A1(n27205), .A2(n44228), .ZN(N53174));
    INVX1 U40303 (.I(N8790), .ZN(N53175));
    INVX1 U40304 (.I(n45156), .ZN(N53176));
    NOR2X1 U40305 (.A1(N5485), .A2(n19312), .ZN(N53177));
    NOR2X1 U40306 (.A1(n20008), .A2(n13773), .ZN(N53178));
    NANDX1 U40307 (.A1(n29051), .A2(N929), .ZN(N53179));
    NANDX1 U40308 (.A1(n30956), .A2(n14283), .ZN(N53180));
    NANDX1 U40309 (.A1(n26291), .A2(n31264), .ZN(N53181));
    INVX1 U40310 (.I(n47546), .ZN(N53182));
    INVX1 U40311 (.I(n45864), .ZN(N53183));
    INVX1 U40312 (.I(N6907), .ZN(N53184));
    NANDX1 U40313 (.A1(N8722), .A2(N2552), .ZN(N53185));
    NOR2X1 U40314 (.A1(N5954), .A2(n16807), .ZN(N53186));
    INVX1 U40315 (.I(n36359), .ZN(N53187));
    INVX1 U40316 (.I(n36796), .ZN(N53188));
    INVX1 U40317 (.I(n32630), .ZN(N53189));
    INVX1 U40318 (.I(N3267), .ZN(N53190));
    INVX1 U40319 (.I(n18291), .ZN(N53191));
    NOR2X1 U40320 (.A1(n21744), .A2(n40835), .ZN(N53192));
    NANDX1 U40321 (.A1(N1111), .A2(n25146), .ZN(N53193));
    NOR2X1 U40322 (.A1(n27401), .A2(N4821), .ZN(N53194));
    INVX1 U40323 (.I(n44975), .ZN(N53195));
    INVX1 U40324 (.I(n42954), .ZN(N53196));
    NANDX1 U40325 (.A1(n45351), .A2(n24585), .ZN(N53197));
    NANDX1 U40326 (.A1(n17930), .A2(N11624), .ZN(N53198));
    INVX1 U40327 (.I(n34736), .ZN(N53199));
    NOR2X1 U40328 (.A1(N809), .A2(N10293), .ZN(N53200));
    NOR2X1 U40329 (.A1(n36750), .A2(n12951), .ZN(N53201));
    NOR2X1 U40330 (.A1(N10044), .A2(n35616), .ZN(N53202));
    NOR2X1 U40331 (.A1(N11312), .A2(N5771), .ZN(n53203));
    NOR2X1 U40332 (.A1(n36555), .A2(n28497), .ZN(N53204));
    NANDX1 U40333 (.A1(n19726), .A2(N4309), .ZN(N53205));
    NANDX1 U40334 (.A1(n38432), .A2(n49283), .ZN(N53206));
    NOR2X1 U40335 (.A1(n29797), .A2(n50647), .ZN(N53207));
    NOR2X1 U40336 (.A1(N2793), .A2(N9144), .ZN(N53208));
    INVX1 U40337 (.I(n36033), .ZN(N53209));
    NOR2X1 U40338 (.A1(n25445), .A2(n39296), .ZN(N53210));
    NOR2X1 U40339 (.A1(N5765), .A2(n27767), .ZN(N53211));
    NANDX1 U40340 (.A1(n18715), .A2(n20755), .ZN(N53212));
    NANDX1 U40341 (.A1(n24358), .A2(n23678), .ZN(N53213));
    INVX1 U40342 (.I(n30128), .ZN(N53214));
    INVX1 U40343 (.I(n30733), .ZN(N53215));
    INVX1 U40344 (.I(n33161), .ZN(N53216));
    INVX1 U40345 (.I(n32961), .ZN(N53217));
    NOR2X1 U40346 (.A1(n37301), .A2(N683), .ZN(N53218));
    NOR2X1 U40347 (.A1(n37126), .A2(n51330), .ZN(N53219));
    NANDX1 U40348 (.A1(N9946), .A2(n30501), .ZN(N53220));
    NOR2X1 U40349 (.A1(n45978), .A2(N4095), .ZN(N53221));
    NANDX1 U40350 (.A1(n33686), .A2(n21729), .ZN(N53222));
    INVX1 U40351 (.I(n31480), .ZN(N53223));
    INVX1 U40352 (.I(n31013), .ZN(N53224));
    NANDX1 U40353 (.A1(n37362), .A2(N3783), .ZN(N53225));
    NOR2X1 U40354 (.A1(N9924), .A2(n33910), .ZN(N53226));
    INVX1 U40355 (.I(N10685), .ZN(N53227));
    NOR2X1 U40356 (.A1(n13385), .A2(n31170), .ZN(N53228));
    NOR2X1 U40357 (.A1(N8736), .A2(n38499), .ZN(N53229));
    NANDX1 U40358 (.A1(n34692), .A2(n24036), .ZN(N53230));
    NANDX1 U40359 (.A1(n33429), .A2(N4009), .ZN(N53231));
    NANDX1 U40360 (.A1(n22874), .A2(n20015), .ZN(n53232));
    INVX1 U40361 (.I(n29408), .ZN(N53233));
    NOR2X1 U40362 (.A1(N10764), .A2(n41706), .ZN(N53234));
    INVX1 U40363 (.I(n35287), .ZN(N53235));
    INVX1 U40364 (.I(n25880), .ZN(N53236));
    NOR2X1 U40365 (.A1(n24912), .A2(n41847), .ZN(N53237));
    INVX1 U40366 (.I(n28850), .ZN(N53238));
    NOR2X1 U40367 (.A1(n33312), .A2(N9851), .ZN(N53239));
    NOR2X1 U40368 (.A1(n12893), .A2(n45428), .ZN(N53240));
    NOR2X1 U40369 (.A1(n21419), .A2(n30099), .ZN(N53241));
    NANDX1 U40370 (.A1(n45454), .A2(n36128), .ZN(N53242));
    INVX1 U40371 (.I(n19491), .ZN(N53243));
    NOR2X1 U40372 (.A1(n45268), .A2(n39505), .ZN(N53244));
    INVX1 U40373 (.I(n44703), .ZN(N53245));
    INVX1 U40374 (.I(N12511), .ZN(N53246));
    NANDX1 U40375 (.A1(n15262), .A2(n17825), .ZN(N53247));
    NOR2X1 U40376 (.A1(N11169), .A2(N8912), .ZN(N53248));
    NOR2X1 U40377 (.A1(N1427), .A2(n31539), .ZN(N53249));
    NANDX1 U40378 (.A1(n23498), .A2(n13262), .ZN(N53250));
    NOR2X1 U40379 (.A1(n50597), .A2(n47771), .ZN(N53251));
    INVX1 U40380 (.I(n34843), .ZN(N53252));
    NOR2X1 U40381 (.A1(N1993), .A2(N2192), .ZN(N53253));
    NANDX1 U40382 (.A1(n38120), .A2(n24586), .ZN(N53254));
    INVX1 U40383 (.I(n29216), .ZN(N53255));
    NANDX1 U40384 (.A1(N10517), .A2(N9347), .ZN(N53256));
    INVX1 U40385 (.I(n22160), .ZN(N53257));
    NOR2X1 U40386 (.A1(n16226), .A2(N7449), .ZN(N53258));
    INVX1 U40387 (.I(n42202), .ZN(N53259));
    NANDX1 U40388 (.A1(n18621), .A2(N11530), .ZN(N53260));
    INVX1 U40389 (.I(n20187), .ZN(N53261));
    NANDX1 U40390 (.A1(n13569), .A2(n33449), .ZN(N53262));
    NANDX1 U40391 (.A1(N12577), .A2(n51247), .ZN(N53263));
    NOR2X1 U40392 (.A1(n47419), .A2(n17259), .ZN(N53264));
    INVX1 U40393 (.I(n19638), .ZN(N53265));
    NANDX1 U40394 (.A1(n51356), .A2(n44223), .ZN(N53266));
    NOR2X1 U40395 (.A1(n28984), .A2(n32515), .ZN(N53267));
    INVX1 U40396 (.I(N8358), .ZN(N53268));
    INVX1 U40397 (.I(n45672), .ZN(N53269));
    NOR2X1 U40398 (.A1(N174), .A2(N1532), .ZN(N53270));
    INVX1 U40399 (.I(N12404), .ZN(N53271));
    INVX1 U40400 (.I(n20215), .ZN(N53272));
    NOR2X1 U40401 (.A1(N10220), .A2(n40402), .ZN(N53273));
    NANDX1 U40402 (.A1(n45404), .A2(n43878), .ZN(N53274));
    INVX1 U40403 (.I(n28008), .ZN(N53275));
    NOR2X1 U40404 (.A1(n24289), .A2(n23838), .ZN(N53276));
    NOR2X1 U40405 (.A1(n37525), .A2(n43475), .ZN(N53277));
    NANDX1 U40406 (.A1(N7320), .A2(N6138), .ZN(N53278));
    INVX1 U40407 (.I(n36303), .ZN(N53279));
    NOR2X1 U40408 (.A1(n44468), .A2(n14689), .ZN(N53280));
    NANDX1 U40409 (.A1(N8579), .A2(n36547), .ZN(N53281));
    NANDX1 U40410 (.A1(N10111), .A2(n16525), .ZN(N53282));
    NOR2X1 U40411 (.A1(N287), .A2(N6768), .ZN(N53283));
    NOR2X1 U40412 (.A1(n32122), .A2(n47169), .ZN(N53284));
    NANDX1 U40413 (.A1(n25937), .A2(n39458), .ZN(N53285));
    NANDX1 U40414 (.A1(N2356), .A2(N1433), .ZN(N53286));
    NANDX1 U40415 (.A1(n47809), .A2(n32254), .ZN(N53287));
    NOR2X1 U40416 (.A1(N9723), .A2(N1884), .ZN(N53288));
    NOR2X1 U40417 (.A1(n15860), .A2(n44455), .ZN(N53289));
    NOR2X1 U40418 (.A1(n24540), .A2(N7362), .ZN(N53290));
    NOR2X1 U40419 (.A1(n17168), .A2(n15940), .ZN(N53291));
    INVX1 U40420 (.I(N9969), .ZN(N53292));
    NANDX1 U40421 (.A1(n39210), .A2(n36790), .ZN(N53293));
    NOR2X1 U40422 (.A1(n45977), .A2(N5983), .ZN(N53294));
    NOR2X1 U40423 (.A1(n41557), .A2(n30431), .ZN(N53295));
    NANDX1 U40424 (.A1(n51042), .A2(n37951), .ZN(N53296));
    NANDX1 U40425 (.A1(n22502), .A2(n48144), .ZN(N53297));
    NOR2X1 U40426 (.A1(N3167), .A2(n35916), .ZN(N53298));
    NOR2X1 U40427 (.A1(n26667), .A2(N9392), .ZN(N53299));
    INVX1 U40428 (.I(n19533), .ZN(N53300));
    NANDX1 U40429 (.A1(n13201), .A2(n48510), .ZN(N53301));
    NANDX1 U40430 (.A1(n30368), .A2(n34477), .ZN(N53302));
    NOR2X1 U40431 (.A1(n40337), .A2(n30555), .ZN(N53303));
    NANDX1 U40432 (.A1(n47154), .A2(n26918), .ZN(N53304));
    INVX1 U40433 (.I(N1548), .ZN(N53305));
    NOR2X1 U40434 (.A1(n21587), .A2(n31978), .ZN(N53306));
    INVX1 U40435 (.I(n21040), .ZN(N53307));
    INVX1 U40436 (.I(n46711), .ZN(N53308));
    NOR2X1 U40437 (.A1(n36511), .A2(n39762), .ZN(N53309));
    NANDX1 U40438 (.A1(n42455), .A2(n42536), .ZN(N53310));
    INVX1 U40439 (.I(N258), .ZN(N53311));
    INVX1 U40440 (.I(N2989), .ZN(N53312));
    NANDX1 U40441 (.A1(n44398), .A2(n51498), .ZN(N53313));
    INVX1 U40442 (.I(n44794), .ZN(N53314));
    INVX1 U40443 (.I(n44374), .ZN(N53315));
    NANDX1 U40444 (.A1(n34969), .A2(N8400), .ZN(N53316));
    NANDX1 U40445 (.A1(n31914), .A2(n18402), .ZN(N53317));
    INVX1 U40446 (.I(N5756), .ZN(N53318));
    INVX1 U40447 (.I(n32659), .ZN(N53319));
    INVX1 U40448 (.I(n31055), .ZN(N53320));
    NANDX1 U40449 (.A1(n42401), .A2(n44623), .ZN(N53321));
    INVX1 U40450 (.I(n30574), .ZN(N53322));
    NANDX1 U40451 (.A1(n18431), .A2(n43138), .ZN(N53323));
    INVX1 U40452 (.I(n40304), .ZN(n53324));
    INVX1 U40453 (.I(n17830), .ZN(N53325));
    INVX1 U40454 (.I(n37172), .ZN(N53326));
    INVX1 U40455 (.I(n37784), .ZN(N53327));
    NANDX1 U40456 (.A1(n22154), .A2(n30569), .ZN(N53328));
    INVX1 U40457 (.I(N5534), .ZN(N53329));
    NANDX1 U40458 (.A1(n33080), .A2(N7475), .ZN(N53330));
    NANDX1 U40459 (.A1(N3789), .A2(n13231), .ZN(N53331));
    NOR2X1 U40460 (.A1(n36447), .A2(N8921), .ZN(N53332));
    INVX1 U40461 (.I(n27501), .ZN(N53333));
    NOR2X1 U40462 (.A1(N1556), .A2(n25093), .ZN(N53334));
    NOR2X1 U40463 (.A1(N2968), .A2(n43523), .ZN(N53335));
    INVX1 U40464 (.I(n17809), .ZN(N53336));
    NOR2X1 U40465 (.A1(n36245), .A2(n35639), .ZN(N53337));
    INVX1 U40466 (.I(n21829), .ZN(N53338));
    NOR2X1 U40467 (.A1(n39836), .A2(n22233), .ZN(N53339));
    INVX1 U40468 (.I(n40432), .ZN(N53340));
    NANDX1 U40469 (.A1(n21120), .A2(n49427), .ZN(N53341));
    INVX1 U40470 (.I(n28594), .ZN(N53342));
    INVX1 U40471 (.I(n33103), .ZN(N53343));
    NANDX1 U40472 (.A1(n24318), .A2(n39577), .ZN(N53344));
    NOR2X1 U40473 (.A1(n32839), .A2(n37105), .ZN(N53345));
    NANDX1 U40474 (.A1(n34394), .A2(N10609), .ZN(N53346));
    NOR2X1 U40475 (.A1(N7390), .A2(N2543), .ZN(N53347));
    INVX1 U40476 (.I(n25198), .ZN(N53348));
    NOR2X1 U40477 (.A1(n18993), .A2(N9248), .ZN(N53349));
    NOR2X1 U40478 (.A1(n40821), .A2(N2681), .ZN(N53350));
    NOR2X1 U40479 (.A1(n33081), .A2(n48239), .ZN(N53351));
    NOR2X1 U40480 (.A1(n29315), .A2(n39386), .ZN(n53352));
    NOR2X1 U40481 (.A1(N7041), .A2(n38008), .ZN(N53353));
    NOR2X1 U40482 (.A1(N10171), .A2(n49859), .ZN(N53354));
    INVX1 U40483 (.I(n19775), .ZN(N53355));
    NOR2X1 U40484 (.A1(n17497), .A2(N5292), .ZN(N53356));
    NANDX1 U40485 (.A1(n21919), .A2(n15900), .ZN(N53357));
    NANDX1 U40486 (.A1(n29308), .A2(n40059), .ZN(N53358));
    NOR2X1 U40487 (.A1(N2917), .A2(n14895), .ZN(N53359));
    NANDX1 U40488 (.A1(n33781), .A2(n43371), .ZN(N53360));
    NANDX1 U40489 (.A1(n36461), .A2(N8507), .ZN(N53361));
    NANDX1 U40490 (.A1(N3140), .A2(n14075), .ZN(n53362));
    INVX1 U40491 (.I(n42525), .ZN(N53363));
    INVX1 U40492 (.I(n44134), .ZN(N53364));
    INVX1 U40493 (.I(n51025), .ZN(n53365));
    NANDX1 U40494 (.A1(n48831), .A2(n35683), .ZN(N53366));
    NOR2X1 U40495 (.A1(N7929), .A2(N1592), .ZN(N53367));
    NANDX1 U40496 (.A1(n39118), .A2(n45126), .ZN(N53368));
    NOR2X1 U40497 (.A1(N9585), .A2(n22845), .ZN(N53369));
    NANDX1 U40498 (.A1(n14387), .A2(n47377), .ZN(N53370));
    NANDX1 U40499 (.A1(n38181), .A2(n29569), .ZN(N53371));
    INVX1 U40500 (.I(n42851), .ZN(N53372));
    INVX1 U40501 (.I(N9006), .ZN(N53373));
    NOR2X1 U40502 (.A1(N9225), .A2(n23080), .ZN(N53374));
    NOR2X1 U40503 (.A1(n21777), .A2(n32204), .ZN(N53375));
    NOR2X1 U40504 (.A1(n20749), .A2(n31640), .ZN(N53376));
    INVX1 U40505 (.I(n39607), .ZN(N53377));
    INVX1 U40506 (.I(n23912), .ZN(N53378));
    NOR2X1 U40507 (.A1(n38942), .A2(n21720), .ZN(N53379));
    NOR2X1 U40508 (.A1(n32479), .A2(n27072), .ZN(N53380));
    NANDX1 U40509 (.A1(n25351), .A2(n20894), .ZN(N53381));
    INVX1 U40510 (.I(n21139), .ZN(N53382));
    NOR2X1 U40511 (.A1(n37270), .A2(n20736), .ZN(N53383));
    INVX1 U40512 (.I(n28532), .ZN(N53384));
    INVX1 U40513 (.I(n39114), .ZN(N53385));
    NANDX1 U40514 (.A1(n36045), .A2(n32221), .ZN(N53386));
    NANDX1 U40515 (.A1(N6233), .A2(n34452), .ZN(N53387));
    NANDX1 U40516 (.A1(n26981), .A2(n36119), .ZN(N53388));
    NOR2X1 U40517 (.A1(n14999), .A2(n21881), .ZN(N53389));
    NANDX1 U40518 (.A1(N10945), .A2(N9234), .ZN(N53390));
    NANDX1 U40519 (.A1(n46009), .A2(N11740), .ZN(N53391));
    NANDX1 U40520 (.A1(N9096), .A2(N7118), .ZN(n53392));
    INVX1 U40521 (.I(N8186), .ZN(N53393));
    NOR2X1 U40522 (.A1(n48987), .A2(n45455), .ZN(N53394));
    NOR2X1 U40523 (.A1(n27507), .A2(n22399), .ZN(N53395));
    NOR2X1 U40524 (.A1(n36648), .A2(n49971), .ZN(N53396));
    NANDX1 U40525 (.A1(n38896), .A2(n18856), .ZN(N53397));
    NOR2X1 U40526 (.A1(n21759), .A2(n46392), .ZN(N53398));
    NANDX1 U40527 (.A1(N6290), .A2(N2146), .ZN(N53399));
    INVX1 U40528 (.I(n49786), .ZN(N53400));
    NANDX1 U40529 (.A1(N7892), .A2(n29048), .ZN(N53401));
    INVX1 U40530 (.I(n23928), .ZN(N53402));
    NANDX1 U40531 (.A1(N3294), .A2(N3051), .ZN(N53403));
    INVX1 U40532 (.I(n22671), .ZN(N53404));
    INVX1 U40533 (.I(n46189), .ZN(N53405));
    NANDX1 U40534 (.A1(N5103), .A2(n13620), .ZN(N53406));
    NOR2X1 U40535 (.A1(n49117), .A2(N7871), .ZN(N53407));
    NOR2X1 U40536 (.A1(n47499), .A2(N8194), .ZN(N53408));
    NANDX1 U40537 (.A1(n14766), .A2(n44721), .ZN(N53409));
    NANDX1 U40538 (.A1(N9570), .A2(n26669), .ZN(N53410));
    INVX1 U40539 (.I(N11715), .ZN(N53411));
    NOR2X1 U40540 (.A1(n51092), .A2(n45112), .ZN(N53412));
    NANDX1 U40541 (.A1(n28551), .A2(n49922), .ZN(N53413));
    INVX1 U40542 (.I(n39365), .ZN(N53414));
    NANDX1 U40543 (.A1(n50128), .A2(N5709), .ZN(N53415));
    INVX1 U40544 (.I(N9776), .ZN(N53416));
    NOR2X1 U40545 (.A1(n36009), .A2(n36494), .ZN(N53417));
    NOR2X1 U40546 (.A1(n23640), .A2(n34022), .ZN(N53418));
    NANDX1 U40547 (.A1(n17947), .A2(n29932), .ZN(N53419));
    NANDX1 U40548 (.A1(n51149), .A2(n44697), .ZN(N53420));
    NOR2X1 U40549 (.A1(n46165), .A2(n24294), .ZN(N53421));
    INVX1 U40550 (.I(n47471), .ZN(N53422));
    NOR2X1 U40551 (.A1(n35079), .A2(n46974), .ZN(N53423));
    INVX1 U40552 (.I(N6641), .ZN(N53424));
    NOR2X1 U40553 (.A1(n19509), .A2(n32102), .ZN(N53425));
    INVX1 U40554 (.I(N12779), .ZN(N53426));
    INVX1 U40555 (.I(N9065), .ZN(N53427));
    NANDX1 U40556 (.A1(N10445), .A2(n30989), .ZN(N53428));
    NANDX1 U40557 (.A1(n46938), .A2(n14945), .ZN(N53429));
    NOR2X1 U40558 (.A1(n50987), .A2(n50002), .ZN(N53430));
    NOR2X1 U40559 (.A1(n29330), .A2(n20049), .ZN(N53431));
    NANDX1 U40560 (.A1(n44054), .A2(n26460), .ZN(N53432));
    NOR2X1 U40561 (.A1(n14059), .A2(n29815), .ZN(N53433));
    NANDX1 U40562 (.A1(N2970), .A2(n43796), .ZN(N53434));
    NOR2X1 U40563 (.A1(n48310), .A2(n41275), .ZN(N53435));
    NANDX1 U40564 (.A1(N11892), .A2(n25119), .ZN(N53436));
    NOR2X1 U40565 (.A1(n25361), .A2(N10543), .ZN(N53437));
    NANDX1 U40566 (.A1(n16589), .A2(n31423), .ZN(N53438));
    NANDX1 U40567 (.A1(n31774), .A2(n32043), .ZN(N53439));
    INVX1 U40568 (.I(N2296), .ZN(N53440));
    INVX1 U40569 (.I(n53027), .ZN(N53441));
    INVX1 U40570 (.I(n18253), .ZN(N53442));
    INVX1 U40571 (.I(n44138), .ZN(N53443));
    NOR2X1 U40572 (.A1(n34551), .A2(N7261), .ZN(N53444));
    NANDX1 U40573 (.A1(N12798), .A2(n53076), .ZN(N53445));
    NOR2X1 U40574 (.A1(N3161), .A2(n25921), .ZN(N53446));
    NANDX1 U40575 (.A1(n46300), .A2(n27503), .ZN(N53447));
    INVX1 U40576 (.I(n17986), .ZN(N53448));
    NOR2X1 U40577 (.A1(n49316), .A2(n28528), .ZN(N53449));
    NOR2X1 U40578 (.A1(N12472), .A2(N6518), .ZN(N53450));
    INVX1 U40579 (.I(n44245), .ZN(N53451));
    INVX1 U40580 (.I(N2686), .ZN(N53452));
    NANDX1 U40581 (.A1(n13177), .A2(N4144), .ZN(n53453));
    NANDX1 U40582 (.A1(n31429), .A2(n22106), .ZN(N53454));
    NANDX1 U40583 (.A1(n27860), .A2(N5088), .ZN(N53455));
    INVX1 U40584 (.I(n36485), .ZN(N53456));
    INVX1 U40585 (.I(n14753), .ZN(N53457));
    NANDX1 U40586 (.A1(n22910), .A2(n42537), .ZN(N53458));
    INVX1 U40587 (.I(n15777), .ZN(N53459));
    NANDX1 U40588 (.A1(n28803), .A2(n33762), .ZN(N53460));
    NANDX1 U40589 (.A1(n26550), .A2(N8857), .ZN(N53461));
    NOR2X1 U40590 (.A1(n40187), .A2(n30701), .ZN(N53462));
    NOR2X1 U40591 (.A1(n32523), .A2(n48218), .ZN(N53463));
    NANDX1 U40592 (.A1(n45651), .A2(n49010), .ZN(N53464));
    NOR2X1 U40593 (.A1(N5299), .A2(n39412), .ZN(N53465));
    INVX1 U40594 (.I(N6811), .ZN(N53466));
    INVX1 U40595 (.I(n48403), .ZN(N53467));
    NOR2X1 U40596 (.A1(n22533), .A2(n34444), .ZN(N53468));
    NANDX1 U40597 (.A1(N12163), .A2(n29532), .ZN(N53469));
    NANDX1 U40598 (.A1(n15775), .A2(n14649), .ZN(N53470));
    NOR2X1 U40599 (.A1(n20865), .A2(n49775), .ZN(N53471));
    NOR2X1 U40600 (.A1(n14985), .A2(n41370), .ZN(N53472));
    NOR2X1 U40601 (.A1(N1710), .A2(n18609), .ZN(N53473));
    NANDX1 U40602 (.A1(n25494), .A2(n13365), .ZN(N53474));
    INVX1 U40603 (.I(N8944), .ZN(N53475));
    INVX1 U40604 (.I(n40451), .ZN(N53476));
    NOR2X1 U40605 (.A1(n39585), .A2(n21110), .ZN(N53477));
    NOR2X1 U40606 (.A1(N6203), .A2(N7313), .ZN(N53478));
    NANDX1 U40607 (.A1(n19996), .A2(n41756), .ZN(N53479));
    NOR2X1 U40608 (.A1(n23419), .A2(N9087), .ZN(N53480));
    NANDX1 U40609 (.A1(n39193), .A2(n14997), .ZN(N53481));
    NANDX1 U40610 (.A1(N6596), .A2(N2571), .ZN(N53482));
    NANDX1 U40611 (.A1(N12841), .A2(n43941), .ZN(N53483));
    INVX1 U40612 (.I(N5811), .ZN(N53484));
    INVX1 U40613 (.I(N336), .ZN(N53485));
    INVX1 U40614 (.I(n13714), .ZN(N53486));
    NOR2X1 U40615 (.A1(n31509), .A2(n13887), .ZN(N53487));
    NOR2X1 U40616 (.A1(n37012), .A2(N11), .ZN(N53488));
    NANDX1 U40617 (.A1(n40586), .A2(n50935), .ZN(N53489));
    NANDX1 U40618 (.A1(n49134), .A2(n17469), .ZN(N53490));
    NOR2X1 U40619 (.A1(n32520), .A2(n40887), .ZN(N53491));
    INVX1 U40620 (.I(N8461), .ZN(N53492));
    NOR2X1 U40621 (.A1(N9019), .A2(n30397), .ZN(N53493));
    NOR2X1 U40622 (.A1(N11589), .A2(n18077), .ZN(N53494));
    NOR2X1 U40623 (.A1(N2068), .A2(N294), .ZN(N53495));
    INVX1 U40624 (.I(N2417), .ZN(N53496));
    INVX1 U40625 (.I(N3489), .ZN(N53497));
    NOR2X1 U40626 (.A1(n52799), .A2(n34997), .ZN(N53498));
    INVX1 U40627 (.I(n29758), .ZN(N53499));
    NOR2X1 U40628 (.A1(N12548), .A2(n27826), .ZN(N53500));
    NANDX1 U40629 (.A1(N10021), .A2(n24467), .ZN(N53501));
    NOR2X1 U40630 (.A1(n18750), .A2(N9402), .ZN(N53502));
    NOR2X1 U40631 (.A1(n50897), .A2(n48146), .ZN(N53503));
    INVX1 U40632 (.I(n15314), .ZN(N53504));
    INVX1 U40633 (.I(n46502), .ZN(N53505));
    NANDX1 U40634 (.A1(n51275), .A2(N2378), .ZN(N53506));
    NANDX1 U40635 (.A1(n44603), .A2(N2672), .ZN(N53507));
    INVX1 U40636 (.I(n38280), .ZN(N53508));
    NANDX1 U40637 (.A1(n26556), .A2(n45670), .ZN(N53509));
    NANDX1 U40638 (.A1(n52813), .A2(N4747), .ZN(N53510));
    NANDX1 U40639 (.A1(N420), .A2(n17294), .ZN(N53511));
    INVX1 U40640 (.I(n42073), .ZN(N53512));
    NANDX1 U40641 (.A1(N5008), .A2(n17199), .ZN(N53513));
    NANDX1 U40642 (.A1(N5671), .A2(n16105), .ZN(N53514));
    INVX1 U40643 (.I(n45077), .ZN(N53515));
    NANDX1 U40644 (.A1(n41335), .A2(n40041), .ZN(N53516));
    INVX1 U40645 (.I(N10183), .ZN(N53517));
    NANDX1 U40646 (.A1(n18889), .A2(n52326), .ZN(N53518));
    NANDX1 U40647 (.A1(N12821), .A2(n21932), .ZN(N53519));
    NANDX1 U40648 (.A1(n52104), .A2(n48487), .ZN(N53520));
    NOR2X1 U40649 (.A1(n37263), .A2(n39099), .ZN(N53521));
    NOR2X1 U40650 (.A1(n43441), .A2(n39518), .ZN(N53522));
    NOR2X1 U40651 (.A1(n23982), .A2(n19391), .ZN(N53523));
    INVX1 U40652 (.I(n20251), .ZN(N53524));
    INVX1 U40653 (.I(N4283), .ZN(N53525));
    INVX1 U40654 (.I(n43954), .ZN(N53526));
    INVX1 U40655 (.I(N8797), .ZN(N53527));
    NOR2X1 U40656 (.A1(N9439), .A2(n40098), .ZN(N53528));
    INVX1 U40657 (.I(N10882), .ZN(N53529));
    NANDX1 U40658 (.A1(n49361), .A2(N9746), .ZN(N53530));
    NANDX1 U40659 (.A1(N8720), .A2(n22939), .ZN(N53531));
    NOR2X1 U40660 (.A1(N7362), .A2(n17964), .ZN(N53532));
    NOR2X1 U40661 (.A1(n35886), .A2(n48324), .ZN(N53533));
    INVX1 U40662 (.I(n17126), .ZN(N53534));
    INVX1 U40663 (.I(n24758), .ZN(N53535));
    NANDX1 U40664 (.A1(n36292), .A2(n45177), .ZN(N53536));
    INVX1 U40665 (.I(N10680), .ZN(N53537));
    INVX1 U40666 (.I(N7599), .ZN(N53538));
    NANDX1 U40667 (.A1(N8824), .A2(N7657), .ZN(N53539));
    NANDX1 U40668 (.A1(N9523), .A2(n39015), .ZN(N53540));
    INVX1 U40669 (.I(N11665), .ZN(N53541));
    INVX1 U40670 (.I(n32767), .ZN(N53542));
    NOR2X1 U40671 (.A1(n19833), .A2(n41487), .ZN(N53543));
    INVX1 U40672 (.I(n43435), .ZN(N53544));
    NANDX1 U40673 (.A1(n44834), .A2(N10858), .ZN(N53545));
    NANDX1 U40674 (.A1(n39696), .A2(n25032), .ZN(N53546));
    INVX1 U40675 (.I(N11875), .ZN(N53547));
    INVX1 U40676 (.I(n18565), .ZN(N53548));
    INVX1 U40677 (.I(n24026), .ZN(N53549));
    INVX1 U40678 (.I(n50107), .ZN(N53550));
    INVX1 U40679 (.I(N7842), .ZN(N53551));
    INVX1 U40680 (.I(N11369), .ZN(N53552));
    NOR2X1 U40681 (.A1(n40195), .A2(N12152), .ZN(N53553));
    NOR2X1 U40682 (.A1(n23601), .A2(n23816), .ZN(N53554));
    NOR2X1 U40683 (.A1(N2907), .A2(n36486), .ZN(N53555));
    NANDX1 U40684 (.A1(n35654), .A2(n18634), .ZN(N53556));
    NOR2X1 U40685 (.A1(n22301), .A2(N10006), .ZN(N53557));
    INVX1 U40686 (.I(n36095), .ZN(N53558));
    NOR2X1 U40687 (.A1(n21832), .A2(n13552), .ZN(N53559));
    INVX1 U40688 (.I(N682), .ZN(N53560));
    INVX1 U40689 (.I(n30063), .ZN(N53561));
    NOR2X1 U40690 (.A1(n23620), .A2(n26709), .ZN(N53562));
    NOR2X1 U40691 (.A1(n31461), .A2(N7048), .ZN(N53563));
    NANDX1 U40692 (.A1(n38219), .A2(n38503), .ZN(N53564));
    NOR2X1 U40693 (.A1(n39269), .A2(N8643), .ZN(N53565));
    NANDX1 U40694 (.A1(n24146), .A2(N11549), .ZN(N53566));
    NOR2X1 U40695 (.A1(n28854), .A2(n38463), .ZN(N53567));
    NANDX1 U40696 (.A1(n23536), .A2(n52024), .ZN(N53568));
    INVX1 U40697 (.I(n20336), .ZN(N53569));
    INVX1 U40698 (.I(n30054), .ZN(N53570));
    INVX1 U40699 (.I(n39470), .ZN(N53571));
    NOR2X1 U40700 (.A1(n25370), .A2(N646), .ZN(N53572));
    NANDX1 U40701 (.A1(n41338), .A2(n15526), .ZN(N53573));
    NANDX1 U40702 (.A1(N6389), .A2(n46986), .ZN(N53574));
    NANDX1 U40703 (.A1(n18792), .A2(n31743), .ZN(N53575));
    NOR2X1 U40704 (.A1(n52084), .A2(N8812), .ZN(N53576));
    NOR2X1 U40705 (.A1(n38253), .A2(n24218), .ZN(N53577));
    INVX1 U40706 (.I(n16185), .ZN(N53578));
    NANDX1 U40707 (.A1(n48522), .A2(n48733), .ZN(N53579));
    NOR2X1 U40708 (.A1(n47085), .A2(n37825), .ZN(N53580));
    NANDX1 U40709 (.A1(n19541), .A2(N5678), .ZN(N53581));
    INVX1 U40710 (.I(n50271), .ZN(N53582));
    INVX1 U40711 (.I(n22599), .ZN(N53583));
    NOR2X1 U40712 (.A1(n14917), .A2(N10475), .ZN(N53584));
    NOR2X1 U40713 (.A1(n21437), .A2(N8125), .ZN(N53585));
    INVX1 U40714 (.I(n35004), .ZN(N53586));
    NOR2X1 U40715 (.A1(N12031), .A2(n24874), .ZN(N53587));
    NOR2X1 U40716 (.A1(n20842), .A2(n23385), .ZN(N53588));
    NANDX1 U40717 (.A1(n36320), .A2(n33445), .ZN(N53589));
    NOR2X1 U40718 (.A1(n27191), .A2(n19766), .ZN(N53590));
    INVX1 U40719 (.I(n32857), .ZN(N53591));
    NOR2X1 U40720 (.A1(n24652), .A2(N5398), .ZN(N53592));
    NANDX1 U40721 (.A1(n30329), .A2(N2627), .ZN(N53593));
    NANDX1 U40722 (.A1(n47956), .A2(n16486), .ZN(N53594));
    NANDX1 U40723 (.A1(N672), .A2(n18222), .ZN(N53595));
    NANDX1 U40724 (.A1(n22109), .A2(n17607), .ZN(N53596));
    NANDX1 U40725 (.A1(n48373), .A2(n35783), .ZN(N53597));
    INVX1 U40726 (.I(N11046), .ZN(N53598));
    NANDX1 U40727 (.A1(N9640), .A2(n34431), .ZN(N53599));
    INVX1 U40728 (.I(n45959), .ZN(n53600));
    NOR2X1 U40729 (.A1(n36988), .A2(n19688), .ZN(N53601));
    NANDX1 U40730 (.A1(n32555), .A2(n52545), .ZN(N53602));
    NOR2X1 U40731 (.A1(n48467), .A2(n49203), .ZN(N53603));
    INVX1 U40732 (.I(n25335), .ZN(N53604));
    NANDX1 U40733 (.A1(n40323), .A2(N11090), .ZN(N53605));
    NANDX1 U40734 (.A1(n32561), .A2(N11761), .ZN(N53606));
    NOR2X1 U40735 (.A1(n20301), .A2(n25130), .ZN(N53607));
    INVX1 U40736 (.I(N5807), .ZN(N53608));
    INVX1 U40737 (.I(n15523), .ZN(N53609));
    NOR2X1 U40738 (.A1(n22348), .A2(n50626), .ZN(N53610));
    NANDX1 U40739 (.A1(n48039), .A2(n33857), .ZN(N53611));
    NANDX1 U40740 (.A1(N252), .A2(N8644), .ZN(N53612));
    NOR2X1 U40741 (.A1(n16953), .A2(n41198), .ZN(N53613));
    NOR2X1 U40742 (.A1(n38303), .A2(n36204), .ZN(N53614));
    NOR2X1 U40743 (.A1(n12904), .A2(n52799), .ZN(N53615));
    INVX1 U40744 (.I(n44487), .ZN(N53616));
    NOR2X1 U40745 (.A1(n25499), .A2(n14847), .ZN(N53617));
    INVX1 U40746 (.I(n49833), .ZN(N53618));
    NANDX1 U40747 (.A1(n29839), .A2(n20835), .ZN(N53619));
    NOR2X1 U40748 (.A1(n32402), .A2(n36357), .ZN(N53620));
    INVX1 U40749 (.I(n46010), .ZN(N53621));
    NOR2X1 U40750 (.A1(n31060), .A2(n40588), .ZN(N53622));
    NOR2X1 U40751 (.A1(N10322), .A2(n32100), .ZN(N53623));
    INVX1 U40752 (.I(N9272), .ZN(N53624));
    NANDX1 U40753 (.A1(n46279), .A2(N7304), .ZN(N53625));
    INVX1 U40754 (.I(n20282), .ZN(N53626));
    INVX1 U40755 (.I(n29318), .ZN(N53627));
    NANDX1 U40756 (.A1(N11723), .A2(n20344), .ZN(N53628));
    INVX1 U40757 (.I(n37221), .ZN(N53629));
    NANDX1 U40758 (.A1(n26015), .A2(n24854), .ZN(N53630));
    INVX1 U40759 (.I(n47114), .ZN(n53631));
    NOR2X1 U40760 (.A1(n49089), .A2(n17315), .ZN(N53632));
    INVX1 U40761 (.I(n22445), .ZN(N53633));
    NOR2X1 U40762 (.A1(n53365), .A2(n44766), .ZN(N53634));
    NOR2X1 U40763 (.A1(N5080), .A2(N1626), .ZN(N53635));
    NOR2X1 U40764 (.A1(N10161), .A2(N10897), .ZN(N53636));
    NANDX1 U40765 (.A1(N2979), .A2(N9462), .ZN(N53637));
    NOR2X1 U40766 (.A1(n23260), .A2(n46522), .ZN(N53638));
    NOR2X1 U40767 (.A1(n34140), .A2(n49505), .ZN(N53639));
    INVX1 U40768 (.I(n46706), .ZN(N53640));
    INVX1 U40769 (.I(n46266), .ZN(N53641));
    NANDX1 U40770 (.A1(n49379), .A2(N941), .ZN(N53642));
    NOR2X1 U40771 (.A1(n41605), .A2(n50029), .ZN(N53643));
    INVX1 U40772 (.I(N7987), .ZN(N53644));
    NOR2X1 U40773 (.A1(n13871), .A2(n52612), .ZN(N53645));
    NOR2X1 U40774 (.A1(n46842), .A2(n48953), .ZN(N53646));
    INVX1 U40775 (.I(N4991), .ZN(N53647));
    INVX1 U40776 (.I(n50083), .ZN(N53648));
    INVX1 U40777 (.I(n53352), .ZN(N53649));
    NANDX1 U40778 (.A1(n18329), .A2(n23151), .ZN(N53650));
    NOR2X1 U40779 (.A1(N9061), .A2(N3829), .ZN(N53651));
    NOR2X1 U40780 (.A1(n20137), .A2(n50534), .ZN(N53652));
    INVX1 U40781 (.I(n12941), .ZN(N53653));
    INVX1 U40782 (.I(n51611), .ZN(N53654));
    INVX1 U40783 (.I(N3025), .ZN(N53655));
    NANDX1 U40784 (.A1(N1709), .A2(n15772), .ZN(N53656));
    NANDX1 U40785 (.A1(N11982), .A2(n29642), .ZN(N53657));
    INVX1 U40786 (.I(N4820), .ZN(N53658));
    NANDX1 U40787 (.A1(n16165), .A2(n44006), .ZN(N53659));
    INVX1 U40788 (.I(n13078), .ZN(N53660));
    NANDX1 U40789 (.A1(n13987), .A2(n12968), .ZN(N53661));
    INVX1 U40790 (.I(n23576), .ZN(N53662));
    NOR2X1 U40791 (.A1(n19634), .A2(n32636), .ZN(N53663));
    INVX1 U40792 (.I(n42063), .ZN(N53664));
    INVX1 U40793 (.I(n19541), .ZN(N53665));
    INVX1 U40794 (.I(N3512), .ZN(N53666));
    NOR2X1 U40795 (.A1(n42445), .A2(N8653), .ZN(N53667));
    NOR2X1 U40796 (.A1(n19999), .A2(N10362), .ZN(N53668));
    NANDX1 U40797 (.A1(n50261), .A2(n13604), .ZN(N53669));
    NOR2X1 U40798 (.A1(n17473), .A2(N9685), .ZN(N53670));
    NANDX1 U40799 (.A1(n24899), .A2(n44951), .ZN(N53671));
    NOR2X1 U40800 (.A1(n37976), .A2(n32116), .ZN(N53672));
    NANDX1 U40801 (.A1(n50943), .A2(n52607), .ZN(N53673));
    NANDX1 U40802 (.A1(n24861), .A2(n18779), .ZN(N53674));
    INVX1 U40803 (.I(N2606), .ZN(N53675));
    NOR2X1 U40804 (.A1(n28015), .A2(n22146), .ZN(N53676));
    NOR2X1 U40805 (.A1(n22787), .A2(n40539), .ZN(N53677));
    NOR2X1 U40806 (.A1(n31440), .A2(N8496), .ZN(N53678));
    NANDX1 U40807 (.A1(n33062), .A2(n45684), .ZN(N53679));
    NANDX1 U40808 (.A1(n37926), .A2(n50314), .ZN(N53680));
    NOR2X1 U40809 (.A1(n38871), .A2(n15765), .ZN(N53681));
    NOR2X1 U40810 (.A1(n30360), .A2(n45211), .ZN(N53682));
    NOR2X1 U40811 (.A1(N275), .A2(n35182), .ZN(N53683));
    NANDX1 U40812 (.A1(n52881), .A2(n39989), .ZN(N53684));
    INVX1 U40813 (.I(N9459), .ZN(N53685));
    INVX1 U40814 (.I(N12131), .ZN(N53686));
    INVX1 U40815 (.I(n34506), .ZN(N53687));
    NOR2X1 U40816 (.A1(n51035), .A2(n48554), .ZN(N53688));
    NANDX1 U40817 (.A1(n20754), .A2(n17793), .ZN(N53689));
    INVX1 U40818 (.I(N1732), .ZN(N53690));
    INVX1 U40819 (.I(n13333), .ZN(N53691));
    NOR2X1 U40820 (.A1(n26579), .A2(N10185), .ZN(N53692));
    NOR2X1 U40821 (.A1(N11989), .A2(n25949), .ZN(N53693));
    NANDX1 U40822 (.A1(n42348), .A2(n17698), .ZN(N53694));
    NOR2X1 U40823 (.A1(n42623), .A2(n44140), .ZN(N53695));
    NANDX1 U40824 (.A1(n42042), .A2(n21928), .ZN(N53696));
    NOR2X1 U40825 (.A1(n51501), .A2(n28419), .ZN(N53697));
    NOR2X1 U40826 (.A1(n50861), .A2(N725), .ZN(N53698));
    NOR2X1 U40827 (.A1(n48434), .A2(n49278), .ZN(N53699));
    NANDX1 U40828 (.A1(n15727), .A2(n13609), .ZN(N53700));
    NANDX1 U40829 (.A1(n17458), .A2(N2262), .ZN(N53701));
    INVX1 U40830 (.I(n41689), .ZN(N53702));
    NANDX1 U40831 (.A1(n44970), .A2(n52430), .ZN(N53703));
    NANDX1 U40832 (.A1(N8718), .A2(n21118), .ZN(N53704));
    INVX1 U40833 (.I(n17676), .ZN(N53705));
    NOR2X1 U40834 (.A1(n46120), .A2(N8354), .ZN(N53706));
    NANDX1 U40835 (.A1(n25961), .A2(n21542), .ZN(N53707));
    INVX1 U40836 (.I(n15261), .ZN(N53708));
    NOR2X1 U40837 (.A1(n16382), .A2(N12660), .ZN(N53709));
    INVX1 U40838 (.I(N4111), .ZN(N53710));
    NANDX1 U40839 (.A1(n37762), .A2(N4455), .ZN(N53711));
    NANDX1 U40840 (.A1(n51370), .A2(n25909), .ZN(N53712));
    NOR2X1 U40841 (.A1(n44892), .A2(N7233), .ZN(N53713));
    NANDX1 U40842 (.A1(N11531), .A2(n43464), .ZN(N53714));
    NOR2X1 U40843 (.A1(n43620), .A2(n52181), .ZN(N53715));
    INVX1 U40844 (.I(n47117), .ZN(N53716));
    NOR2X1 U40845 (.A1(n53362), .A2(n39775), .ZN(N53717));
    INVX1 U40846 (.I(n33089), .ZN(N53718));
    NANDX1 U40847 (.A1(n28813), .A2(n25077), .ZN(N53719));
    INVX1 U40848 (.I(n25312), .ZN(N53720));
    INVX1 U40849 (.I(n31455), .ZN(N53721));
    NANDX1 U40850 (.A1(n28091), .A2(n39087), .ZN(N53722));
    INVX1 U40851 (.I(n32545), .ZN(N53723));
    NOR2X1 U40852 (.A1(n40726), .A2(N4992), .ZN(N53724));
    NOR2X1 U40853 (.A1(n32156), .A2(N12225), .ZN(N53725));
    NANDX1 U40854 (.A1(n34947), .A2(N2227), .ZN(N53726));
    NANDX1 U40855 (.A1(n25105), .A2(n45668), .ZN(N53727));
    NOR2X1 U40856 (.A1(N10021), .A2(n53324), .ZN(N53728));
    NOR2X1 U40857 (.A1(n41056), .A2(N7134), .ZN(N53729));
    NOR2X1 U40858 (.A1(n44591), .A2(n35946), .ZN(N53730));
    NOR2X1 U40859 (.A1(n18664), .A2(n52518), .ZN(N53731));
    INVX1 U40860 (.I(n50118), .ZN(N53732));
    INVX1 U40861 (.I(n19369), .ZN(N53733));
    INVX1 U40862 (.I(n46930), .ZN(N53734));
    NANDX1 U40863 (.A1(N9771), .A2(n34194), .ZN(N53735));
    NOR2X1 U40864 (.A1(n24614), .A2(N4149), .ZN(N53736));
    NOR2X1 U40865 (.A1(n24805), .A2(n39095), .ZN(N53737));
    INVX1 U40866 (.I(n35528), .ZN(N53738));
    NOR2X1 U40867 (.A1(n46084), .A2(N6962), .ZN(N53739));
    INVX1 U40868 (.I(n37207), .ZN(N53740));
    NOR2X1 U40869 (.A1(n44337), .A2(n44340), .ZN(N53741));
    NOR2X1 U40870 (.A1(n35466), .A2(n26824), .ZN(N53742));
    NOR2X1 U40871 (.A1(N668), .A2(n25880), .ZN(N53743));
    NOR2X1 U40872 (.A1(n42046), .A2(n21253), .ZN(N53744));
    NOR2X1 U40873 (.A1(N6850), .A2(n14721), .ZN(N53745));
    NANDX1 U40874 (.A1(n16621), .A2(n40175), .ZN(N53746));
    INVX1 U40875 (.I(n32495), .ZN(N53747));
    NOR2X1 U40876 (.A1(n23977), .A2(N3838), .ZN(N53748));
    NOR2X1 U40877 (.A1(n24392), .A2(n30626), .ZN(N53749));
    NANDX1 U40878 (.A1(N8275), .A2(n28848), .ZN(N53750));
    NOR2X1 U40879 (.A1(n45482), .A2(n51866), .ZN(N53751));
    INVX1 U40880 (.I(n36360), .ZN(N53752));
    NOR2X1 U40881 (.A1(n52837), .A2(N984), .ZN(N53753));
    NANDX1 U40882 (.A1(n44765), .A2(n18124), .ZN(N53754));
    NANDX1 U40883 (.A1(n24611), .A2(n39377), .ZN(N53755));
    NANDX1 U40884 (.A1(n22721), .A2(N636), .ZN(N53756));
    NOR2X1 U40885 (.A1(n39341), .A2(n32072), .ZN(N53757));
    NANDX1 U40886 (.A1(N9636), .A2(n22933), .ZN(N53758));
    INVX1 U40887 (.I(N4734), .ZN(N53759));
    INVX1 U40888 (.I(N12355), .ZN(N53760));
    INVX1 U40889 (.I(N5166), .ZN(N53761));
    INVX1 U40890 (.I(N10746), .ZN(N53762));
    INVX1 U40891 (.I(N3911), .ZN(N53763));
    NANDX1 U40892 (.A1(n40295), .A2(n31531), .ZN(N53764));
    NANDX1 U40893 (.A1(n30932), .A2(n23775), .ZN(N53765));
    INVX1 U40894 (.I(n13496), .ZN(N53766));
    NANDX1 U40895 (.A1(N2032), .A2(n38106), .ZN(N53767));
    NANDX1 U40896 (.A1(n42289), .A2(n52088), .ZN(N53768));
    NOR2X1 U40897 (.A1(n51429), .A2(n29228), .ZN(N53769));
    NANDX1 U40898 (.A1(n32894), .A2(n38863), .ZN(N53770));
    INVX1 U40899 (.I(n29596), .ZN(N53771));
    INVX1 U40900 (.I(n47924), .ZN(N53772));
    NANDX1 U40901 (.A1(N8017), .A2(n44351), .ZN(N53773));
    NOR2X1 U40902 (.A1(N10023), .A2(n13813), .ZN(N53774));
    NANDX1 U40903 (.A1(N10434), .A2(n45368), .ZN(N53775));
    NOR2X1 U40904 (.A1(n19210), .A2(n22838), .ZN(N53776));
    NANDX1 U40905 (.A1(n13614), .A2(n36334), .ZN(N53777));
    INVX1 U40906 (.I(N6906), .ZN(N53778));
    NANDX1 U40907 (.A1(n49627), .A2(n49194), .ZN(N53779));
    INVX1 U40908 (.I(N7137), .ZN(N53780));
    NANDX1 U40909 (.A1(n40093), .A2(n50178), .ZN(N53781));
    NANDX1 U40910 (.A1(n16755), .A2(N491), .ZN(N53782));
    NANDX1 U40911 (.A1(n42873), .A2(n39676), .ZN(N53783));
    NANDX1 U40912 (.A1(n50889), .A2(n30565), .ZN(N53784));
    INVX1 U40913 (.I(N7451), .ZN(N53785));
    NANDX1 U40914 (.A1(N5649), .A2(n17884), .ZN(N53786));
    NANDX1 U40915 (.A1(n32729), .A2(n28354), .ZN(N53787));
    NOR2X1 U40916 (.A1(n21383), .A2(n33228), .ZN(N53788));
    INVX1 U40917 (.I(n51936), .ZN(N53789));
    NOR2X1 U40918 (.A1(n36753), .A2(n39362), .ZN(N53790));
    INVX1 U40919 (.I(n38879), .ZN(N53791));
    NOR2X1 U40920 (.A1(n20826), .A2(n16771), .ZN(N53792));
    INVX1 U40921 (.I(n29941), .ZN(N53793));
    NANDX1 U40922 (.A1(n34966), .A2(n15189), .ZN(N53794));
    NANDX1 U40923 (.A1(n21180), .A2(n33648), .ZN(N53795));
    NANDX1 U40924 (.A1(n51744), .A2(n43747), .ZN(N53796));
    NANDX1 U40925 (.A1(n33920), .A2(n40656), .ZN(N53797));
    INVX1 U40926 (.I(N8003), .ZN(N53798));
    INVX1 U40927 (.I(N3112), .ZN(n53799));
    INVX1 U40928 (.I(n32566), .ZN(N53800));
    NOR2X1 U40929 (.A1(n29437), .A2(n22301), .ZN(N53801));
    NOR2X1 U40930 (.A1(N3989), .A2(N8202), .ZN(N53802));
    INVX1 U40931 (.I(n42867), .ZN(N53803));
    INVX1 U40932 (.I(N8762), .ZN(N53804));
    NOR2X1 U40933 (.A1(n35713), .A2(n38702), .ZN(N53805));
    NANDX1 U40934 (.A1(N8479), .A2(n45152), .ZN(N53806));
    NOR2X1 U40935 (.A1(n20919), .A2(n16599), .ZN(N53807));
    INVX1 U40936 (.I(N10463), .ZN(N53808));
    NOR2X1 U40937 (.A1(N4919), .A2(n44382), .ZN(N53809));
    INVX1 U40938 (.I(n33137), .ZN(N53810));
    INVX1 U40939 (.I(N5261), .ZN(N53811));
    INVX1 U40940 (.I(N3845), .ZN(N53812));
    NOR2X1 U40941 (.A1(N1648), .A2(n24542), .ZN(N53813));
    NANDX1 U40942 (.A1(N7180), .A2(n28531), .ZN(N53814));
    NOR2X1 U40943 (.A1(n48577), .A2(N9197), .ZN(N53815));
    INVX1 U40944 (.I(n48599), .ZN(N53816));
    NANDX1 U40945 (.A1(n34339), .A2(n33840), .ZN(N53817));
    NOR2X1 U40946 (.A1(n34078), .A2(n16791), .ZN(N53818));
    NANDX1 U40947 (.A1(N1536), .A2(n33389), .ZN(N53819));
    NOR2X1 U40948 (.A1(N3259), .A2(n31534), .ZN(N53820));
    NOR2X1 U40949 (.A1(n47640), .A2(n16872), .ZN(N53821));
    NANDX1 U40950 (.A1(n37824), .A2(n13394), .ZN(N53822));
    NANDX1 U40951 (.A1(n32929), .A2(n42481), .ZN(N53823));
    NOR2X1 U40952 (.A1(N4010), .A2(n40407), .ZN(N53824));
    NOR2X1 U40953 (.A1(n23801), .A2(n46535), .ZN(N53825));
    INVX1 U40954 (.I(n32997), .ZN(N53826));
    NOR2X1 U40955 (.A1(n36082), .A2(n39630), .ZN(N53827));
    NANDX1 U40956 (.A1(N7721), .A2(n15024), .ZN(N53828));
    INVX1 U40957 (.I(n24511), .ZN(N53829));
    NANDX1 U40958 (.A1(n44173), .A2(N4438), .ZN(N53830));
    NANDX1 U40959 (.A1(n47431), .A2(n27232), .ZN(N53831));
    NANDX1 U40960 (.A1(n32870), .A2(n44104), .ZN(N53832));
    NOR2X1 U40961 (.A1(N8493), .A2(N4036), .ZN(N53833));
    NOR2X1 U40962 (.A1(n41422), .A2(n46516), .ZN(N53834));
    NOR2X1 U40963 (.A1(n36692), .A2(n24722), .ZN(N53835));
    NOR2X1 U40964 (.A1(n51753), .A2(n17795), .ZN(N53836));
    INVX1 U40965 (.I(n31288), .ZN(N53837));
    INVX1 U40966 (.I(n29962), .ZN(N53838));
    INVX1 U40967 (.I(n26793), .ZN(N53839));
    INVX1 U40968 (.I(n23741), .ZN(N53840));
    INVX1 U40969 (.I(n53453), .ZN(N53841));
    NOR2X1 U40970 (.A1(N6680), .A2(n49152), .ZN(N53842));
    INVX1 U40971 (.I(n45371), .ZN(N53843));
    NANDX1 U40972 (.A1(n49704), .A2(n24779), .ZN(N53844));
    NOR2X1 U40973 (.A1(n32805), .A2(n33272), .ZN(N53845));
    NANDX1 U40974 (.A1(N8186), .A2(N12493), .ZN(N53846));
    NOR2X1 U40975 (.A1(n13477), .A2(n49184), .ZN(N53847));
    INVX1 U40976 (.I(n19875), .ZN(N53848));
    NANDX1 U40977 (.A1(n26952), .A2(n13756), .ZN(N53849));
    INVX1 U40978 (.I(n27707), .ZN(N53850));
    INVX1 U40979 (.I(n25279), .ZN(N53851));
    INVX1 U40980 (.I(N10460), .ZN(N53852));
    NANDX1 U40981 (.A1(N8267), .A2(N10451), .ZN(N53853));
    INVX1 U40982 (.I(n14946), .ZN(N53854));
    NANDX1 U40983 (.A1(N6572), .A2(N6855), .ZN(N53855));
    NANDX1 U40984 (.A1(N2814), .A2(n22894), .ZN(N53856));
    INVX1 U40985 (.I(n26879), .ZN(N53857));
    INVX1 U40986 (.I(n16530), .ZN(N53858));
    NOR2X1 U40987 (.A1(n15196), .A2(N965), .ZN(N53859));
    NANDX1 U40988 (.A1(N2179), .A2(N10122), .ZN(N53860));
    NOR2X1 U40989 (.A1(n40914), .A2(n37074), .ZN(N53861));
    NANDX1 U40990 (.A1(N4015), .A2(N11319), .ZN(n53862));
    INVX1 U40991 (.I(n20554), .ZN(N53863));
    NOR2X1 U40992 (.A1(N11946), .A2(N7373), .ZN(N53864));
    INVX1 U40993 (.I(n13657), .ZN(N53865));
    NOR2X1 U40994 (.A1(n18089), .A2(N11059), .ZN(N53866));
    INVX1 U40995 (.I(n16204), .ZN(N53867));
    INVX1 U40996 (.I(n19198), .ZN(N53868));
    NOR2X1 U40997 (.A1(n30312), .A2(n46076), .ZN(N53869));
    NANDX1 U40998 (.A1(n38102), .A2(n18940), .ZN(N53870));
    NANDX1 U40999 (.A1(n30328), .A2(n50002), .ZN(N53871));
    NOR2X1 U41000 (.A1(n40449), .A2(N2755), .ZN(N53872));
    INVX1 U41001 (.I(n15322), .ZN(N53873));
    INVX1 U41002 (.I(n15685), .ZN(N53874));
    NOR2X1 U41003 (.A1(n15472), .A2(n27500), .ZN(N53875));
    NOR2X1 U41004 (.A1(n18678), .A2(n34872), .ZN(N53876));
    INVX1 U41005 (.I(n32334), .ZN(N53877));
    INVX1 U41006 (.I(n25270), .ZN(N53878));
    INVX1 U41007 (.I(n16346), .ZN(N53879));
    INVX1 U41008 (.I(n48556), .ZN(N53880));
    INVX1 U41009 (.I(n18370), .ZN(N53881));
    NANDX1 U41010 (.A1(n19419), .A2(n42692), .ZN(N53882));
    NOR2X1 U41011 (.A1(n29619), .A2(n20009), .ZN(N53883));
    NANDX1 U41012 (.A1(n26159), .A2(n52966), .ZN(N53884));
    NOR2X1 U41013 (.A1(n28913), .A2(N11176), .ZN(N53885));
    INVX1 U41014 (.I(n34159), .ZN(N53886));
    NANDX1 U41015 (.A1(n34367), .A2(n40891), .ZN(N53887));
    INVX1 U41016 (.I(n47144), .ZN(N53888));
    NANDX1 U41017 (.A1(n18292), .A2(N9604), .ZN(N53889));
    INVX1 U41018 (.I(n18254), .ZN(N53890));
    INVX1 U41019 (.I(N2154), .ZN(N53891));
    NANDX1 U41020 (.A1(n14146), .A2(n41971), .ZN(N53892));
    INVX1 U41021 (.I(n23776), .ZN(N53893));
    NOR2X1 U41022 (.A1(n18621), .A2(n13006), .ZN(N53894));
    NOR2X1 U41023 (.A1(n48239), .A2(n33014), .ZN(N53895));
    NOR2X1 U41024 (.A1(n20936), .A2(n23780), .ZN(N53896));
    NANDX1 U41025 (.A1(n41109), .A2(n34955), .ZN(N53897));
    NANDX1 U41026 (.A1(n21807), .A2(n44336), .ZN(N53898));
    NOR2X1 U41027 (.A1(N9236), .A2(n36495), .ZN(N53899));
    NOR2X1 U41028 (.A1(N6604), .A2(N1325), .ZN(N53900));
    INVX1 U41029 (.I(n27566), .ZN(N53901));
    NOR2X1 U41030 (.A1(n39835), .A2(n29719), .ZN(N53902));
    NANDX1 U41031 (.A1(n45241), .A2(n18228), .ZN(N53903));
    NANDX1 U41032 (.A1(n15555), .A2(n23404), .ZN(N53904));
    NOR2X1 U41033 (.A1(n19821), .A2(N12410), .ZN(N53905));
    NOR2X1 U41034 (.A1(n44096), .A2(n33050), .ZN(N53906));
    NANDX1 U41035 (.A1(n14414), .A2(N10112), .ZN(N53907));
    NANDX1 U41036 (.A1(n40629), .A2(n48361), .ZN(N53908));
    INVX1 U41037 (.I(n31503), .ZN(N53909));
    NOR2X1 U41038 (.A1(n45226), .A2(N5797), .ZN(N53910));
    NOR2X1 U41039 (.A1(n43090), .A2(n51843), .ZN(N53911));
    NOR2X1 U41040 (.A1(n17194), .A2(N481), .ZN(N53912));
    NANDX1 U41041 (.A1(n38174), .A2(n28440), .ZN(N53913));
    INVX1 U41042 (.I(N2940), .ZN(N53914));
    NANDX1 U41043 (.A1(N8083), .A2(n17605), .ZN(N53915));
    NOR2X1 U41044 (.A1(n27904), .A2(n30014), .ZN(N53916));
    NOR2X1 U41045 (.A1(n18538), .A2(N9602), .ZN(N53917));
    NANDX1 U41046 (.A1(n32951), .A2(N10974), .ZN(N53918));
    NOR2X1 U41047 (.A1(N11379), .A2(n50595), .ZN(N53919));
    INVX1 U41048 (.I(n42881), .ZN(N53920));
    NANDX1 U41049 (.A1(n41291), .A2(n48678), .ZN(N53921));
    INVX1 U41050 (.I(n30920), .ZN(N53922));
    NOR2X1 U41051 (.A1(n52454), .A2(n39374), .ZN(N53923));
    NANDX1 U41052 (.A1(n53203), .A2(n24086), .ZN(N53924));
    NANDX1 U41053 (.A1(n45731), .A2(n27026), .ZN(N53925));
    INVX1 U41054 (.I(N352), .ZN(N53926));
    INVX1 U41055 (.I(n37619), .ZN(N53927));
    NANDX1 U41056 (.A1(N12443), .A2(n46418), .ZN(N53928));
    INVX1 U41057 (.I(n13305), .ZN(N53929));
    NOR2X1 U41058 (.A1(N8803), .A2(n15539), .ZN(N53930));
    NANDX1 U41059 (.A1(N11442), .A2(N12672), .ZN(N53931));
    NOR2X1 U41060 (.A1(N862), .A2(n15121), .ZN(N53932));
    NANDX1 U41061 (.A1(n40800), .A2(n44460), .ZN(N53933));
    INVX1 U41062 (.I(n25658), .ZN(N53934));
    NOR2X1 U41063 (.A1(n51293), .A2(N2258), .ZN(N53935));
    INVX1 U41064 (.I(n21917), .ZN(N53936));
    NANDX1 U41065 (.A1(n17985), .A2(n48942), .ZN(N53937));
    INVX1 U41066 (.I(N9597), .ZN(N53938));
    NANDX1 U41067 (.A1(n52093), .A2(n29113), .ZN(N53939));
    INVX1 U41068 (.I(n45049), .ZN(N53940));
    INVX1 U41069 (.I(n39639), .ZN(N53941));
    NOR2X1 U41070 (.A1(N5029), .A2(N1716), .ZN(N53942));
    NANDX1 U41071 (.A1(n16470), .A2(N5649), .ZN(N53943));
    INVX1 U41072 (.I(N8592), .ZN(N53944));
    NOR2X1 U41073 (.A1(n17371), .A2(n40652), .ZN(N53945));
    INVX1 U41074 (.I(n29289), .ZN(N53946));
    INVX1 U41075 (.I(n37741), .ZN(N53947));
    INVX1 U41076 (.I(N6367), .ZN(N53948));
    INVX1 U41077 (.I(n40298), .ZN(N53949));
    INVX1 U41078 (.I(N10501), .ZN(N53950));
    NOR2X1 U41079 (.A1(n28138), .A2(n20098), .ZN(N53951));
    NANDX1 U41080 (.A1(n18030), .A2(n40471), .ZN(N53952));
    NOR2X1 U41081 (.A1(N879), .A2(n36696), .ZN(N53953));
    INVX1 U41082 (.I(n20757), .ZN(N53954));
    INVX1 U41083 (.I(N1698), .ZN(N53955));
    NOR2X1 U41084 (.A1(n49455), .A2(n52068), .ZN(N53956));
    INVX1 U41085 (.I(n49307), .ZN(N53957));
    NOR2X1 U41086 (.A1(n20542), .A2(n27759), .ZN(N53958));
    INVX1 U41087 (.I(n41092), .ZN(N53959));
    NANDX1 U41088 (.A1(n51404), .A2(N6011), .ZN(N53960));
    NOR2X1 U41089 (.A1(n52660), .A2(n46308), .ZN(N53961));
    NOR2X1 U41090 (.A1(N960), .A2(n19886), .ZN(N53962));
    INVX1 U41091 (.I(n21057), .ZN(N53963));
    NOR2X1 U41092 (.A1(n18386), .A2(N8066), .ZN(N53964));
    NOR2X1 U41093 (.A1(n38804), .A2(n34139), .ZN(N53965));
    NOR2X1 U41094 (.A1(N8859), .A2(n36670), .ZN(N53966));
    NOR2X1 U41095 (.A1(n33717), .A2(n19702), .ZN(N53967));
    INVX1 U41096 (.I(n16362), .ZN(N53968));
    NANDX1 U41097 (.A1(n16099), .A2(n33070), .ZN(N53969));
    NANDX1 U41098 (.A1(n20673), .A2(n40328), .ZN(N53970));
    NOR2X1 U41099 (.A1(n32478), .A2(N12124), .ZN(N53971));
    INVX1 U41100 (.I(n34126), .ZN(N53972));
    INVX1 U41101 (.I(n19919), .ZN(N53973));
    NANDX1 U41102 (.A1(n37589), .A2(n21174), .ZN(N53974));
    NANDX1 U41103 (.A1(n44287), .A2(n47758), .ZN(N53975));
    INVX1 U41104 (.I(n29280), .ZN(N53976));
    NANDX1 U41105 (.A1(n14271), .A2(n33581), .ZN(N53977));
    NOR2X1 U41106 (.A1(N10585), .A2(n32022), .ZN(N53978));
    NANDX1 U41107 (.A1(n27943), .A2(n49219), .ZN(N53979));
    NOR2X1 U41108 (.A1(n23234), .A2(n36375), .ZN(N53980));
    NANDX1 U41109 (.A1(N8454), .A2(n42998), .ZN(N53981));
    NANDX1 U41110 (.A1(n32003), .A2(n26969), .ZN(N53982));
    INVX1 U41111 (.I(n39769), .ZN(N53983));
    NOR2X1 U41112 (.A1(n13735), .A2(N5716), .ZN(N53984));
    NOR2X1 U41113 (.A1(n51323), .A2(n26890), .ZN(N53985));
    INVX1 U41114 (.I(N10109), .ZN(N53986));
    INVX1 U41115 (.I(n20156), .ZN(N53987));
    NOR2X1 U41116 (.A1(n18586), .A2(N2897), .ZN(N53988));
    NOR2X1 U41117 (.A1(N3112), .A2(n13481), .ZN(N53989));
    NOR2X1 U41118 (.A1(N868), .A2(N9895), .ZN(N53990));
    NOR2X1 U41119 (.A1(n19914), .A2(n33128), .ZN(N53991));
    NANDX1 U41120 (.A1(n26011), .A2(n41581), .ZN(N53992));
    INVX1 U41121 (.I(n27456), .ZN(N53993));
    INVX1 U41122 (.I(N4047), .ZN(N53994));
    INVX1 U41123 (.I(n27852), .ZN(n53995));
    NOR2X1 U41124 (.A1(N9374), .A2(n33567), .ZN(N53996));
    NOR2X1 U41125 (.A1(N6726), .A2(n28927), .ZN(N53997));
    NOR2X1 U41126 (.A1(n16834), .A2(n40515), .ZN(N53998));
    NOR2X1 U41127 (.A1(n24693), .A2(N5130), .ZN(N53999));
    INVX1 U41128 (.I(n43690), .ZN(N54000));
    INVX1 U41129 (.I(N2566), .ZN(N54001));
    NOR2X1 U41130 (.A1(N21), .A2(n34902), .ZN(N54002));
    NANDX1 U41131 (.A1(n19934), .A2(n14058), .ZN(N54003));
    INVX1 U41132 (.I(n14415), .ZN(N54004));
    NOR2X1 U41133 (.A1(n33958), .A2(n41870), .ZN(N54005));
    INVX1 U41134 (.I(N6475), .ZN(N54006));
    NOR2X1 U41135 (.A1(n40043), .A2(N8557), .ZN(N54007));
    NANDX1 U41136 (.A1(n42081), .A2(n36142), .ZN(N54008));
    NANDX1 U41137 (.A1(n39478), .A2(N2176), .ZN(N54009));
    NOR2X1 U41138 (.A1(n26022), .A2(n42335), .ZN(N54010));
    NOR2X1 U41139 (.A1(n31151), .A2(n53862), .ZN(N54011));
    NOR2X1 U41140 (.A1(n30304), .A2(n24898), .ZN(N54012));
    NANDX1 U41141 (.A1(n30324), .A2(N5828), .ZN(N54013));
    INVX1 U41142 (.I(n50257), .ZN(N54014));
    INVX1 U41143 (.I(n39678), .ZN(N54015));
    NANDX1 U41144 (.A1(n43993), .A2(n19664), .ZN(N54016));
    NANDX1 U41145 (.A1(n24656), .A2(n48580), .ZN(N54017));
    NANDX1 U41146 (.A1(N10727), .A2(N3166), .ZN(N54018));
    INVX1 U41147 (.I(n21278), .ZN(N54019));
    NOR2X1 U41148 (.A1(n42010), .A2(N6785), .ZN(N54020));
    NANDX1 U41149 (.A1(n26951), .A2(n32806), .ZN(N54021));
    INVX1 U41150 (.I(N5055), .ZN(N54022));
    NANDX1 U41151 (.A1(n20649), .A2(n26848), .ZN(N54023));
    NOR2X1 U41152 (.A1(n45546), .A2(n48761), .ZN(N54024));
    NOR2X1 U41153 (.A1(n51373), .A2(n31559), .ZN(N54025));
    INVX1 U41154 (.I(n17286), .ZN(N54026));
    NOR2X1 U41155 (.A1(N5450), .A2(n29749), .ZN(N54027));
    INVX1 U41156 (.I(n48931), .ZN(N54028));
    NANDX1 U41157 (.A1(n22450), .A2(n21980), .ZN(N54029));
    INVX1 U41158 (.I(n48057), .ZN(N54030));
    NOR2X1 U41159 (.A1(n23350), .A2(N1863), .ZN(N54031));
    NOR2X1 U41160 (.A1(n30134), .A2(N11816), .ZN(N54032));
    NANDX1 U41161 (.A1(n31410), .A2(n32574), .ZN(N54033));
    INVX1 U41162 (.I(n32307), .ZN(N54034));
    INVX1 U41163 (.I(n48186), .ZN(N54035));
    NANDX1 U41164 (.A1(n44796), .A2(n42975), .ZN(N54036));
    INVX1 U41165 (.I(N10668), .ZN(N54037));
    NOR2X1 U41166 (.A1(n43367), .A2(n27953), .ZN(N54038));
    NOR2X1 U41167 (.A1(n48816), .A2(n26172), .ZN(N54039));
    NANDX1 U41168 (.A1(n43776), .A2(n49047), .ZN(N54040));
    INVX1 U41169 (.I(n34226), .ZN(N54041));
    NOR2X1 U41170 (.A1(n19144), .A2(n22165), .ZN(N54042));
    INVX1 U41171 (.I(n21006), .ZN(N54043));
    INVX1 U41172 (.I(n19102), .ZN(N54044));
    NANDX1 U41173 (.A1(n14425), .A2(n50511), .ZN(N54045));
    INVX1 U41174 (.I(n35763), .ZN(N54046));
    NOR2X1 U41175 (.A1(N1586), .A2(n29977), .ZN(N54047));
    INVX1 U41176 (.I(n14852), .ZN(N54048));
    NANDX1 U41177 (.A1(n46383), .A2(n25519), .ZN(N54049));
    NANDX1 U41178 (.A1(n35778), .A2(n21942), .ZN(N54050));
    NANDX1 U41179 (.A1(n53065), .A2(n16585), .ZN(N54051));
    NOR2X1 U41180 (.A1(N11340), .A2(N11660), .ZN(N54052));
    NOR2X1 U41181 (.A1(n45565), .A2(n31249), .ZN(N54053));
    INVX1 U41182 (.I(n36200), .ZN(N54054));
    INVX1 U41183 (.I(n41510), .ZN(N54055));
    NANDX1 U41184 (.A1(n39317), .A2(N11273), .ZN(N54056));
    NOR2X1 U41185 (.A1(n35857), .A2(n45137), .ZN(N54057));
    INVX1 U41186 (.I(N1645), .ZN(N54058));
    NOR2X1 U41187 (.A1(n19917), .A2(N8497), .ZN(N54059));
    NANDX1 U41188 (.A1(N7367), .A2(N908), .ZN(N54060));
    INVX1 U41189 (.I(n37822), .ZN(N54061));
    NANDX1 U41190 (.A1(n14447), .A2(n43045), .ZN(N54062));
    NANDX1 U41191 (.A1(n31031), .A2(n19348), .ZN(N54063));
    NANDX1 U41192 (.A1(n42690), .A2(n52238), .ZN(N54064));
    INVX1 U41193 (.I(n42409), .ZN(N54065));
    NANDX1 U41194 (.A1(N2765), .A2(n40183), .ZN(N54066));
    NANDX1 U41195 (.A1(n50460), .A2(n25528), .ZN(N54067));
    INVX1 U41196 (.I(n27080), .ZN(N54068));
    NANDX1 U41197 (.A1(n53631), .A2(n17020), .ZN(N54069));
    INVX1 U41198 (.I(n37295), .ZN(n54070));
    INVX1 U41199 (.I(N8467), .ZN(N54071));
    NOR2X1 U41200 (.A1(n35216), .A2(n31816), .ZN(N54072));
    NOR2X1 U41201 (.A1(n41508), .A2(N5443), .ZN(N54073));
    INVX1 U41202 (.I(n53023), .ZN(N54074));
    NANDX1 U41203 (.A1(n19821), .A2(n18399), .ZN(N54075));
    NOR2X1 U41204 (.A1(N8540), .A2(n16665), .ZN(N54076));
    NOR2X1 U41205 (.A1(n50948), .A2(N3906), .ZN(N54077));
    INVX1 U41206 (.I(N5630), .ZN(N54078));
    NANDX1 U41207 (.A1(n49337), .A2(n53600), .ZN(N54079));
    NOR2X1 U41208 (.A1(n44887), .A2(n51925), .ZN(N54080));
    NANDX1 U41209 (.A1(N7936), .A2(n51895), .ZN(N54081));
    NOR2X1 U41210 (.A1(n35784), .A2(n28832), .ZN(N54082));
    NOR2X1 U41211 (.A1(n39470), .A2(n29118), .ZN(N54083));
    NOR2X1 U41212 (.A1(n27006), .A2(N3032), .ZN(N54084));
    INVX1 U41213 (.I(n26057), .ZN(N54085));
    INVX1 U41214 (.I(n33808), .ZN(N54086));
    NOR2X1 U41215 (.A1(N10742), .A2(n42347), .ZN(N54087));
    INVX1 U41216 (.I(n38383), .ZN(N54088));
    INVX1 U41217 (.I(n33495), .ZN(N54089));
    INVX1 U41218 (.I(n35866), .ZN(N54090));
    NOR2X1 U41219 (.A1(N1096), .A2(N3965), .ZN(N54091));
    NOR2X1 U41220 (.A1(n45982), .A2(N1919), .ZN(N54092));
    INVX1 U41221 (.I(n22388), .ZN(N54093));
    NOR2X1 U41222 (.A1(n37036), .A2(n26643), .ZN(N54094));
    INVX1 U41223 (.I(n33918), .ZN(N54095));
    NOR2X1 U41224 (.A1(n48703), .A2(N5144), .ZN(N54096));
    INVX1 U41225 (.I(n51734), .ZN(N54097));
    INVX1 U41226 (.I(N11232), .ZN(N54098));
    NOR2X1 U41227 (.A1(n52939), .A2(N1716), .ZN(N54099));
    NOR2X1 U41228 (.A1(N9785), .A2(n31305), .ZN(N54100));
    NOR2X1 U41229 (.A1(n40021), .A2(n33271), .ZN(N54101));
    NOR2X1 U41230 (.A1(n44358), .A2(N4834), .ZN(N54102));
    NANDX1 U41231 (.A1(n48322), .A2(n17546), .ZN(N54103));
    INVX1 U41232 (.I(n18711), .ZN(N54104));
    NANDX1 U41233 (.A1(N8687), .A2(N9465), .ZN(N54105));
    NANDX1 U41234 (.A1(N3800), .A2(n29050), .ZN(N54106));
    NANDX1 U41235 (.A1(n15941), .A2(n46224), .ZN(N54107));
    NOR2X1 U41236 (.A1(N1116), .A2(N12457), .ZN(N54108));
    NOR2X1 U41237 (.A1(N12347), .A2(n36297), .ZN(N54109));
    NOR2X1 U41238 (.A1(n36504), .A2(n16907), .ZN(N54110));
    NOR2X1 U41239 (.A1(n36280), .A2(N4371), .ZN(N54111));
    NANDX1 U41240 (.A1(n15579), .A2(n51535), .ZN(N54112));
    INVX1 U41241 (.I(n20412), .ZN(N54113));
    NOR2X1 U41242 (.A1(n33069), .A2(N6428), .ZN(N54114));
    NOR2X1 U41243 (.A1(n20250), .A2(n14435), .ZN(N54115));
    NOR2X1 U41244 (.A1(n29715), .A2(N5506), .ZN(N54116));
    INVX1 U41245 (.I(n27235), .ZN(N54117));
    INVX1 U41246 (.I(n51462), .ZN(N54118));
    NANDX1 U41247 (.A1(n42452), .A2(n52577), .ZN(N54119));
    NANDX1 U41248 (.A1(n51099), .A2(n33394), .ZN(N54120));
    NOR2X1 U41249 (.A1(n27183), .A2(n15927), .ZN(N54121));
    NANDX1 U41250 (.A1(n13052), .A2(n52206), .ZN(N54122));
    NOR2X1 U41251 (.A1(N7413), .A2(n36255), .ZN(N54123));
    NOR2X1 U41252 (.A1(n46130), .A2(N2695), .ZN(N54124));
    NOR2X1 U41253 (.A1(n47669), .A2(n31564), .ZN(N54125));
    NOR2X1 U41254 (.A1(n13948), .A2(n45998), .ZN(N54126));
    INVX1 U41255 (.I(N12133), .ZN(N54127));
    NOR2X1 U41256 (.A1(n52181), .A2(n39367), .ZN(N54128));
    NOR2X1 U41257 (.A1(n49671), .A2(n27325), .ZN(N54129));
    INVX1 U41258 (.I(n48276), .ZN(N54130));
    INVX1 U41259 (.I(n17901), .ZN(N54131));
    NOR2X1 U41260 (.A1(n42007), .A2(n45083), .ZN(N54132));
    NANDX1 U41261 (.A1(N10124), .A2(N4164), .ZN(N54133));
    NOR2X1 U41262 (.A1(n36582), .A2(n34018), .ZN(N54134));
    NANDX1 U41263 (.A1(n29075), .A2(n26176), .ZN(N54135));
    NOR2X1 U41264 (.A1(n13419), .A2(n42316), .ZN(N54136));
    NOR2X1 U41265 (.A1(n52328), .A2(n24734), .ZN(N54137));
    INVX1 U41266 (.I(n15016), .ZN(N54138));
    NOR2X1 U41267 (.A1(n29781), .A2(n35667), .ZN(N54139));
    NOR2X1 U41268 (.A1(n39632), .A2(n31366), .ZN(N54140));
    NANDX1 U41269 (.A1(n37963), .A2(n48112), .ZN(N54141));
    NOR2X1 U41270 (.A1(N1892), .A2(n44280), .ZN(N54142));
    NANDX1 U41271 (.A1(n15445), .A2(N2404), .ZN(N54143));
    INVX1 U41272 (.I(n42050), .ZN(N54144));
    INVX1 U41273 (.I(n17477), .ZN(N54145));
    INVX1 U41274 (.I(n50228), .ZN(N54146));
    INVX1 U41275 (.I(n16743), .ZN(N54147));
    INVX1 U41276 (.I(n28440), .ZN(N54148));
    NOR2X1 U41277 (.A1(N257), .A2(n49238), .ZN(N54149));
    NOR2X1 U41278 (.A1(N10064), .A2(n32724), .ZN(N54150));
    NOR2X1 U41279 (.A1(n39845), .A2(n14419), .ZN(N54151));
    NOR2X1 U41280 (.A1(n47947), .A2(n14255), .ZN(N54152));
    NOR2X1 U41281 (.A1(n31938), .A2(N8395), .ZN(N54153));
    NOR2X1 U41282 (.A1(N2300), .A2(n21146), .ZN(N54154));
    INVX1 U41283 (.I(n40186), .ZN(N54155));
    NOR2X1 U41284 (.A1(N786), .A2(n28265), .ZN(N54156));
    INVX1 U41285 (.I(n40704), .ZN(N54157));
    INVX1 U41286 (.I(n23449), .ZN(N54158));
    INVX1 U41287 (.I(N4044), .ZN(N54159));
    NANDX1 U41288 (.A1(n52635), .A2(n31572), .ZN(N54160));
    INVX1 U41289 (.I(n47902), .ZN(N54161));
    NOR2X1 U41290 (.A1(n38685), .A2(n49096), .ZN(N54162));
    NANDX1 U41291 (.A1(n47000), .A2(n31986), .ZN(N54163));
    NANDX1 U41292 (.A1(n40975), .A2(n46240), .ZN(N54164));
    INVX1 U41293 (.I(n41383), .ZN(N54165));
    NANDX1 U41294 (.A1(n39675), .A2(N12153), .ZN(N54166));
    INVX1 U41295 (.I(n28037), .ZN(N54167));
    NANDX1 U41296 (.A1(n36270), .A2(n51264), .ZN(N54168));
    NANDX1 U41297 (.A1(N9491), .A2(n37996), .ZN(N54169));
    NOR2X1 U41298 (.A1(N1411), .A2(n39749), .ZN(N54170));
    INVX1 U41299 (.I(n29776), .ZN(N54171));
    NANDX1 U41300 (.A1(n18019), .A2(N4426), .ZN(N54172));
    NOR2X1 U41301 (.A1(n16352), .A2(N11581), .ZN(N54173));
    INVX1 U41302 (.I(n40752), .ZN(N54174));
    NANDX1 U41303 (.A1(n18836), .A2(n27981), .ZN(N54175));
    NANDX1 U41304 (.A1(N11104), .A2(n18536), .ZN(N54176));
    NANDX1 U41305 (.A1(N2680), .A2(N4240), .ZN(N54177));
    INVX1 U41306 (.I(n46930), .ZN(N54178));
    INVX1 U41307 (.I(N2899), .ZN(N54179));
    NANDX1 U41308 (.A1(n52010), .A2(n51972), .ZN(N54180));
    NOR2X1 U41309 (.A1(n36034), .A2(N2847), .ZN(N54181));
    NANDX1 U41310 (.A1(n44253), .A2(n43265), .ZN(N54182));
    INVX1 U41311 (.I(n19606), .ZN(N54183));
    NANDX1 U41312 (.A1(N11271), .A2(n42861), .ZN(N54184));
    NANDX1 U41313 (.A1(n22851), .A2(N7269), .ZN(N54185));
    INVX1 U41314 (.I(n49902), .ZN(N54186));
    NOR2X1 U41315 (.A1(n29337), .A2(N9986), .ZN(N54187));
    NANDX1 U41316 (.A1(n47873), .A2(n33894), .ZN(N54188));
    NOR2X1 U41317 (.A1(n20583), .A2(n15983), .ZN(N54189));
    INVX1 U41318 (.I(n43771), .ZN(N54190));
    NOR2X1 U41319 (.A1(n43899), .A2(n41809), .ZN(N54191));
    NOR2X1 U41320 (.A1(n51088), .A2(n46313), .ZN(N54192));
    NANDX1 U41321 (.A1(n28158), .A2(N5065), .ZN(N54193));
    NOR2X1 U41322 (.A1(n35003), .A2(n24670), .ZN(N54194));
    NOR2X1 U41323 (.A1(n53232), .A2(n49762), .ZN(N54195));
    NANDX1 U41324 (.A1(N2652), .A2(n16181), .ZN(N54196));
    NOR2X1 U41325 (.A1(N1836), .A2(N2872), .ZN(N54197));
    NOR2X1 U41326 (.A1(n51196), .A2(n13455), .ZN(N54198));
    INVX1 U41327 (.I(N10886), .ZN(N54199));
    INVX1 U41328 (.I(N2766), .ZN(N54200));
    NANDX1 U41329 (.A1(n46062), .A2(n45239), .ZN(N54201));
    INVX1 U41330 (.I(n23864), .ZN(N54202));
    NOR2X1 U41331 (.A1(n38534), .A2(N6555), .ZN(N54203));
    INVX1 U41332 (.I(n23301), .ZN(N54204));
    INVX1 U41333 (.I(n18497), .ZN(N54205));
    INVX1 U41334 (.I(n49029), .ZN(N54206));
    NOR2X1 U41335 (.A1(N3078), .A2(N1669), .ZN(N54207));
    NOR2X1 U41336 (.A1(n19643), .A2(N4320), .ZN(N54208));
    NANDX1 U41337 (.A1(n16343), .A2(n13952), .ZN(N54209));
    INVX1 U41338 (.I(N5599), .ZN(N54210));
    INVX1 U41339 (.I(n34509), .ZN(N54211));
    NOR2X1 U41340 (.A1(n29634), .A2(n19133), .ZN(N54212));
    NOR2X1 U41341 (.A1(n13604), .A2(n18796), .ZN(N54213));
    NANDX1 U41342 (.A1(n30814), .A2(n50455), .ZN(N54214));
    NANDX1 U41343 (.A1(n22949), .A2(N10611), .ZN(N54215));
    NANDX1 U41344 (.A1(n46250), .A2(N3049), .ZN(N54216));
    INVX1 U41345 (.I(n50917), .ZN(N54217));
    NOR2X1 U41346 (.A1(N5669), .A2(n53995), .ZN(N54218));
    NOR2X1 U41347 (.A1(n54070), .A2(n27239), .ZN(N54219));
    INVX1 U41348 (.I(n18059), .ZN(N54220));
    NANDX1 U41349 (.A1(n34617), .A2(N9449), .ZN(N54221));
    NANDX1 U41350 (.A1(N11055), .A2(n42891), .ZN(N54222));
    INVX1 U41351 (.I(N3811), .ZN(N54223));
    NOR2X1 U41352 (.A1(N12722), .A2(n37132), .ZN(N54224));
    NANDX1 U41353 (.A1(n46033), .A2(n48520), .ZN(N54225));
    INVX1 U41354 (.I(n32242), .ZN(N54226));
    NOR2X1 U41355 (.A1(N6775), .A2(n17139), .ZN(N54227));
    NANDX1 U41356 (.A1(n18038), .A2(n50199), .ZN(N54228));
    INVX1 U41357 (.I(N7737), .ZN(N54229));
    NANDX1 U41358 (.A1(n41163), .A2(n33148), .ZN(N54230));
    INVX1 U41359 (.I(N6101), .ZN(N54231));
    INVX1 U41360 (.I(n35297), .ZN(N54232));
    INVX1 U41361 (.I(n20498), .ZN(N54233));
    NOR2X1 U41362 (.A1(n33333), .A2(n31552), .ZN(N54234));
    NOR2X1 U41363 (.A1(N317), .A2(n43254), .ZN(N54235));
    NANDX1 U41364 (.A1(N2092), .A2(N11849), .ZN(N54236));
    NOR2X1 U41365 (.A1(N7411), .A2(N2569), .ZN(N54237));
    NOR2X1 U41366 (.A1(n45785), .A2(N5403), .ZN(N54238));
    NANDX1 U41367 (.A1(n40814), .A2(n43202), .ZN(N54239));
    NOR2X1 U41368 (.A1(N3932), .A2(n18525), .ZN(N54240));
    INVX1 U41369 (.I(n50423), .ZN(N54241));
    NOR2X1 U41370 (.A1(n51337), .A2(n45306), .ZN(N54242));
    NOR2X1 U41371 (.A1(n33172), .A2(n52605), .ZN(N54243));
    NANDX1 U41372 (.A1(N636), .A2(n26648), .ZN(N54244));
    NOR2X1 U41373 (.A1(n39114), .A2(n47717), .ZN(N54245));
    NOR2X1 U41374 (.A1(n44720), .A2(n26607), .ZN(N54246));
    NANDX1 U41375 (.A1(N7808), .A2(n40690), .ZN(N54247));
    NANDX1 U41376 (.A1(n42709), .A2(n15912), .ZN(N54248));
    NOR2X1 U41377 (.A1(n19572), .A2(n21683), .ZN(N54249));
    NANDX1 U41378 (.A1(N8535), .A2(N9212), .ZN(N54250));
    NOR2X1 U41379 (.A1(n42783), .A2(n50568), .ZN(N54251));
    NANDX1 U41380 (.A1(n44490), .A2(N9153), .ZN(N54252));
    NOR2X1 U41381 (.A1(n14395), .A2(n42324), .ZN(N54253));
    NANDX1 U41382 (.A1(n24282), .A2(n42960), .ZN(N54254));
    NANDX1 U41383 (.A1(n39072), .A2(n43559), .ZN(N54255));
    NOR2X1 U41384 (.A1(n53392), .A2(n49764), .ZN(N54256));
    NANDX1 U41385 (.A1(n24934), .A2(N3333), .ZN(N54257));
    INVX1 U41386 (.I(n13537), .ZN(N54258));
    NANDX1 U41387 (.A1(n19903), .A2(n53799), .ZN(N54259));
    NOR2X1 U41388 (.A1(N3072), .A2(n42122), .ZN(N54260));
    INVX1 U41389 (.I(N12283), .ZN(N54261));
    NANDX1 U41390 (.A1(N1387), .A2(n24336), .ZN(N54262));
    NOR2X1 U41391 (.A1(N7362), .A2(n33488), .ZN(N54263));
    NOR2X1 U41392 (.A1(n21756), .A2(n37298), .ZN(N54264));
    NANDX1 U41393 (.A1(N7524), .A2(n26019), .ZN(N54265));
    NOR2X1 U41394 (.A1(n46595), .A2(n31063), .ZN(N54266));
    NOR2X1 U41395 (.A1(N7235), .A2(n26589), .ZN(N54267));
    NANDX1 U41396 (.A1(n32168), .A2(n45645), .ZN(N54268));
    NOR2X1 U41397 (.A1(n45704), .A2(n14658), .ZN(N54269));
    NANDX1 U41398 (.A1(n45264), .A2(N3241), .ZN(N54270));
    NANDX1 U41399 (.A1(n23827), .A2(N6988), .ZN(N54271));
    INVX1 U41400 (.I(n28390), .ZN(N54272));
    NOR2X1 U41401 (.A1(n43627), .A2(n13251), .ZN(N54273));
    NOR2X1 U41402 (.A1(n18652), .A2(n26927), .ZN(N54274));
    INVX1 U41403 (.I(N8324), .ZN(N54275));
    NANDX1 U41404 (.A1(N1216), .A2(n35685), .ZN(N54276));
    NOR2X1 U41405 (.A1(N8081), .A2(n32612), .ZN(N54277));
    INVX1 U41406 (.I(n34269), .ZN(N54278));
    INVX1 U41407 (.I(N2343), .ZN(N54279));
    INVX1 U41408 (.I(n35157), .ZN(N54280));
    INVX1 U41409 (.I(n31090), .ZN(N54281));
    NANDX1 U41410 (.A1(n32248), .A2(n47375), .ZN(N54282));
    NOR2X1 U41411 (.A1(n43017), .A2(n16931), .ZN(N54283));
    NANDX1 U41412 (.A1(n45943), .A2(n25572), .ZN(N54284));
    INVX1 U41413 (.I(n15551), .ZN(N54285));
    INVX1 U41414 (.I(N796), .ZN(N54286));
    NOR2X1 U41415 (.A1(n26253), .A2(n36324), .ZN(N54287));
    NANDX1 U41416 (.A1(n14002), .A2(n37539), .ZN(N54288));
    INVX1 U41417 (.I(N1317), .ZN(N54289));
    NANDX1 U41418 (.A1(n17056), .A2(n16271), .ZN(N54290));
    INVX1 U41419 (.I(n13984), .ZN(N54291));
    NANDX1 U41420 (.A1(n31952), .A2(n29393), .ZN(N54292));
    NANDX1 U41421 (.A1(n43293), .A2(N3112), .ZN(N54293));
    NOR2X1 U41422 (.A1(n36397), .A2(n27006), .ZN(N54294));
    NOR2X1 U41423 (.A1(n33580), .A2(n38140), .ZN(N54295));
    INVX1 U41424 (.I(N4881), .ZN(N54296));
    NANDX1 U41425 (.A1(N9431), .A2(n23955), .ZN(N54297));
    NOR2X1 U41426 (.A1(n43633), .A2(n50207), .ZN(N54298));
    NANDX1 U41427 (.A1(n46663), .A2(N9938), .ZN(N54299));
    NANDX1 U41428 (.A1(n50854), .A2(n45777), .ZN(N54300));
    INVX1 U41429 (.I(n13639), .ZN(N54301));
    INVX1 U41430 (.I(n23027), .ZN(N54302));
    NOR2X1 U41431 (.A1(N6641), .A2(N708), .ZN(N54303));
    INVX1 U41432 (.I(N7604), .ZN(N54304));
    NOR2X1 U41433 (.A1(n40378), .A2(N6292), .ZN(N54305));
    INVX1 U41434 (.I(n47635), .ZN(N54306));
    INVX1 U41435 (.I(n23061), .ZN(N54307));
    INVX1 U41436 (.I(n33913), .ZN(N54308));
    INVX1 U41437 (.I(n17478), .ZN(N54309));
    INVX1 U41438 (.I(n29689), .ZN(N54310));
    NANDX1 U41439 (.A1(n33048), .A2(n51192), .ZN(N54311));
    NANDX1 U41440 (.A1(n51227), .A2(n39476), .ZN(N54312));
    NOR2X1 U41441 (.A1(N5057), .A2(n28284), .ZN(N54313));
    INVX1 U41442 (.I(n46259), .ZN(N54314));
    INVX1 U41443 (.I(n33883), .ZN(N54315));
    NANDX1 U41444 (.A1(n50686), .A2(n35867), .ZN(N54316));
    NOR2X1 U41445 (.A1(N9616), .A2(N9858), .ZN(N54317));
    INVX1 U41446 (.I(n36658), .ZN(N54318));
    INVX1 U41447 (.I(n47132), .ZN(N54319));
    NOR2X1 U41448 (.A1(n45596), .A2(N1806), .ZN(N54320));
    NANDX1 U41449 (.A1(n47715), .A2(n27674), .ZN(N54321));
endmodule
